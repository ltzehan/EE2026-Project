`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ihvl9qvl6mtGSCn2QmTq24p+4WK+wehYw2BbTxVxOCa6AomXDDHWk3N+fCT7Ec6ymOwaE84zl0AE
FfZ+2lebag==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AHSEaMSHfcPE7ySf3fWQlVVbNBrSBwx7+2AARSD3OQbYwQqttf2jqz1AS0VS/c8hbcCH5/xEo6wc
0YCLC0TLjuP2NG+0xTTkINJp9RP36eLtRQ2gjEU9+Pygg4ojLhxKahp/JEhqwbC1zJ0m6z6tXz28
bTJx42bN7mGmsF/5Vgo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eUgf8tzJSzGYR4YGwogvvkQDrltsQcVA9ax6H/7FMeGxBK2ExpkrnTayKuSWcrEPmKPLWojzX4Rp
jrntLR03FJ33vvdw2iwqsMr+YZSn0FiWqFMgiPpkhPbKlP4d15bbtMD1Gko6ThnUYsNe1Uokkn4j
XnzAaz7aLS/P1FfaZrZVJLZBmqw+M4M3WTQh3kHKZi1NfWDWFanvoTIJ8umhWll7zTiRIxxlj2sf
1AcaTjGRqpbPx1fswKwB7zjTxMYAB6XDrFCMn5GWHrXicRi1BSZ1dc9X0RaAEy2+fbCe/QSMIv19
MDudZjBjTBvKNBHTvAxVaCQR/r6TjwYyPHNUow==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fCE0iqQqQmMaiqxfu+lTOtYiRgejwUsC7ex66qrLPjZOeOOR6VFQe0j18JJeWW1cqE1CqiDHXXhL
6qtSICA9OSpeVggF9+AotqgyKE2nkxSN+OH8BinQb+BCes2TzJdC0Q8T8bvLRGMoliywPlIhdI6M
pVGSFhdws+piimMdaiPwhMLA0wE+YYK+4mN+QesiOMEQp3/Cv4ACToB5iiqSUx8R1uBNs+IBsaLd
CAPHniHtsT0elqUJOwqg9qiDbSvuE6UgMnvSrPAsFvL62QdWpPybBWyfKrhItzQnrneRgsJNsmbD
TdnUyZ73dN5jp+L64ScrCI3oJTqLgQ/GAoegqQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KP8tDEaMtNiHb7fLSQNSmIn6f3quyU2/8znjyIPJk9gEjSsUmr7PpaLzh7KITyetyAykLNDy0+If
oi9FlchUdYS1S8pIc+xKb4AysqoPNQ+I+BYMgLboZ2BRi67NmSNSZYIhupYI3kmhhdoBdG0KzW7A
Aa4Qz9i9rgI0nLPReO8LZ1al6lYDHDry02cDN+z+OiGpkpvQiPH1p/hGXvKiTMWnkZNiRGteD3q8
NidKjK7vDwMwTVfAhWlaTHlCguRO0FMdED3Flrh0oUCH2MyAsCHNAsNEF/4qI+Lk3OL1BLUoHCO/
hHnZPWSiBfVLKyuWqMN3Hqm/+H7K+iaKo2cU/A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VYINJP/X0xCgvLZxQq9WoLczB1D4IDZ/fiNpsohtGnTSTTQAZTTkHNgUYHINe8Hnm+sHY/z+79mf
SZmevlmaMyfQ/bruVpg7xkGk0kbsRE0657dK7+oA8vBZP50PGrnmyAUz9JthH6ARIL//Z+jFQIOm
3AEyJSkfolORpd6jmrA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BCuflP0+YszOWk6oPUbw/aQvnws00cRjSsHJnmgdFgTaszbu6AWa6hxrBP5OsH4RBPYxnsCAzzmv
F5qT51GZNkOOZdTFTAcngBKxoMJSIxiAaRhxchN7P0V+S0FF7xLP/fGcJOqyFT6KpjP/RTwm3vUe
xD8zDgnEwlNjVHzIqTKpFHYOSL3LJUDoF1rbjBDNfrVak1lMu0CVMwqb+wnGLhRZ1UjS/sXTSCp+
vZNSonNgI1muW5JsxMZapVVzl8zcz4B4MQirD3E8dZylgZJrpaW5nyfCS6axpHQXarqv+DjNU4u9
nolZ1lTfG/mT8DJpdiBfhnV1wNBkgF9/OFqaIw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1558368)
`protect data_block
hJ65tJJqeWzVMBLB/s8+gBjBymuiuUUS5Hia0vJDVvdsI4gpBjtF2sNkpKQA630bxxk+RdyfcoAd
yRAvNDU2CyLROUlas6DJamSfHzyrn0QiFmfGvmvOe00TmuI72LIH4UrF9p9BHiHnR3HHmst/Gp27
atJvXJsBWojZGN68rD1tNaTkmwi94IZWfoP2T1eAY3foEyOU2HVyp8PGqepx170KkdMj82jXfRVM
69wF3oOdnjpM9bEtbCYeWlSot+zZo34plic1pyAkUI3pUhcjVehE9p58c2/UywV0g3poqIVF0iQ1
0zcSchXUbeEeeZWj4qdc+L7UeAZn6HTtkLZ4M8Sz+nP9K9jGAEpuQy4Im05d2EqRGkCQkGp0Tfci
7sov+sBSNrKVol7bflNemMZn/6D5to8reGXqv0PM1GCYY5Ggssajew0VqRUln3cfvrT0201oP/2h
YAgJUJgRqauKrBUbr1/2lZ+aIYles94+LqnFCwDN22JhC88UAJqfxN9pTeKsUEX3pyw3RxaQlPHl
E/Uox+gfVU2oKlGV1QRToyoPwj8xTIhaG9SMrwO3WgmtAaEbkOZcN4RbkwCjyM1D6FIwZqWEK0ia
d1woO8g2DF2Pv0sU6qV8ACCNhvg1/eVEY30M68wOU/+j8dT8mDBivjNS9FZVNQjEDbrLnUbkArKC
PuRnb75QZOI8NYMnvuQ0nyTwH/Iqnp3IrjMjRNcAekL54+LqLvoahTRbE77jJngq77gBnDAtrRXr
W/UKp5ZBGGWT8mkL4/mo/IBzcbebv20Db0b8S/hxpRlwa06M5fpMXo4OKJU5ZNxfXNVZPTJHmOle
LpBonVPBjw8+w5xLc2GlnhvPDCoPCbspo9A7FifIVOGIU8/pk1XRbp0C1Mpn6TEngqLoHSbQsdnQ
frMVaxZ9IjnYSdyvtp9M0kf+F5YbDX809BNdCU+/n6sD9FtmksBrP12oT3ODQuWOTV4WLLL+wmvl
crW0WPOZYXqStXpNSyjYKyjcTEsdThPKAO2hrzcyGkYkMQF9YacFPgkWdWxGFCtfP982SQzxl+FG
ygIp5U7RCbeTzxpXBwyYGm+p0m/PsHnieyAmkesbJHowvMvlSQUw5Q7SoVnUSpyVV5vqG3DwnSDO
/4OnfZKi4jkwbUEnKgmpqAI/c80HaJCiprACPrZw5vbfvrqw/cT6OHLPXMwssddVGBQdz9gh4Brt
Yjq3vHZrC0puS/xZ7t5RiTJEAEpE/C/dGm+cWvyaVyON9xTLJthe7yWx0AYHFoKCFRDfFQkkK0w7
8//iDjrKqh1j6vihiri8y44+X4iNk79vGThvZ1VAFzIFqg7yVfyp3d3ci4hPA2B+bLCuzpUCUr2p
xG7IXyQo49iEE+aoCk29ZNpdYXYPPqTS3KY1S9wa6wEkQXd+U4IPAUAWP03Y6hdGBiV8A4XtOOsX
eRzgz6C9S2ppYnrDWA+lUYU9T+MLgwyeTuCLqmA4v4xiAivEs3DPy6mKSE/VFEKVGEa6GmAv4mgi
Ykm8ycCpWGTz8cPVKu6vVWkoLDhm/yFkOLKJ2RrX+SIlvjFqTUsga+ef6UTLFwfKbXGiC+znbK8P
K70Q8Zft97sZ030ETCKnm4J+mjKHTglgW1vYGQGYp1gGibT+G1aIuHBNbfkC1YwSULuXo03IVWPo
xpikPAlJIuwCv81oa0BINBeoeiT/P4LO5/iZHzDDbGdyqPSC5DSoiMpz/wVqXk7yJn5wmkqhDiyf
HrOnqXD6N2iAyegqIv0nwcbG9opNn6j4rqD5bpsE2h8Iq4tx2ItCPX2xq7hTudAphyzbxoJW1dqx
Gev7ROTo6pRonqdiNjuGDGx8PW6EZtttexuak/5yLVDyt0X6f79DJsnnUgVGs6KY2vzD9XJFJEY9
4aFv8FHC9dvPcWIJwr7GmT6IHz4lIyVz4mXqoa4UcuZ7MVxPgp/5L9bkwRO78vrGKkMo8uo9Kx5f
of46SGRt5OQ3L49/jd82gNvo7f72y4sfVC7zllSiOLUio+dlXPEsqyC8hEbx7dR/bu4ftrE5LShV
NnrOkoMZjZWDPH44ceU+g5jUaC72OR3t46GP2OkImFCO1ST4C9Qmb+2DCdCa/cKup9LUlp8VGhAz
JlnaPA/TsoIbhrsNJiJv3kzBtzR/AeV5GjyoMYja0YxFE6oEtZ9116kPJd+vf18/0fBwtIx7Sz4f
5MizOQ8lwXvuZuAttyq08bhvuLC125/p/teabuA4ZmIdKlUcJWawxfO1//CrU3r84nYZpXy9ZwaE
+9+JTj6LdLCSPLX4W+UMe7XJ0y/cBM/YyHGj7GXmTtIWCZygkUXfFQwqk+sg+jIp4yF5kz79HrkL
9sqNNzXv7CqWv5Ha6GbhCxAOME1PHk+qDfA46fJWUOPSiX/0xYM2qJbxqqB+bulnsfH4dfSayLNq
V6W/ijJQ8jvkIwUnFNmbLU0j8200yQrP9QdUoS7jAok07m4SXjsqifPo16Wus7qZX/o8V0YAQ7U2
gjc2FBAgWUJdK6Y2lcf7lwMK5M8yiXakriytXdgKfy0mbOR8RsSSTXTetlHNppPwd6YtX1StmJoV
NzunCEI/DTgqV3BiXpnhDL/8t+TWuel1kHP0iVe1EEtJFUUecQCISpa4vihPXwQm5SleskVumhoB
IHcA4ohd4AvlEKc8Jzg51aYWlc4fgqIPALYPNp8nvrU+yyNsGbKo1EDExc6oc4BPQT24Fsu/fob+
wbEjWhWLFSkPiPf75Wi7bIglpBlxvN1rictae+MBsGUrIt44RB+kyjSJIKckaLG9Fr/vLDs4UTmG
a3ZakZZG7VaOkdkQc63IIZTjkfymxOHmVwncfo88gNwmLuZgcj5cIDg7TRVOq3Zvd6i9oS841qvk
sn5Z+mszKq2lP/s7JoFZRXyA9hc9SxRA0h+2RfEbs1mTUmfc+rJbKpvT+wvfQ/NsQVjvyU9wdrm5
3iffvgzJjiOv2IrDVEQBF7AWAGd7axi4+erZQ95rUxIZ1++mtdcBMdCr0HqL2EmDVv9kk+jbXcMV
1In0SLJn5Gg3Amc5DnwzzZbkz5YzH/qLidsmk1xGYuD9KlJa8xK9yDpJB8vAUFiuohvBqFkEpmDO
UqB1ahLMqjO0/tbWmLN3hwfH84pt+VKzejM3njolgwNDXcunGeCRG2LnUoQAqZvZyEJb3WWv+aGi
M52eiLThy22WUoFJv8qI3GLIyiIHs0Vka9zVdH+UYbKJhjeBkQq3qWlAwBTa0tWl/AbWqTYg9JJQ
IgW2EXcDj0peke6lVKE1kJmJUuMCZGeZhMZ/VXnzAtX4RXgz6lgTCsOKGqoUrf0BaiMR1xyoAjLM
JCw8x7n1G0ifMmZufU3Vdun4noA6hyiVjtYGgyoSBDaUl96oB6PBb77mFhXnZH+b8WYrS4n8Zxg0
QhIJlGaMCH0mIccvp61t9rUQrI0F2fNMwQPbViso4FINhoW/5zvkNqPAxg5BHh29iLpdW5XcELMl
Luayz+pBG/xRxt7jaE6WzoiudAtZA97jNF6LyYBfFOAKurF6fTShZxzqY8xOoln4t/bepEtkiAlN
LCTu6wcjlnvYhe9hJODMgmAySJP56CajPOP3kYUgQXeaS8Lhoi6HnFY2UKSK8812fuU/G/fx0JBI
lWcGHR0arSRM5FB8KIsEC1TVTnl0coXPrQ2HiNvTXybxpyx+n2auBsUj+nb86aNAZH+JG2dZvL6z
5Y+LRb5ZVGRhCrKKgYMPRRGLiw/Qgv2UpKrHzmPavDgALUqWZI+ZUoi69R36s6+TqjehVWPsiQ03
iAQ6Gt8o7iWeN+PJwK58MVPEVyxw8ij+GgNF5ZE115FfKC+p557BJ1cF+GVH6wlzcnQm9PVphGE7
l503ysPTLwCgN9GEPWnskgj0ce6QZEHLpMjQaccIQx5i3C28lyOvPxaSX2/5Ahu2D+0/9M+7OxmV
8FeklR5EG0TbixtP4nawsQb0xRRpbxUBd/u4CLHcL6prelv/FrxXWNCrr3+WzjTBBiO3H2htCrhJ
ERhtlj6aWjuQOP433RM3ZQfA0v9nPI52MacE2c+nWbMtLCQD5fHj3lwxwbl2TRUQxLrP3iVO7YCs
/UCYMrgx7jEVYJgnn0hjA3Osg9VnqnxveYEG3V4gMoO4EUxnMxHs1MzyEMb6lbM2BQSZU7ojFfoI
6E9Y5v0IAF/caqt4kvRCEMZgm5vCosX/PfodiKbFKb9f+e94+axdKAUZonpcjK0EJCBfYrpdrtu6
3ci6KtxY0MARHj1d+kqNADyh2zJbJ4SU2CP2ROse7b6CHVQBCc+ZfaUtbTMSJd+e4FHBkE2csECd
49NPWQ2dlwPcOIRaQxFB58MkB5gmlqgMIZiChDeLAGs+Hzdj5tp6wPXn/T8r9WTDbalXuSf7Cgz2
2V4bGkc8xevSqnotgicuTl27yfy2XzNP53C02zVOttWS+5DO5IgvGo6rxInG2FgG7jzFtZEGXInY
GMMtrXP1Xp4VZUZi+VVrys/yD/wrIRSvz1B3giyFNj2hxRNZGEIkeaw9PVz4GFrk0ECPcURa+0jL
p52p72W8x7k+VNzictOzSdsljVu+4AJydYrbYBsskB7w3xsEUlzz8aEA+ILWp7ccd1jT3XWh/3H4
IwQcjaf/bhefjyh/Zo3F+cP7OEoQPLfcm22lVL/vLddSvX/obf+/Xz8dw/qMG4tiIKqAvG3IoGS5
Qz1mh6468XxLe7ThJ0B7pNVhbTDE5j3K2oCWd++ZK9EgWQ+oOffc4zKo1y9OxYFnjQDmcQIWw5hf
goVr04Uu/MYRn/5PgiEYHdPreJVwGDZTO5WJm4oi2hMV0Ddiamg0D/ZFsZJrHicSHVHhS83qeuTB
fVY0goVaQS41yipvHkSDP/3IQ6V0dh9WIxQhoJufgPz2Q2qLeY/O2tW4KN7g6vxfjEofFJ9dRqYG
/aDzGnnyKynuHnZN3VjxON/rxwqBKaRdXfhbzZzWci8fr1x+RexSENDoeLfA/Sag/C1QVjwfy4sg
iZXPWa7+UG0PY3qs/jIdJqJwFlhHztkVwc7pEAx+3dS6MsH10b4CTgqa1EVAxLjIn1wIMVMB0rQg
iWNKTD3W1AeDTciFAaVZoWqytfM+TUPwGLMu7vC9BUipnaQZTY+GtOqyL33HOUhbQLrAAwGdUA0A
t8x5BX5oKkJ7M5EB2KLo++gNCRHjdtBWm4OiNuOh1cgIMTynGGEilMaqdz+H/xEAoC8aZiB57JDM
ZD59jjgf87gJLFgTr4A4OlXceimRB6gYLWerm2ER13Di7bSAQeuiBP7s8uvVkFLGwe/+uGoOwPEX
KXFZNRsgQtqx6UsVzDRMJBkw2ylBeqEfidVFTkgKaN+fqL8B1go6iPpD7Eo2Mi5u2M5A/p2EQemj
WShCcGJldRNEyrJxaI+Drtc8NAT/MWU2yHyBrQIqLj6gm6aQRdVToTrVWx7QvL2bbhxQSbE3jJ9B
yk7GBOa2TkOi7F+Eg+bElqNrZk+Ltxp5Gki9ka8JxS35EDw4MjDSFgjFlXJjhX95iGAh62u12YdM
x11GpYI6Kscx4RZqES7yxgl3t3bu6/Eruot1RE92wtzWEIxFMepnltrsVj/sRnYH6iNwEAqKi47K
GsNZXg+qJNpvSqkFcNxZugewx8gS1abTzCKaHOGBmCrSuPZupN0XRnWEAtPkIEz/sFFK43JMG27v
m2ir8qeylkA2ljSRxQ8rjDSPkCkp52lVH5OeYHRyXiFccvt5q3LLo9xmPCG4eh54FErN6TCCsip1
X9RRdOk258RbqrMfoAbPi1fjLKZ+4hDyNOm272QTPN105lggN1Fw9u9+w3blRH2nDgWRUXWpEOhM
4FO7+UdCerJX0uwfANCRYP0HMurMR18EKnUpi4IfSWhJNRrf8Kvn77ftw0LoA7awkMhbA5qQprZ5
QBZmMX8hKpOs0DcuRE+5fEST59aEL+wL5+Eznq+5677pI+O82WKb6tWlbTct4Bs1wZpnSIQ+EyVq
xofX9zh75i6914zBRnFmJq0Yiqd9bgB6VsJfszf3yRDsr/EqAFbTdPaXaR3azdvyLsjobXutVG9Z
hqweJ5xnHXsokl7c5HKNBy2pIR23nCEO7xou2pmaDbPubDQqy5pDdNONFmrkyMLCGeUxQXOzqrhF
GrXyd1txlbbuYIkk4RcibPQ+wt3Kz1i7K+go/DWSVlDXgIq8nh124UVRP2h31AUh/fVVtFOnrLfk
93tRsLfNKIN1IYry2nv7l5aCTHqngj2VEquuvimfolNnqZMa+zLo5xiFZ0GHr/n1ewtpiH46Krov
GsA4zhUAKue8ISSXh5eUX9A+lo8rE3/zdOmCpXwNbEtF9cllVVuTyUOJyy2NFL22rfBWcO5r40Dr
IrhZunQ7HUdX7TkekGBppO/EtUw2E5lC11VCI6DiUsJbXLWbObpNZ8w/hI4/n6cToDXmUvq3Qn8I
86Sf89EqqyN2hOM0Qw9CK6wqGWxH5TOvUMNoUiYSxmnb0hzFsIs6YvGQ1+nnExCTeOHiem5nV5P2
4kDP3rapHhl0HX5/KuhzukY/4Yaad1DZrxK0Sul1ZsMV3pykW7B9fMPYpx8+Ny/HXs/fcmeVO75J
ve6VI9Hczq2NOh16wI13IbIA0Fti8uriLzHXknIC1p1JODXtEI5QeNFf+Oe0+wpgE3BAfRr1lfpm
vgPEpiIwME701FwmojrCV9wa8547uH5zIxunpifxIP0Jn/BS1GVBH1TXwtViu9zY6P3EGMXq3+5M
zLqajvav9gdsBhMKhvS24Gj38cQpZRdBdDK+udP2oy9v/M1TK9pYhubSDrol6h0XF/cW5k0xkgC0
iX4ByIf8MqeLFH5ZYVmhNessE4gI5uOUu1v3vcFK6YqOVg4HeN+/Ft+ew91um48sxfT3TQKBLnEw
rBRx3yFQ+CK5kEMzZdncj4ymUo8H/Q1ol4o169TbqT0/HiAiycVExgbSslWCCPBe/0guJKaj54Fq
HeedOxDqPMB6SyLq4dVU5z87D5x++CFPS2z6X5+YPN1lKCxcf+xOZQ1SjxW2JErMhRkaS1iVu1XW
aYl5jto05h46hlMAVcahrn+1fixkjijMFBgdl2BTuoC2p2Jbh3KIHsoQarMU7xGXT2Y9s5n4/6Yo
LiPABFHcjTpdceTl4KDtAypLLwDgv9VlnKVUNUY9ejNNWbgBJhfW/oVDwS/6a218L8NTcMV7TWOM
LuIjSehFUE6ILjxoXLKvA31KcFkQltWUn7GjcikbliUceAMJD3pYXggvxJQ5VPQSuTSeTx+tgvyo
ys94FhQ5KbVoCtuCaC9YTAL8i7uh0BMzBrijx46/ks19F4GBpHWBF9YETnLeRkepv5Q2mSHLYJAV
bB9xyUugD0FpiVvUo/U50wVXyKQ2zclHldRfmMYvP2hRJv8UgbHu6i5Zp8hOlh4RcRU/RjHx1Bun
cp0da86/dlf5Fhc+bAzYIDzh2qVjDkjI4qX0GMPHvsENiVeKHezsJcwZlXBIWMYxYjNbHxkTiXMa
Wr/e/AdHu0Z0ADUVN6bzz2xeLE4ySLHUx0CvKCluLr0ILoz3B8AAPx6sVz1dWBNKBI56eek6eG0T
9gPsSZyBMUT6qPVczvXyIyzZGUTTu1SEP5eFnjI3T4lb4MP4/+gpFmv5W8hBInlscfslEmArslqd
LUoAWhhInaGAZ43Do0tKw/0/7d7YREFBMrdzdhE4XzaYGLmXk1bbBTmaRTHQNsKvT0XQPaXKITT+
yD+s/VaqgvyHmcuv5BDhOTELmjYVX/LLTZkzlywWqr7J7ae6ft0kyd87S7d9Bcdu4BEQfsUwbLGC
4mhf12/6vnULTGn8svvndyNsybi0bf4+CmAs8ckgbKUU8D5SXTTe3N3MTmp2ZCI6jy3bS7b3JsRF
TjZGkdyePrrjtzfssC/X3b/6EnEH9uiKrqigF++saO5luZ5tPmARk8A0s7/xhwWfC8a8BWMp9APe
li3ciXLMYckgRNKT6ifGy7fRcxp7SUIBN9wbokKiH5Tq9Eo2WFMGXLmyHd+M+Pao1F+TTBPfU4UL
PSPk8at3FjKyhtZqWCsuBeIQfbNDajdtpKUOPXJNYuqISTJGcFnWdGocDBpwCgEfASFbpwvpZ/GG
Zd6XcOrAvlPlh3MoXT9szCaON7imJ/kyUYr6lowPz7g8s0eE4jpwLaymdYrIdG/3tc1sf5wtqE1/
x0Vos0PMH5+fVxiGtIeHBW+P0vNXqTrdpBX4rQhr6muQGbl6CkygeySnXtQz3j0i3AbPSVN8jUUF
SYvEMpslKG7+z4v36fPvwW7m1mXgLrFMFVr3Ea6/fndRF7s4soqcnqaCeMfHJbkQFHhVziGbbSYz
iYDxbrCaUc/xQkS06SCYwFUA0i5BDk/AmoaHNqeWJf+K2XA3NJGoqNM2+9GoAzYw9u7OoVh+NBw1
CHHURgIWgZDf6a5NYb1/khGo/NoG2CFDrcMEj7/PX2CJCwmhl51yi1vIMR1vvlGNkNunG8m0yCfY
D+1JVAnx8Hur/26oQBZTNUdcnofrboFi5gy64lAj14ZYk6MGNIpX6dboAI9k9yqdbDc7IuaAr8qO
RBARlpwavctDiubWjqNZduopQ6kyAkDsie614oA0b4Q4d2vqWl0EoLh0KZSKxPp/zWwdVwrnQOMU
qgKRqiAhxgf+dl5kh/gMbBON2xkCgRyCJDsVAADREKuGTw+Qy8Yv6T6u94HTB/ezGGa1BCD3939M
Kp4c+4LunGSBk/Cbhkpi7YuqIsLfTLQTQJQbN3vcGQ7y8yqCzT+fXapNskEfkDStDi/mOjJ3Vrcx
0u5dbP7M1PLcr1tXMgKANgwX2IrljK6wSn8rRUY8rCR+nxWS7WPVLGwF7T0Upk8di9+adCok3SwV
PEx5LnLXYmAACqDs7imWHQBzxAwoTsr9BYhqiUIJ2DuwoUtIG9Ae1AKLpEjdikG7mRpeUx57D4yT
+bEcP7VCpiGrAgHTDzFe0yApS6WYo6zrj6ncAJUL+f+ybVjCHe6DhZsOhe9BaXqerKuY0J2dRgal
FIcEY01SrLq8VYPG4GuNc6FHy14Fy0tOT6iOVlIOZI/ytw1Glo+LRINPid1CWFLA4E5zDJnmxIzg
jhM/pQ/yxeE4I7FXj3PtQDTN8f/Amgw63gOUkWY/kcutYiL8Ga3OfzdvcPnNCxF4hWeBVQnT1ezS
3ZuScxmS0YRtgWOs/pwOthdolc4qKhif6nGk/YGEND+Bo0YCXp46KKATBDWyZt4yThWaw1fJ+N4E
a3fl2VWA3FA7hr0d2Bh+M/3c/d8N8t0XV/sbn09nuap9sr15WH/0EdGQPTTB+wd/y5oOHW52WCUT
AF4OEZjVL7YWCa1QVsqRu38vwtc/GiBLvXeu0QbG79Jakuu7jvcwoEwRpiRD6HpX5Nz7GTBnmAwD
K/chENvr4Znr7G7lso0FlOryEhlnIxLrIV1jeddIXz5TKsHq3DDlA6VMaaC6pyuPQgif+QYofrWy
RWLaJkFTX/giomdUUaslvb6sCj1D6yDU9f4wDwoD3IEckzHokdw1V3KAXhpfEViioIZeaI4MoBHa
onj5KivPfjYxYCNpWnuPnycW9y0xwvAjReoMykBigshbF7eszZQY6yHJ5D8bd8QJFb9PcTyf+O4u
KOF+0zHwmhVDY7mYIkkDblt6dEqcEJhfKix1I3JcCduuictaCoAh3bf6DfjzRnw/fyAfIJWNFf+5
o+gJvw3ymeovgxCwbQL+6WACCx/k9EOzFBDuc+FvS6EF0HDM7DCfVvN0DTEFgwJZze6LWYUeKZyo
EJHblTpitxpVpPULZyaFCEnNHhHyFeM7Oel0RxsXh2RE1cVnqSMTb1RyVcZx6YlO+xqiaF960yHh
J7NBSAO9nLlD0nWNPh/UaSobSwhDfhirW481yiMuumVOKp0wUh0/Ia5mm2bU/cPUjouYlYLOvosl
bvhkg1FAG0DMF5wFquniFnRtXK2cYtgFd2ytAzMm30JecSLyF6m4tY4e8bl+hb/skUXvZ87SMevQ
g1RsJOgIaZaJ+zBjcuqMPRgx/XR+He1/YHAQ8ErljffEt2MrYfsMDhUXRAvv/+W2Earfc6jfeqce
gWXwYXNV273SJKMkKOPflQ3tRl9Il626ZFnjCbOFpJwsYMKPCkrTVezKHdyyArQDET2ZSsyG+9hH
HVKsye45woaywp/yDDN+bLn7N/2Hqpdg/Ps9Gj2motrH0eBCrNuJ2iY9I9LWin25r4p1BHFFDzTf
dW2jem7CJMWvF5wr3UAWCW4VkYtM9jxzVBXxYUG/Wbpa6j9iurxc7CS64jSPxP+JpxEIBqLlxIwo
F5YjbPu1AzfC5PkVzlTQM3uTfHmk3WFixubBJZNLQNjsapxlggm9PlEYs0gQ4ZaAX1PBN0iQfSlz
DTZi1sS2bHrsIQ5Y1IBwDmoxbqI6SbVEiubmfl+OinUsIR4/K2pxq4JwgaXtZTpLmeEjaI9jg4QG
uTRizzpkVXBVvp6XP0otCynw9A4uSHV7WHwwTd22PcwfChiK+jWSmNMKu2jtfinIfa0DrzjmSH/3
2QNiRvv2dAeMG9+tn9BPUiztgXtR3IgYMbauRD36LomwioLi1aHSdxLfTCybpDqlDk1k/spQJLVD
gVcxfrrApJQD9+AsX9/JymlWOh16qaE2ptTLznuDnLDxI3onpPsvFpDIvzbwcH5SRhmZUcIaPYEy
G6TcaK9joWrNoWI46uVknjm121HeqSc7Q20HlZ8cw+f17T8GTcM3mVsVLSyUQuZHPM9ENB5Bg3K8
B1VasE8tRU81L3jzeJc/VlDVFRPShMS4B5M7M81PDETNoPQyVEGgPB74v9ZnNC1GFzI0ekY1auwX
lQdUBtzAEvGD9MC7E86GGt51c5f4n9OI64+7I0OQDooVmATppmYhIPjyqEcvAkuZ+LkXHSBJEn4U
UnvHgjdyHLtSAT6OdHVkCtgAadbxdRHltDqL9jFfSQ2LhiCPrewhEvKzEqVuOt4LDEE8ru+sFas3
QzVIeb/zhX05TmSVzZGUi/nsCO/xLhTF0J+CC7Q09AV0a7b82DZcN0zhe/zfcwOPYlnnsltVb/Lk
om5kRTuzaqpnKR1xpq62YCtiClkb/1oV5Agtv4LQBX4DNqDGGCYVmFcb8cQnxzfkMnTqF5csEs4o
s6ZI8xLSggvPP5Pje7x1NS84rPndpHIdyPdbZSBoBWJ29/KDSge+esgn9bSsyzQW+59Nu/l+MObA
nT3A2+ZyXl4aqGBNjIRKOtONAuJ3JJjwFpa4kHxHE9csfC3Nxvm1NRT8rKM+I++KWAyf8YFygKIy
v5jSJJPRPI+jBxjhX3ARgPEkO25IIxFoFbqPw/wf8gthu7uZ6Ot0VKUx9uEeNsFP3xUYz5FeH+A4
d7XqPX6d6sRTQluloJOG0+b2R8f73U4HOc/QApQFNTGlug7KLnsPA5U1sxt/Xo5H4pHT5LXmFWle
uZSu8/MGTZa8meT/CY5pkv9MdijhVNv1OhJBharvw47DlxlZ/OF8Y1mMpQHQ7/AVTFNbrHTojxJ8
zRyugP/yg81yFMTxpIwRUTukZXHBAyPdGSbB39lZQegCZvJi+rDzhXII6fwfLPfp+w8WcQ/aZWZY
8wYh8NPrANUOaCQe5dq5q18/ma+ecmwTrh9MKgHWnl3VpS1AaClgWapfTRU3RPewFl/+sX3rc/CJ
ZdtbmcAFMjNpTWUw7CqsqFH+Ev2FpIWmpMHqqUk+JBALuYZ90quS6V7aTsdssWG7E/s7wPxpZBvz
MB9kYhUEUt61t1FKc/RcCe/4BYHsAqnXyG1LARzpH1aBfgYXzHEin8dvK3tBa610aa6ejoqx/+HV
OsFO6fBt59u8Qh79QFcihFGxHLELUIKXfTikXCPl8I4scAwaCMTUfLX6fxucMI100QMfsQZYJ6qj
hzlRMnuVbsxpScQffXA6K5I0UoonZc9Foax2VdFkvjel7ijZROg69GkMwOygrQMGmHI9788Wsbf0
34Qg8rvLlvANXWnbyp3vsQdlW8szscfhRcRY3YZ/q4yqXWOTDPpP7yAtpWr+0BtLsAnNXlE1C+Hw
H2p7GS0p6GvJ8+6L6ATmcS0kpo0QBqs2Msjt7hz/9bQQEtIc5XxBClYKa7yG2GrzfZg7jtnrsVYX
nueaxYdSZqX1y0v5zvKEwokV8e/mZt0a4p3wIC0rzaO8ztw13vv5mRGaI08z/0u8fXSr9JEJn9SJ
ssjppLPUwOx1R6n74gqZn4AecgMmMyE62ir+Kdn/xymVQkE5+sxNmYHb36uE46awM/tGPdxSl82p
CwThjkus6R5NYrIYDb6+F/a1KAvdPlfHpUmC8e90K4CoUxxpAdILfahj8wNaYPrMU731UGOffAM8
cktQ4AVdn4nHPJFTiAim4Be+Lgz6w77cVC0PGG263S4lb7eXjIEtYO3FcXIygITb7sq08egPnWMj
x+g+LIz+15Xm/bKfgrFE3/23rZ9s6IR/qim9whMTOAU3Q9+neAdElhoH4dR7gcd6iICPtDRDcs4O
nfdnBxzm36JTCtd0pLKD4VVv4IzidufOY/IiYJDDPCJqMfGMjpZA21p2+y+F5+65DNZfoYnOWS8m
pA7x2UIrbtIiegda5NkVmdhPUy2DeFk0V3JAezJHJH/A7ygsSE5s5PvNP4W34yBp5tcX4N1TFNgz
0gPeCoyh6s8LXzNIEEvZxUr5sMObzmyg6a4zAJm0rJIXyemoZVlumoPsumi5OP042QklBsWdWmNt
GlrGu3G0GPF2kXdkWtVPXt9dB2GVO2LuiuUoezHb6GgoKTv4uubWPQzC4vwgpJRxopo3Ce2oOhMv
qUoSf0pHw9gKtUGLWvxH1N0xp8yeUMsUixL1lWMIjrMOlPj8BcEHmOCRUxpAqE7K3g2cGiGG5yor
hyM0cL5uq+6TdNTmknftvXdWNegXBNKgYf9QkWj9UKxtMFjiwiEdcawPwzbeADvI6J6KorLuhuV2
7TMdffcCo8Vqzec+mOMxc5nnLhdvpRlCOBzyOPC845Iu5wiJN1qKpoUUcLu0CfHExTtuBXdyL01E
pEBwywxYxapVDNkKXfvKYqSLPkv9Dyim4WDanWzG9QsPHDkoaA+REFBHpoMkAz3P2l7UgNgvdObS
oDmkRWbtX6JNo9Nv6npmuABIYhB9zZmUF9RGo4poIpdglvUuEYKpdRaaeEuQCxGqqExbtm6nthOa
1D722ew4mRh+F1TjbNHloUhRTmiOm29zzzE2aF5DFuooEWuy2MYeGaQq2W1Pvg6NvyY1vqb3ldWV
nbPu18f/YUfkEIWXbPIrWD0Y+A1cDq4mj8S18gCC3uBLaUySVB7Zp2HmDmYwV2mYNHoEDPoK2Ahk
/4oOzwov94UqHHANmIro7nGKFBwS4mJ3xUwpGzvqnYYlu9s3pd+VZr01QBlYf02POeUZVnqKo+Sy
sTmthZfrUlLqUMW7un+BSNU6SoUuL/IBZSsR9/VFSEc8tBQCW4y38IM//UpaiJBwsyVmPEmUj2CM
CXr4OQbzI3m86FSFPkHRwNKcC4YwOQX1pA42kM44YAFyXrXLqZJHYCYohm7hsMuwC5+ddUP1NKgK
rvfjJp5QLpL84zwa/R/BBW64FlW/sI9IieM+tonaXOlZT3+z8OKYQhUQ39SbpmbvxXxXLpviN00w
03KRrEMghoGv8DRipAf0bsoZ074YGGKe2trs1dlmd44UTU6zheSWB17jRICcnue4AdwQ7uEmnQIc
8szBz/VqPKOehvYnfg/r1z8SBou7k3am/Q6lHEIAuyVGEKhQUAsjrfXhFEV4c7D4U2oeVSkL1pei
n74IUePTfO/Xkt7ez/wjl3iyv1uTgsm2QnuvFmoWfEvn/U0TeFVTrT7MewSO0Z93HvzkKMJA9E9o
Mfhtrh/ySaPPmZ2MedeKUnJaoADbW3jAs+2EgYuFNjeXD9PQ1UgsVZzjIlYO7FnUgHjETsEfJh4h
ACAiRlQrtdtU251/nvGQbZ3AqvpkuFGeLC64m0TnBt/NJhuEZ/aShDljCLjfwoxRkxi0o5pZv5AI
it3KR4UpiJ/x7pUne/pDpimTRv4NVEz9OgkBimn2DYFduSfTfIqjIRnczWl4bFk+N+6kNBj0Hc56
ylRKzF/jHfXXCbRQ8Wh+1NEdjocpIgsWm+FgTTb/sAvB8h+Bm65sZeFUcFzi3ePhKnLedrE0CdK4
XUxr4R9jmML14Ee/jwe/SSy7ytTipEFYGFHvE0tf1XPttZf4giGYFf6UX6HfTwvUUrQA4cdyaYQK
XI9wk4oyNsFmjdlKaSgokaIbZvQOn1NX1ynSL0X3bgwBUpK/GDQgLGX2F9KPCUknHH9dDUS8ERsZ
E5A/XkDCM9sgGrzauI58vK7+fp5Pvp9mewvUeUWGm5yls/u1fCBz6zjbGu5+Cp8h2vn/ssAYSSUZ
yPz2MPiql41zwDBwosbKTnIZZ/Ehm7iLI6tc1utLAn1TS6eSs06Rk7CPSSUFI6vncLAFwiSern9z
Guuo+7bF0MH4SBEdCBfY9CtSOSTPYiuD6wbE3WX9NiYWOMC0GAdASy1s9W7pVEst5anLPo+GGWvb
rHBMbYQFYncLTmVLy/YjcfbKbyvC7tO7VLyS6o0baXDoC5k1nX+qHKVlV1Qgr4/2zmxi5d5OF65r
dYGnTTkqvkRuAndH9fJYL5c4TmDlq5SZa/MTbnF4bNLSn+qUUy5l56rYEx7rfwVpcsKKuQL6b5s/
2pwVfWmUEKKzuO0duKEVJLYMqBCNw8J9A2nwen5pjd04bUfHDKfqVt1AKZajopDvh9J8p4+yFs3A
w4WkvTojmM4B06vHeakRtL7amsWnybiLYIdMkSAeuH8Lg5iGgLVSrhDbqqBNcFNWTJ7EvqBXUqqE
oV04gCw+obzFc5AvGBudA96ERBxjzMjfPEICTXUCwplUka1Jc/aGnuGPgrA+hvDpcBGyxey6c8oO
TUDdGfZ7A8Ps4EvoSAHZvUyJEFjpG4o+XYiV9XMmPpTVTrEGLrrdbbVLDhdYlJf0q/tgjqqhQsV9
3HLQxSsYHj07/vkGFfWcVYfxSgryD+b9aLPhYbhoyJebrEj1dq+RJ8SfH8Mthm5p2sLRQcKS227t
Wd8WUMML6gpKLSxP8mXN8g+442mTCPw3HsYZpkhPiFfQkGBtzFPiEIJLGxpwWhxVJE+vZqGXEodq
zYuM4OCNB99r9suoEl79IuUGPxnm6LfBtZ+RX+qFV1Q7fsKySaLtfr3mKSVlrdMRQuxwyI01vPCD
puTFH+fy8lBTggX0ThZbOqjAQp3AH1R26BMzFq2Fg663Bqk5czUpoa2qU8ZvvgoNNCPpWtbm+X/Y
8P/5w4uKlDGL89m78haSVEtWn/LawLYHcAGMUtJ17Iy75c3bSn/KOO7w9OlqzPZyScP63MYWANvb
X2YgnnJ1fyp2/3Vr/aMFMSHVTVO+9QEEg+DfSXXNzGbukmq/OUn94wWAERY7UbvjRvjlcP3zAcKW
T/XFBOANsKlqXz59xHmL3POg/24xdlagxuONz5jQr2MXLP364OcP7rYgg773EFePUAsjsLb7t2gU
IUrmumsM3BWmupWeM3g7uf9+6/XJJQGhYxpEdGiamYv8/owyxjjt7oZJqAHbGKTgXHcE3OXBXiwl
n5U7hW4yAmHR371bk9byGX8Cw3fOiori9ghmHeRI3M8RPO8cYSEKHYPh+p7eWZqJ41CZ3yBLx811
AZewkMQpjqfslKevWljH742iOm6OfPjS1NQBJq/lv1ZW0/6CtYf0nvRRHOay2xL4Kfulrrl2k/MR
29kWTa8tSWBHJcDVQISYi2jCOybhta3JLwK0isYQO0PZsZlm3KJb+8XxLNG50sDpqc5B+OgfyJfW
VeSUeDPeO02d/PzEjNffKrKup4WXEiYG4EqN7yhNG0gGDhWwHhXRWe2JpTBvQRh7w8O06mK0IlBF
u0P35f9/p3E7ORxFHbhzEiSZ25DRioihqjqo3vODIxsURCa5XBkSlUhi9D68sd0tvLb2jV+iPyL0
mbyg/gZyZXeYDJLNgwjOmHEH6EGrzkXGDiEwWQGPAn3PKJR/JvOZ9VWgxpJJmO05h4BDU6VEGL6/
IZEvOg7nvS/gUQflEOYq64K+I0x1B4GA7PkdMnOj43A6j9MVL3ouMats4s6Cm85vMcNfaoQ4g8Hc
C969sUKh+jyUxq5UgssKkmZVrZJOEpkeJ/sJTV+FX8t44Xp5STmYDdN+fYrmpNgGdHcY1ekM3V3n
94p++d8C6BpG22OPJ6UT1N2aOIUyPLSJEsWumokE///6qATTxR2MMqN4dKIlcDYEto7EcJS2DVwS
+Tq1EdLUhmRt7Ngs0itwNqmKOL5OJOcSCsmRBe/GrvD84EvERmkEf3txoHv4Kjm1QyK+cULPeFFX
qAVOVmmFcbS2Zq0FaOkQxK94x1j3+gG7vZZLtsNORNy0FWC3hmGM3PvrVl2gIlLFhK2aMLkjkDRj
UWzWTTrM9oGa8AEbdTd0lckwDp8GXxnAOM6+fmCJK2rGQjeA4ZHgzuIAji4SnhVbfFLue7nFR22k
PwnZEVxxr64ggh2xDwJSss9EFNU7+LgIJq5xG198Dn+wiH5HHVLjkkS8RhE3viH5PDZed0kEU0RO
SHTmQvjHE61RdhKMnXFveJPDOcRcEpXF8dVrqKluJHl9gY8RDG+JZC0n1EZ+uSRP5EJ+M79eSO85
ewb6ZjVdpoeVto5n0aPsSi0lHFeajp+5xJQ2o/3kz1r0R4/LL42hwu5j6RlYJMHu1pOzZRatSJ7T
C5zA2bCU44H4QT0+MmWcKcBc4IBdl4PDR3qxry0aUslVFN9u4i5xKjRpn2NwEzjl8J2PVWlYfdBK
WgohL0rF+2yUvusA0iLZJyYD2c5ADygpL7LDxiPtEf+rNbTMivy7eZUjgMN8xSXszVACyQwB0Ea2
sJoZi+dtU12GQk5SykUJRbnGiTTEtilmvdCyuky905MYlmn8wix8s3MTMwExaEwebfSHtMigefoT
M5FHe2nyJXs72ncYpph1qwH4CxTHzswl/RtsiERKVuZiHBJ+A7tXK4Wxn6qZj8JKfsW1qg5ZPqaa
9ABbzkvqAu+Y6C+FN0QllFDiY1hztHELPkiqkiqDVwDercQzrCZyGjffZN8oRwRb/h5yjWG2IpNm
dMnRqTuF2SqbFyYUQUzpqt+rJgkodOAsqf3oHe7ACKK5Q0rxwDd3JSGE68U1gETKImxqBF2w1dwB
8yIuPfAU6mxs4yeeDzBPEEkML+3K3eNCHlDezyqoZQ0CP1XBfu3vWMO1LswVBKg76G8+aGB7a9iC
ILaP6dVoTy2gDxxJ16Sbn9HgzhnP7adyi/pVh+6weuiOVkQ71pQkQxXu+Kb1jvsWuY/OCcpggAjc
vS+lOLR4ZnwW6sknCJIRXOWKsyodBD21j5sqZnFHPYxgZ4iUdZOlx0xAm66IDLW8iqbMLJkAlWRC
sdKnOb733P786JGrv6rXdbuFbNwTY6NnBofheQiEk4uXCT4r7Va6j8xOQgNX/202l+IwT5LEeC2w
V9NkN1cVfuyBjBj+7zWCPOVT2h5HB9z5tYK+4mWBb26ZbsSwNm/i08Q5NMfy2wdpGhPYXyEpy0SE
+IoFGBmWCtwnOPyKLNrPAd7T17OrEF3LvML5Paq9uejQ7xeq9jNnzVsMYEGcreJnrsFlM5+Y/W/T
pNhOaoVXImgeuYXp2RHUYaizNtmgYzREOAq23gWetS5yWhd6ySc75yT/AiUoFgggCBUmO0pIjQAV
ntpSjgE/5Ls4JElHrVhqcIGwulH/jPbPtJzMlHpSoC0Gs13Yepnz2icPubxi8va5g24rlXN++TQs
DMkcDdE3awNUFbZg9l4F4D5jZm2zzoa+nDrkR0b8knVUPoUxazHEcmqIjvLeOhOjyaGbcTz5gxjn
T7FxQ6LzIMNt/xFR8IWI27R48qmVQba/tNXuwmiabJCP547NVrRAnxi1vop36BvmSHr5ATKZmyez
pmj3hyWgEnADCHF4IMviWGTrYfVgwDHWi2eFTMjkgaJ+sJ7VyfXyVXQhXie3J7JXgPcalacdUJj+
ZG0BXRhEH+UTMr/YKG5t76NdmEfAobspDPEvZ8UWXK4uYf3BnPF0V46XMHK7Q8TmhwDbzcGb/rjU
hav5N2yDk/4FsvNDnQBTSPlIZP2lQgy9ZN9qVqgP5MTKO5FxYuGa3/dqRwFYe+s83Ah0VFqLNUCU
jnLS98u9XiHYzHO1WIb2povymXHN0a3g2GXS1OTce7BXD2McL/RncD1gW4v4Q2NuNxR72laR/wGl
xOYTMten4lPQuLyP28ksN8gMVFWLUankO/5SUi+b2bZTpNrrtGeTJHX13XAzlJKox7SUlRBLYmpm
RpqrxgtMZzk173W9ekrIdz4pEGN9l+h+w8viC2MnEpTEKuj6rW3wtgURZG8WdY/A8ad0Lx/EoPp6
89KbziZjpi8VqKOU2lRalpjFS67v84izLLZsvybc5U91OrPL/1ddekFlEdLXMoCJy/V7pd1r58uV
2ujxwEt280ESRKbjiSqgISHNbrvxrDuSKICSuhTupgI+c99Zro8sui9E1YmphGVLaBE4X3PHtcyV
9TVfBF+kCUrsVEdUatg0Htb7m7vYoLQgPBBy9XygsgnXrZzGf4oOWFr8srOJXhrAjWEPyodFFJh7
3kEx58wBb+ZqRZIOe4MFhnvYTqK0fsMdoKmhE+Iy58DM27rkEPEahGNFj9WRDAYB5oI5+q2iUAA6
TGJl21QvefmXt0CKKFx7BUL9W4Kuxl/8OCUXIQjykwqjk8Cg5YzEWghJd4JujzRY+1BpmFo64qx4
iaBkfA5fYejp8+lrE77XG2vK4wQX93L+ntyPe9/jVcsZeXmZ5CikSYIXprFBBOUGh7fVXiTnjQW6
Ne2+2ICyXSWhvwTyXR06HYAr+wGMfD90cmmB1+KyOGBrJ/Grd8Kz8Ht8SGtKpnRkEXk6zhPwIokC
jfoQg63coGQNzL6c46e5S+ufyP32Q2+7RvlcbqTRev54WV9cKwLa1fmHZdSSjbaz14oZWGLanGix
82yf0+JGXBvfz4piaQiRnPP3UxuD9TgREJG/O3/ZE3IM7TS7+SVH1l2kFBOBYPvNWANB9i43fsS4
Oh6eqoYGOHwnXI5aGuUt3ISMVGsgon6AzBSLIwjgkGzCEcQqCmJxVG9Ls9PBgBU2dCo0APQldBms
G5s7jIwLAM323ynT+ydYtDSUprcMCS7TRhZqaKUXVxMX61bX5q7DjYkbDX9+73uU4qwwfgZXCuiD
KXm0r94fJbSxwWuE5jNU6rjmVPmcV65HRPijTuwnkJcTQ9M72IXUtqvadfuhMnUG8x4E1rRJqGTR
DIUVLEggOluijvntmT43ZxwXheGvGBad0WMqSoGyWj+UM/mfy0xOL+4h9xS+Ipv5HZ9gMAlsY96O
o1Empd/hm6K7qyzIORPWxF5Is2bSBthC8eoCH1432mOkr9fEnSVDoOGchRWbnOBpHy81CnYShfI9
iB6OHnhGhI8y1YAoMjBfZ2E8X6Wloea/FRu6Q9KKmiqWEnqRhBDwnjKI469POuILaOQ/6XXZCyI+
qyTbtx7xnTmnGqNg3RulgyO6PiotkKixz5hZi6OJhlIDk0qoOzwABWuLqo9eZ/GpH/77CUzEy1AB
KkzQ0EVLnuwwDmBmhHMoKlBvL5ST+79wAAR6YerXzRLjNhclrsIK5dWilLWSHpcq3r7vEfI0eO0V
w3A0trWTzajj6MD0+OWiHo3UVtJa3//q56HZRyJz3lh52bkv91BdKVTefwBDHK9CjgTywOt8i/Ah
XkOiSaWL+BXHQJ3g2JsLUSdgk6f5WjMSmKJBmmQtb4Z0rEk7IeISE8VXqx0cIh0g6tp3tk74kRUk
ohJZK8W29or7/MUsvP6u2uT9VCVBrHQGWKNPXcTzV04nMpyKoQjLhiAfgfIXix3V5E9EFJ51s3BT
xPiLJ73eGhiC7zW+KoTlNSs4/Js09X7hiq3tQANDq7uOj/YFvUTXnLaBgamFfEnfDDANA1Hkzpa/
Bl59srLcfTBQwKhLatkG7kg30+vDGKxINFr6kOq0QgEi3JMC6FhNo/vu8FCl5GtLAIRPMBK+SA7x
JZhDNLLfZ5f1RRQi0YMTC++3yBnH6CfbH6TxcenukmiXW2YejqxPtWsIbP5dLiJRDfLGDq89UP83
+RzBs3lRl+WZTE9gK3uAh9DaW24sblu0/QgitXWTWvlQWhU+rCucenhHOYaf8u+ufIexLMWlAEXu
886eHK8zwoGTtrMGkhG5rQft81BzqIXJNyxX0BQWuM7VRTrHb3bLrO8+b//FBcbbaNex+eqkmAne
EFxb6Do1MIC83k+exl07P+UjOx9x1ePkqriblmtxVBYIFC/Mmug8MVMRTGTKb2Gcmr5W1AfXCxYK
WQWkoIbDjT8MuIpJO5uB90hB8Xm1xoJNBpJaIvxQQfpi7gwn75aDIm3E7s/+bwtO+skzay8thmQO
jz/PDNHUbrtF0MXXu8INASnl0k/ycPumNXtzwLzGJSrb31VbDqWC2o1wmvv4Qep4LoSuPTICTSp8
NcCfizGmn7soOdV1oGgnRw3Tblt5ZQnmcf+C2cZkztjkILlutto1Xd21hMy/MF7YbfY4m3NByuSp
SBAMEsOPf+JuJnmvZ+pYSmRv06k8mrZxS6D2tIoqk42hn/Oq6YRdWZxREO7U+ESCpon64BZ6IjTZ
2FcA7VWaEVJR6Gahp9nU34Sj/8Awpf/lRFIOeunZ1kcRbt3lCcMO+bg501TW0bo2fmgqBYvaLFE7
j+cKmSXP9VY4PFL/XJnQuAx+s7NXs4ijncZCdgQw18a0ho+lMiX7c305sU98qn1DCQ6/r7PeZqg+
3FmY816dNZDa4cE0gRPrjXnf9TOJiUrpdLzEpYdHVRX1f29my1cGUFzbyeUrSRtuBXdd2XWqwH5R
DCUUdjAVqkndpMUZefgLwPeSUX3oqwNy+9iT1Vjg63vr4zLDEfbn/OD4N117yioxr49xhys7QwIr
nuCGEW94GyUAemBj+g2yMojrx/gy/GE1P+YL9zIqf9QIrhT3tuO0p+Ke9B8UACBhbE5QJ2LFYw/Y
ir+pbdaIgmkr/9NnWeVag3Zka16fKtp+DvWFUbXfV7EqDnElkCz81ymWyhzMd5uXzHcO6k8Eg/Zy
j1wFcn8rJ3z8tkZkN7I6VXynD0p8UGIuGwrWua9mHTpiWVZZBaAIktpx/HAzUugH4ALk8Cpg7yYf
oV53g9IMWkDeYbd8ejNRbGNzuOhhMWzsm2+oi8PDerGscGJharigEFgRyjnxDgKlecwA8mSzhpI/
OpD+zwNxQ2uox+ux5kYwgsFDXGls+APCdndAHGVdAvQ2hPFQqLhY04HRJ2JyKFB3AWpWD0BEILP3
05SqFW64VT3k9mLKi9uHsuAca9FEAMLd5SxeH/lc2He6Vir7iCWP0B6tPKcb/czz5AWu1oJWvI/E
yTcMdaFO3F5BEH7dsru1jXPR+P3kIDNwi2fQ+7MoPvRFBxg4igtpr/yazGAHDYsc3gDBwWSsVL7R
L1tRwHr1WHjwVHKa/R5oK1f0dF41zPSHZYiYTi9fOBF7i151HLpcV18PviNIFD7LdaMJWH0mY80Q
aFmZ+ecfTIEhQxBVwat87jCm3fjxOHAVD+BO/Rm/huRT6sWLDXvLyt090q29o/dAMEGVGrY4VjVS
/JDUxg1bZ+MTo4R/RB+1O46hUEpWmldlMLAx93yY5k2UxlcR9n46Gzlvsr4R7XCWVJIVLsz9piLn
TjaGpcIwJtQDEkluFZuGL/IWe42rwyemkFH5B7tTN8sU88LtIlk6Bu7vRlo+CQsXZIBuzLDQzPZO
RY9jx24K4b9s5LzX/lMldpv4Qye9XR4yfifMX//vPqxtCiu5dCkcFhbyKcR/rSvHrNkkc2GqCix4
a00iSEzpV41Eju3e4L6Plvhc5DkXQidcvvdQE77XC8T6i1Z1ht2LztKz5tW1JYPpqnkhc8KTliaq
Ov2DkdPD6RLRzw/UXmh0aWPrzf1M9KmMQqR407x6wxRhqg4uKaKgc3lxf+iobdPhZIF15rRkoZnh
Cl8Idjk3kIfG8AZ/V/dffJ+wiw4EzKv3SsINOvjhpraw8X6uLrCeI01jBTM/IgluV9Zyh+8subJ2
NhSIomMa0y+pE/LOD4F687099H9JbhTetIVTUuYhJGVX8jUC66UvCLYop4sttNme/YCZ68VX7144
FODfl6+DAQ2zXCQZXiI8R0hX0ukhqc10IeBk9OaaNgVzjqCX/rqfTXv+6M1jbeZ5018JLcNtdv20
GI+6Bh2yDqTnDyCbsOv6vxtokd2xw/8rvKmt6d6O5mV2eSUd9av51YDh0lIZN34K/Qg2nj+Iup+i
45EM2M6itYC/AqEmTk4A8+XltEhluqCKdXnc6HoMAaLYcKkNutm1sQJGRvTJNIo2Fk0bsoGh/I8Q
JyR6H66/ybKxrQIV7fValBXnmFzZAuzfjd4mpFL4cH2DvGxQ0mhJeprmeoKFLlEkj67DHlkMoBTD
ody6vofTEqcSQDvaqzUMZospV7o0EaYxEnhTTM6wFKKzkvIEq5txkZc9Tmd0CiFJiKl9QWjE5fw0
xBUQE0PKeUIRP6NBWCVerE5oLcoSM9ES1WzbVWcpbOUBRbqrqStoU1+ixgAJpJ7liN0PTarSKJfX
loJFzlPufagbY73FO+bKxkCPgk41efdtWngCI3U6bY3oNCMqQVug9JMsSNula0JSUI3QkkUol8SN
/tk3Vv2Fb5sQWut+ZSaHQs675FmpjVCiRMvBKNpZfPtsnfLvk78jzn4zvfLNZirzehW7dF+ZUjNx
i6EuSXaK6/LiPDPZRJctOK2v3WuDaOt/EMg8if4vYjLrWoCnJaPURpGw6cLonk+FZO8pNxC1H/yj
oLTFzyIhgo8F1f4L0zXTnR5ebq7ffA3gfXpNkC32+dpV6sp7tw1jcia+73txSUsfmnbFAp+s3lAB
9Knu+Q+l2Xy7ofMgDKWAguxliQf3hD2CHOHipTkSph4DF/5ScvLHbt2fSVOmh1J8jCdK6jMbJ6l2
FAgpOpFKjfrZgAgwD52XMqJHbSnbRdhljHHOVLnDHmUCUSMkDLcjjgKtuZ1+D7NUK+BsWcO/fqaA
3t0kIVdl41wIG8fm6wCzv0XytMP72ajRsobsezjItSm28ffNl+1TrpZoHlvBwL9Z8UQ0JWHxEQ7H
E+DF2DVkXfhMoC/lpAXLKIQyOUhhxLAbCAo5u95+tSE4y3gS3lcARSNU5lO0shDn4HVPb/LKQoES
VFEOBt8Ukp5x6uRQB5zqrb5Yy1pBElS62EsxumfJ7jCDNiIJT3zqNTuwpEffFIxMsxkxERqOjZc6
CLIbUvzPvl5Ni9FEC6g1+83oaRr0dKeVkEygRi4K6AMWMamOfaBE8KWPoTH1dLVRml8KEFPuerrk
rx9UxZEvDYEhliqiJZiK1IvlLwZ2c55tTDt9tmNogA+PBZsy+aLq+z9Fd0Go+rBCI54LnRUbvV02
9KVKTBPDa3WMFpU1zjzfvS/TF2ePQyJPEERV+AiypLQWltS3AMBVEHwQ5KLAkYZcLDdZV6OkWVzY
ASF2HUBrt18d6YJtHC/uEItvLPK21Tg8GhLtXdFtimQPT3Bbm6Kmr3LEp2l1/mVSdZ1F5+5Y7kxB
OXE6xx52cEm8SmLyIgPdGDgjguJKRSEKxNKwHrdobt8zIpGoBgc5FAGtEbqkZYxuOz2DBmjbmCoe
vGPsuQ2Htqg9LQdD8NF2vMYw1wMfROdrlHBPUb/GL1ldVuMejV0+zKJCY/O2bpyy4zwTqB0xpceW
ZipxFQdksiy+Sky52pSNt61Z9q+sLAMrE95XIyUTjCIFQXfWRnzt58IBhV2ACC2UmSxUnOCk9SpC
yfinRGuqLqCq3H1vRwYZED4BEU3dGJ1QL8RJ0pnSkJtGnOeCi1I+nLJ+qPxIzR/raldQOrds+MO/
plS4sOqj/yDaMocOybkdmYDk3W/tvWxOjqGbR6QCcGklWO0I5Derkb+PngBBT1O3KLaunYKlQSly
UNXRf5EhScr8qkCH521qUWT8tGCrkQIyYyTi5IPh4j6PH806DPDkTLDinAwnKFjY552cG2LKB1p3
ctFvOH//tMdd4Xj6yZZxFoa+/dYOEIbl0vLUk64yHNqtXB0bEsKPJuQglBwyCHZrxc8CXwMWpEC4
lFlldWfVoGfuWbrtt5ySBLeTDC2TRKAEK/U/dgKhsL8ppAFcTatEhhX0qw9KS/Omi5ih3tS97LvD
q+InmbW+JAE+5WOdRwB8NRwdiwwyEdtBPS7V3a12Luscw/6UPOieLHZAT8xhcV5CCrbpqQ28fqEi
r05EGuIjddrIGzA4hE9aX+zgN8qgxpJ4mFbANfINC0IJd7h47tVVqbAeUVK5nwQHUNnYUlk82gyr
WkI8qtKnVfmDQsrJ9UfGOjaSGT13nrbVzk6bCcKLK1FeYtJFChlA0kxqluTJOntxsqDagVaLPVDv
HaQSG89ksRfNbY+bqHSTsut3NxifATzxsqihtlaTUDDyVWf76XHOdn6GTTtvNFKAvYKzZUu+MYxN
UTN8AKtwuZG1tYSKV7va979Y5Vv+c4uwhJcWGwrELVU8RU/vipw4+q8/XSkehw6RnM8hc36rIIeH
+tNIcz4pqX9nL3adc7SE6MwCCnjKBmoewp9iiu6qu8RO8fyKPNoKYYnZlxAx9APwRwM1iz5iXAP/
zyGzQ/Ns51AtQYm8zNNkuxlGblroRkjp8dIBO2Lnb3t1ZkDFKZDwl6x630hYVP2GRz1836bLGN8z
aEh5YXczhc0kRFwk9bMILSpDgZThELuF7lEbHgGgBrxBfIma9X1S72gXxqxHWuvsmlN0+Ajd2kJc
1cxx0eoBig0yp7RPUmxVzhO7qXGLZ6cHcGWxTu7BM5whJfCXjYPvx3Ow2uD3fvSpFw6LSxdzNZnI
Nrl7o8q/2uMZtt9ohXNsq1jYSuQa/GdRFcbal8q3wUNCPTnrWx88oJa+AO9UItRcZ6zxhK4yqNK/
HNsWO5T8rK/2BMmfmt60PHeKJUl5GrSEVkR3wrBCmPQ/bK1VMzgx4gUAO3Ss/bkDqXzWKY5r+SWS
3rFDWaV5B+J8w9fqDFBom7y7gyGsfb7x55686jpItNfL4Dai3QdoZJKmFpF4DiDGys2RUdaGn+CD
eM2e+5E+/6upP6FRRPuli3HMJaY/MMIPb8mqVtil76bWjJJVzOIQjdgGwd9LkDMK85t5XCInGxuH
ImZeRVOQKxoPuwklPm1eycy8Hxox5eDHH6yu8aysdMFUO9uI47ZPIM+/KCWesFQRo5tmuO/Tpxyq
puajW21KLjfqbY8BJRhD2ymuQXd0IsT3DcJ6vb2jdNjkrKMQULoFobFErG//ZOpvwVAzNB756w2J
l+RfAhRoAdibZHoVP5DTuhFzGvhuuTIy6aq/8/TE9h8zAJwhgggZktsiN6YYjgp2q75k6kHGUYAH
5F9FHzp6LibC/tqY0cPvlVrGyBrSyt29AuPrkPHZB5STE9m6gI1HZOa0lAhLZixc1pmCH6CZ/s7y
xnIYAetVBY6VTR6nI6XMfRf2a1ayGHZzCaLlHGEdjH6gPtjWjqwNN/NDoZ98Q1h9oiO6daclp7sE
0fhzoYoID4Mrv50qlmC3luSdrE1g5Knn3xNgAhq1Vjfj0WAwIh47g25Z9+jaKusLKxEKfRqYk5jt
ZdNU/QdKhbHuyXv1BCynB+cpFUi1M1h/ap2OunremPS8E+UvStpPpJlusWawALGGlloOUPTbotW9
t2sxbY3y2nUULBvFAz6bKxi3bRA6J0YGZFTGonAIApmYipWHgR8Qy11pXwpshL3peKIStL0tVFY1
yIXRNTaNZkKAKpHfi6rDqwyaTL0K4xJddIka6k4zFy7DR66u81vyHk567bV/DIVZ5BMdl9Z7WchK
tGf6f3kki/BLx9EQXsgtoABmRqRA+OFmYnEIzo1/pWC4hs/sx2Nmd6Zg3CQKqpoi2myatGYis8yd
FkvPfQX4+bgrdm/XsmD0VJqlKWA2B4EFbEsivtD+TkUY9V+7XCObKYSFeO2S3QMiXFGw/efX3EZB
CYaQNFl1B+Gm+hclf8OCOBpkbFcWdpJVpFk+h61D8WF9oWaMSOfepBjCyiDJFYbX1wPA5Ryz2VMP
1HfHQfb6B1U1vGRHmlMU5J8LfLTdGewXFqkIF4OTgJK+AoEgOu2qQJ8iTIVScOqlm0vOQiFp80kA
5HKKex1DWfD+tZjUGElKYfhrNMAMxFnGJlK8HBS2crgh6YqbfxkLCs7NQuGuullD890HbzEFkw/h
fkZnBAR5FTNngypQoN21b25gYVX9P9YXSU0hdaYz5OcffhiOSm83+3+rb3OjcAfl3sjlCZJtazfd
mUoGLX3cXADen3jXv8G0Z7d5W8kZffvoRlT4bB4egyiexDJL+oMdJMZbPPEWa3NNaUJkfmUHtW8Z
mZIt45Hjy56jfJNvBYPJrbRNDLJiK+/g2HK3QfCBlrms7IFVsPqcggU/0REck5jw0zNzCqTxEq9Q
ZGjjOKFBp9YRlqhryRpYqtAUdls4XaAyTw082iea0vYm8HcCcNYmogh0vo3G+bhPowuXTIQPOag/
V+MXk537s0cvui+HLCwREaDDgDqo72BA5N74/MSlYhP/GBZVrH0aONO/tdxq+gtKdXkU94ZnYsof
7IK88teHVF+K4mqhuvtjypbBR4XNB6kRM6smPWdTZLdAt2p0kqx4DjRZBIRSBbYSOPtBlJARBBh6
bXrvWn/Bd35vwX7urjoaPOWHrocIKK/mXbKOOBn4vgZD/CMh7t6v5iUxI1sawXZwmkdA2nljXqMa
xcSczCN1F936BeA9B11rRrayA43EKrndrgBzqV/mZztcVFYT85TkU4OgKklCPkyICt6xOs9izgi4
NeSTVAbJjbtxE4a0rGg5TbX0GdqBeKJgOPs8Ec6QldDw5aeK8fh8CwExSgu6geA+d07mwBqvwx/0
DpskhiOh7KTyfgZ3FGEjYhnQGb12wUwrQlvm5pvImNhyuwRd05gjgWj+pRpQ4HJb8/Q87CUcNd4N
EQhp12cM93ZyfpPJPaQJTo86x9LS2/d1hfji1lcCkcJP0wdhB2Ck89cqA6o84XGSLA61gW1D7z0q
ztLw9pTT/eDR1Mca9NnECUasDrVVwxZ2yBr/NCcvYRfnbsj9KrSvcv0KtS/pqqTfQ7dRb3cEG1dK
oKlkWEbUl2lf8kUYyxf7OxWDZlJPMdfy3gQSlLKKEiKBnC1KXLpVUg323blwofFHtcsWg512y35q
jzXBO+9G3YF8/5BP6L8JDFlcOhvOCoKfzuvCg4le5NTOd0IODR1ELlaY4I6sE5YwGIA5iN9t8dVG
g9sTsXiolyLCP28hEI1FBDDrbXLsX0gwbUv0MkOzDSdzK+pDLtUZOdqn2rxfNc75fOQYJXsCK+rO
O5XUs85g2LF3XSKligaU2naVReomXO6VIQaWQn0prCn34ZvkG9DGp8U7foWGqIbtuwx69anKDy+z
XWqEhTzVR+g7sAksziorQCMC2QGQN1nPd7WY1mqgHWU3QAWz3jTNdqX5R/hhSn0y4pe/QqRUFMqa
Lkl9zDs7myywTCnRDlnkE8j8uWYzr5ZKiOWDQjtzjutM8586yvMcGmGsym/6OIdkyLCHPUe+3Wye
psmWHIWvXZ8ZMay2v1U/HnZLc+TkRt1iCYJjafcY66/QfET+77oZTpLaarao3ZhFSibvmG9O0C/E
w7CuQJSGpCY24xCMMqieiFpVdYd4zA0JIVcodbSGSTdW0vmvADhgISL9pKTZaKZ4XXgp/5klf4lm
4rXgyjNV2/AssaQ+Bd3bBWSAx4J3V5YM6gLAMgdmwtRe+ILE27+ooORTYkRZDeauXDT63FQQCqtB
HBDr1KACRXy7Cvo9HZGuT9cdqqDjCcpgZfBvoGiTg9Wrs9jPWkj7eIVPyWuiBxcJ47J45tTsEzLR
tw8YAC3b8KsIMLbtoeRRqKqUYIz5TID/tm7g4CphunLMrTafApS/xyb0WS2kKcqMNywmkTuzhla+
AWeKnCMQ9VUpRFMcEjdk4IPa5o3Fu1WpcCFu+YrYMGq1+li7lRFqW6cPQ+2DcBIOoRrBkL2udx+J
DmEOtDvEHRe/lsyrKZSioOabAYbYIPpiW8yaaNE7YaThxw33cYPKzxSxlo0FMLiw+txvxMJwQL5V
W0b54ieboWZGOlpbwEOimRiAUYuOoxLVXkf400FBLLpLj4PCZjZJTAyCZdqyszKPfe3WzGsMlIri
E5dVLFN2m7OfgTFuAUxxT+fQwDpbfBgMX2ASLqnt8nBxEyOVEs4DDbDfbbvhns+QZo5vHA4b1lNv
cgOVfyEC4jR1kBrGq8hI+f89qH5n+7+u6yB1infmEylXlQaQNqyQ5xTvMVsHoji4WPA0WFFNITib
XKQvbHGvIUnF79tTNnv828m+o+suJNTb//pk/usAWa9MXx1VD4YjRbRcotuJ//Et7y+gHVbgCqP3
xDKElgdhLMLRo7ExY19TUxVM3S6w7X+N7Kz0GcsTLzbpqnjUSvbCsMvlBiqCyFN0r+g66BvkvZ0u
i60GJydNsDkqVh6SHcDuByGdNzDZWmdz4xadQOT7CeLv00pGlHemnbw3G9DdmNmThWmDMxN3LN8c
v6av93r+WFhUMxpmdUVxufZXpH5jFcCMxAdGlF4mRSvjlFqTuwZfEGDYpqpDwYZuEPZ0nTGpWCVP
5F74bDyqjyhAhJpPHzjmFsOuOV3E5K1m5OkMhbdPnVWN3/uu3M4aYP9rHBmy3CMj8sylG/Ukj6rV
1pu70rnd7IC1TmHbxp3Ypo53woxYYEcZyNXCVt1IPGWDUntRqEcX/v+Y0TDjBG+otdUWKAxo5bYw
6ec2gtkQ6zdExbEjdnaSs6zQpNCTYGu7fe8bFTFr5k4uwap4sfwQV6R1JeVnv67c3Ka7GbM+ylnL
Xt7Si4KPhxpZXJMbkX448BtQK7Grq+8E8GFuZVU42PF9fYzx5bcdAEo7QSqmugzHuUKFDfX27xnE
S+3sKyOLrLcWTO1ZcgZ49WPCrMLnQcBJWnhbsDYgeFmP+DGcEXGrMTknwzXxRZG3yYdVacex8dbs
pVhQHbM8xy9x5mRrY4CucaIZE2LdD/nzhLOZ1w7NJX3JdmxMUdHjw6HsOfkcOX8xOMI0/BU5VqQ4
5xcuuQwm47kbKkGqnNk8D0gGnEXqoerVZDRZ7wRzBtYtpLj9wArwdtt6g3yKBRGuobfi6igFCzFB
H7XPWjMyuMn99HUEibq3tLF0NBLr5hTTx8EMOwN1aefK1dTMDSZOtpQYSFA4phrgLlJM8KuVH6fQ
2AsAFV4AUWYkY9/KRfJJdy4BkJfYsFnZSLSkfIEwoRm7NxzjP4XBFpJnv3OIDsu4ymfT7VQ60EuL
sd3AmoN05EUetN6n2+yK3HEtL++SJrgX+ehmZkPym6ww+fo+BPjZywyygkSd2GnN6y+HZ9cfF6od
D/l6GmDw5SFfaStTgPK11XpRUaH78DwaFcF/zSGdh5N9UgAQBul8OF/Ln5sLSx+dPlepm39K9aIt
ucYegIliU1DwXrfO3SdOKAqAaE+J/7FL7U8+fVwFhlFOGlNp/jDuTRKBS+hoyw9JOCk4rp6p/alw
OnHajtcmAzRaKSxZ0DG7xPvz5thFS990U8rMJnHuxN4Fav0wg1nILWOZ1yEXAcwUheagSkJsnkUc
aTPcjSeUkVVJT8506CAyjlWFBZsh1DOvb1+jz5mm2Lkx+O+2dhZ9extItvVWXtKctsHxgW2xkjOW
Zw1vQmoUke6DmwIu1ZNOO44i0bSHLdO8HRjazZtHY35MA9xtK/AggkMqGwlG24z8maWCH/Q4OLW4
GsobwB2QGHWBCKizatvYaJEAUoqMZnPAZ4WjIQVtNlxHnpwz9oOUp7oD8hgq0akeidHWQs8NwTe5
Szuc3vd3jVlJjAi6h/C7ZO8jVD2gUPzCrjhX1Ivbp2VMUixHUf5R63VBF/u9oZqZm1pAu4LMdW4R
38s4nPlQP+RwRxG8opy/EsSOaBq3fjjhzlwZRsjIhqVgvHhfUcbGEOjR8J19TGUitEHb2DG+kYBK
Idt3OTip7FAXH8OwaEjrJIMrqQXGTpWi9C4n80bG5+dpFTzIeRzNSVrvDOjRYF2bTi3MPrQXTtZm
9+qRUfJKrTy629rrfgNTNbBoxZIlCQm27/H4rfzNdTVPckFr4B5R6lVOzuvAw2o7moLDCw8poU6J
oyCA7iUo4bTtnDsXK1ze6GvbZWKUPeix2DY8HuuB8mAapRDxt2SoHy6hHfQpvjRsxvJBbt/6dl9O
5ew0uEzf8vONm0FMSBE/DWUjDqV64uAgi7o5QfKw1DRxYaturBD3JMgBfXSTR3XJFdPqD8w+C1Tk
dtVGvvqG0vTChy+oGQltux6g6SUSNsfTJmIVq46Byu/gjITw41ZLDvOlzhpgmcEHmpQEfymTqF/o
yREVzeBNJgF+OKIPx0pLg4oCZgm9qiwrUApMwU8sPGUx9XkXFtFtu2NbmpiKgJ4ZhSu/yUdXPIQY
TCt4iwfw+pY3LJV4ycFEpsm8DujppdrTVClMDvflxNibjtgVSEfL/kDTIHkRnhxYO4aSOBlG94/I
6TWEnmwoyUWFsMkj/owFVPya0SWlpsH7sErCrAFIevu5laWqLUAllyF/NWRXiuEME3tNwbPf1HBK
TUFHXos2oWEhvRyIPAXZ/rAy+rEdxr7qZ/1BL7l1SOPui0kkVGODeY3f844VnnTtnE/h6/Pcq4QJ
h4EBqqrVf2I+J2FgAAk4XMRbiJ6v1BtuLW+e+J6KduUJLlt2vsQ3XbNbTsH4XWmBCUHqmA9P1cj2
z0hS4W+53ojHcoKhruGeTgKNCV/S6ruIXtrGYwjCtWFIps8Keso7fxaf75Oxl2Gh4MZFr5hBw3qQ
WHhy6SPlBdJVJRzYqhQAPEYARwMV9xfqr7q84egz4AdIU5eJFNjD2quVufzGQSKUyQBkYt/hEvZz
BpWnpHVgE1TxCItix8v+G4Cpn0H40SXyh48hintnBL34XU4Di/aAeWdeSDA6hvDbUvlajdt0/rk7
ELO3Y1zXVwhOmrqI6UrL4JHzjxN5yqi2Px79rSHs3z5fdki1iMOj9GLXk2W0osvLyaGxqm6ymCZn
XC0Th96LlmWl1NsyMWnHZKJiVPi1AmnLmKBgaiaUZ9oqpz56lxrHnrWOD5HCRuN9l78kDDiEWoDe
OuGazNsO3HZKH8ZOpn1DcPnESKYAwJgrIrRhvOg0t8V9Z23OUogbE/Xxlb8OyK2tuVALbc+jUp5n
XbaFo1FeytXFvDAbBoLhuUjDcRBXxq4iDu+Qql9ta0Pp3hi3cjPR/wXfC3fuKi7ATIZnqHgwL9kT
m42JrkfDFJLnIIlK6I3RkrLERrnV4WGA2vyazseiQd3DdJLKxRZBFBxDZDYVeJ8Evbf8gVtTaF7K
60s7K9hkH5mw6MDvKIRcps+Q4pJ01TtdA1uAq3P64TQOvDN6nEEc5v6VCMN0X87oxDtwHHacyw1Q
OYfri9TfaeSWSwBVzxpmDDmrb2vtMv8ht2aIxUDMy3WL+VNDUUoXlE8mf9n7wH7VjgK40kCFziCl
UzPXmk1kglYIezYPFMlmBochUXMpMyCr8VGLM40AaQsabw+NhmHrwUTH6T8VmEu9v+4j6WyBhhSM
cXQrBLmVqBpmeyJ/kmaerJsrgmiocLyIkSfnErpZKNaFpswthxaq53t1GLfl5utvbZO6B8t53sOp
WpOoRgi/2DUgcRw6oMo8aDHol7fLxrs/OWiyqwiY/yeP3Y431ocA2jBrJ//mJt8+a4d9lb5BUJlc
Vff0PH73AFf/KyQyk/kAfIqbHQGGXkaT/IFnCxnxWtd+IsmTjjbvuIdZCCoE7RjfYlLUp2fBmYi8
Ds77fZFX67DmqtD0CnD/An0uIEfFq/GiVRZB+u3XiAh4OjKfdS3rKUPR3gB7gQmS2fSCpeaLw6Ma
eRFcV1C4ZuMpJU9yAVSB5UVXVfNp7iD/MK3fW6IFBqfRmTXM2r7RlKj/FjJrxATEgA8Y3ZQSNkNU
E7vl4gL/KFs4La/kefOAfxbrMGnU7MdjMduNvbH8aRvkz4wsr5e5oqv/CBrmGkyyAHA2bWZEJ3YR
A50kCIWJZkrq8bz7xkIAUCp2CwXNBDQMCO/K+2YalYoBmAuJD0krTiNFLDxc+gkP4VHlBR3PvjLB
ipqgrbyVt2U81/VfRPKEeMMcm9Il2XmnQ30amd3qpWQ11V3KLNbNlAQa6VdGtaNQ/VapEhci/es3
dHiQwVhGtXJ6xB6Box6MP2C9Yxa0loYDPHMJoqoP6olmlFbEV2G5l4S3XDbI7Oypf+UtlHBItBA7
YxzQFTMcafg/++MYlJTGIrcxEQ9V/rTu4laWbcoMmVW1as868aM7ZIfgaK6EoCun6uTSTtXQIrmh
B1d59KLtFktOlsZClIV+g6DUouq667kdHMGiFPMdnIfZ1n7jKifZHpCaK7JlgoM7jvhx4qlW/Z45
gVqRh61CEACn48qyfib2CH3zOyePNuPgH/iKLIiVGh4zLfBnVusbqjM7R6/NP29CIoWofwJ0dOeh
MUawihK6ZPzouEa0b4fheS1e/6YnTDcGcb2hhdBMGw82kayg0Iy3le6jf+MbICba7KAcm7KwemMt
mAhn2Ch1iikLueeS4Ra2ePLfB+UzEiRaPpX5KBJwIschjJ7BrMKIgcHEfwpSkBWt5sJcv8RgxGtE
rEQy5XSUGZWQwUOETnrP51O7dXDM7D3tooE2ZBeJfFf5SvUruEQ/1yJbRir8fdsJ6sd2yTlLPxZD
T+vTSF2YKJwLZkui+XnbgFEFWofaA47F9Nknkknwc2uS7rwQ8h/jLu0DJczscCvjsI9w+vAoJ8E7
WTWsJUl3sutw8ULBArECQhiLh7CfG8ld02TtCJS3SDjpph2X3b0+imOimBvUQ2SIrxArjDxglCcw
C7PS/xytVo48viDj0tq4Q4rIzMtcjJVr14k/mkYH2frCo9UgjvxuRuSVXhoLwdu2kyy5sRVA7BgA
jEkOr1T+F5HNrUnZklx+7Yzh3WY7ozzcnsmmcYWptMIHuH7aYzJ/thrkG10sJiIXwf8YXwQu5Vzn
Vv+jS6oRyKJEM3r0bGm1xlAOAaEmK6T+ecUynJI4Drp+IhJESJHEiZji4qYYvhyr0G3/vhHmwDFw
NMh0q4oQWR0xxP44tV/YKfsSMW1s7b7KUdZPX2Dc68PYZzFhpp+TJQE9Lqzw9VItE7zFc+2f7qkN
m9C0/VE5+NswqOrg8qXCEemqgy1LpKYI/kBF/XIH7iw9tfZh+Jacbvzl6pM7WVUsF+9kRv0QQWD0
tu9oMQ2Uhf09Sx+jZAygBMQiqSFk7IABeu6WhvzRsyk4gEMwvVHdU4znfzqTqiTMgl1x1TSOga/S
fiKereDNID6Am3e9TnMsW+OOeYGlfgOpQ/eY3zmPRHuzT1WtjqgKF/F7d7+gE6fcfnQYtame7ZXp
G40peM8Nmjb+nlDYpvkGP8hPOsCYBh3rKg6FWRVagzuY9uNm3LFscLlCHp+7coOrd84/fTXHH1sD
4P7TjYIjz/CgLaFBNlBQEFlkUUPMFF6Z/ctfWLP51WBho4qNJ5OmsmshYGTUxtwm7p9AIiXju9TH
ft5oSB+c9kJMJ31Y2lmS8iQFZL0l4LMaib6JeNbQLkFJoLQ09ITcp68WE/dg+XHtwmh2zaFlMOGc
T3r8QdT+IQrEGSQiOkzlJuey+yYjnJIUTPfnnWC0DdT8JLpXxRv/WhO9DIeMB7RMWzbne8seDrc3
X2+uYTSYc3EKHLlhAyb7BmUhmxDwecG6YH4x3Rkiheh+ksxbh8vnLaYW82a760osyNQSRbOuXjVt
98mNn2gkgbaZkZJaTiYoG4qoQTeWp3qmcXvVSuC2bBvMUHFS+qa/JMjokACwrrytjObRTXF4iade
SXf9+GRBumoDx8ewdY4fjivnP48PBSkgaMWdjuAofK2U4uIUKmN1FCGTNwU+4Er/1eJZKhNLvzQP
NsOrlboebiH+n3uaLVoo/9PWJx71ugsnf+NGTYhMh4vSz6RoEJUwejiZqByimrU8GLwKb8CBnl0u
XWj1IdQs6wAlHQvdkSQXqBVsJjiKN5hxn+vI+9H9eNUq2hX0hYmaqoewaMWFF9Tzk5MgKvZO7PEs
63pZocsgZgHBkSlNPg6xGpUA8aAnasrg/t2qn0qwU+A74mvWvWKnNcnsTqllVDrzcAP7f/g47Ft+
4XZ8j0OnSlDIGnL1JFlpJdpjEt7sLUto0KppQ6JpfP2f654QM6IkunD6iMpKv3FdVq499v3DJ0Yj
eRzGP6mx28v+a6/wXOquQea5mwCINpPpXmrojBUK/wbp6eRYW5Kf4afK6P+lrOyeRSBD1dISN0Z2
MJ7UGvG9YCIN9Qy7sjCwYoNr5x3wmknXH81WNpa+ysNwH7O6zfwJQna5EnW1+5elluu5Q93tDLih
9IAOGvIcg93qFHdRV4rzGnMbWK9aVmPIDk1l61kWkY4xycLQEcEWLGOKXpvqUBn4+rs9qZ9mkV/y
c4jH889AZA9LamDZKTayb0mvHKg+Hpgu1if0U8pIHsMGWo+ym03Nia13I9LF53MfYBSgVQhT0Nye
RVQ0+EPztGqd3sVWYgtlXQpT2PMXK6wZAdBn6K4i2UCFjMS9nSQoFW8rDi13WJ5QdX2KvtaRJjtn
hwghSqWmpQwWDvjKJPf37Q26B7NvX/kCsA/W3q5eWM6lpS7aA4uYo+F9A25ucaeVHYYQvEqMuIOB
LWqTEjQF0rDee7IPKf/dpWOaQn7Pk4t74N83L1g35PUYOKLhtesmT/DJ5W+SsckSd/rWzDkyZUm1
Nte33vf8TCor4ZgjZNpxoj+ktqd7iRK4I31UFxvK96Jp3yotGf1l2SFm61jZ4eEhZZTSSK4y55Iy
8AYYUod0yvNH3fJ+5kR6UanazGhRPZx4FTyhDgVKbwpsmKWawL4ntbwx2YJFOw/g4jmIRURi7W9l
Jjk5Ta+WS556YmIHRsLg4CeOGP/39wXo6fxA0FDnf4bb+iO867CNGMff2rg0ry6AZq6S/bGzaery
gG24v0fDgjubnomOywA3Wu/Amys2SyltnS6LUdbUiAuyzW0u3z3X0ig4vycrlnI7vNDg92Gy2oNp
ycz/v37juXJDzCBPPYzdsTIx+XVI7/VPMwXg0fWnMlhXKYQhoUCVkgolw6LdKlqWOfECuojGqy59
Ba3L9W1/7AkdahHZDivY3SdeJ/OKAdwON1ZGV8YwAvp7rRLmDhDnVM/a1HKGIuT838KCQ8OQRBGD
z5hukO482vMB244A3IM9DVb4ulTudwuYnqVIZCDvIz+0yzCQrkvt70gZkIOsEDYAGwa5pd2G/SBQ
MFK/gTCW09i5l0GeJ0YJSWHo4JVMFl/Gza3sY8ru9UWCuk+7KH9xpGLVPGXMJD9Y3HCQ7IYykA9z
KquwuOPeYMEo/LCi5UsbwInq0N8IXyiA+SBICrZ3UiqU2scxrFgrCYs0yEObuF4GpMMQiB5J9KSm
+M7u4IjeCp67jzWawQ2M6BXWhAIxgbZHrpdxlC73vs24MKnFY0zJSILsZJNHF5c25vaDo7QD3QlJ
OPAnrLoa3yUeDRwyvRTonG8rfJt9+qRYB4m+Pg+UesAraDLXPhtQ8sumQKOVLjHuhFBsPPi2o+wB
WKZvF+PHyWAJe3GA4khp57yBNTjB16sVA1bIH3DKAiYoeRwgXA6BD418ROmvb60JOg/v8UXJVnSn
AdTekGaW8W1j7w4mAXgWHNPrk8WU8hrTn3f82eKUrYniTFtYfyZFV7mz9Fo/Zw6u7Dwjp8s3ttZ7
6b8QDmDg4VPc3a7r+tU5QoZSetkFuOoNn9gW5D8EP4l0vvHsPz6eXc/WV8Z6iqmHR4ULhstRpgi7
4UfGnjcOPa+a7Jgh1wn1NR9falPH3PYzfTErmzBXt2SDJyxAJoGr1Wb+Km3rb/2qRRfydq/G0m4a
CMELAxOFY15SeA6aCmEBKHLID4zXnn+U7FU/kJEX6eMHfy8buu1yqQm6itgZNi/K3doLqG9pmAHg
2+i1Rza964iPH/b8XcFY28952tAdyprsVfkQqYMF+CYIGH6Dbj0sC/d3vMxlCMv62IfwvbHM7nIC
4NY+64BxRHjlgnqy62gf+1U6X8d18tE/T1nTVuZHadxNBtmR0rFFIVM/+Yn5GLWSja+3iPEyYXN5
BN+TVjQEiJNAA7rWdWN7dCNPGeyB5xaLh1+e0RjaABJ2pYp7qgjyAIl60LP9PtnNb6ZfMqwsnhwn
7wAHFytBWbqDhnmpqY8zYy2bzg8aJPcgVAVFHsfNVEu9y5jqONP6ttifgulfJ5Io5MZ5QlHTkz20
Be5QhOXDb78cvTBg6J1tZZq8wpcRyGnOACw/g9ZN+HbaY0kcO3gKCwmT+R7ERzMJLgETAw/jtEPF
8OxGMS3UPvoH797Rg5bb5COkh7r/L/Ukg/OMOglkzRZrCfGlkj+tFNVZZp5ActKqSAyfN9OJVw9j
r6lvbuRmLP+c444yFH/mOupM9GspYPcF7erdRC9cJ3P+xyfSa2mEl+Pfq+xGvW7H7FJQEx2mvmBa
YaR7glNR/QuI2S+m1cepIpA/pWN9PfmiISiW90bQt8BSsj1PAdtXNFl2LJpY5IoiOK5y1Co9gLFd
zjsIhfAu6ih8/F8ImXAtZME+z9PT88+dgAU2+W1F/AInyNKWgtubY7vIvbfrdi7LANunQXMvEpNu
KMaxXJ1tmQWEayYihYzwcwb6NZAzwgcW3QRoSDydXvwKk7laf2nMKPRLkOrWTwF4lRPGIilbwwXA
wfHUYMFMMU0XRWY4aA0GgXbxSHpo1r6xP2+KUFgBns6IGqDKrGz8NMrMMQVGvtpwUXFJDqdJwdW4
65hMNUphwOATLNQpbXpZmbTlci8pW0iWRJhZlO7K3lfrycP9yG0yub93B0a9pHk0ovpWyC7Y1hBv
licEzPvFr3RmeFM4sT0tYLtuV3XKdqkw5MYGZWuYAsgISjuWXH9MmjzDw2bY7HtP04xaPw6eiIsZ
lN1EgxomZlUzmuQNrQM3VmmY815XOKOINhSfFcdGbbw2j1USSA5nJFYLlTwyrUgmSVoyi2MHBbWr
nXMPfQ1KkvGDTqsgkHv+S0FrvuqmHoHNZDFgZLqOFjMPgMRLn3CCJ5MpuA9EosLr8/C7yBBi3zJR
xeADzsM93OZ3I2CILsq4cXdihIKek1wcfRPXEo4LZIgJFvz6+AvDIE3M+jEJzpg4cbtbnh01UHJl
haN1W9LVTZR2pFg/Mas1DNE1xVWa5sEglGXhSXB5+MN0/tuq7RZFSm5o3NLec6MxK7mwYvzD0swK
xS5yq28+OzdF6I4mzwTIgND3PgLMUYDQxHa3TopcEvqBM9bSArZXeXEZ37TFmEGSXuzPl4hAP6gZ
gkIcD9pEY79T5qawYOmZ7XHXmdR5WCm90LuqijR4MevovJD4FkD71kB0sEaGlNIFZPqltXH6GW6L
NM7utMAZxnxTtPrYBLrZg8l8ESKGh1k6TqnRnibwosePO+NXe9xz1ZYkylK6MwyIkWayOrI86Z68
o10QD5wiDze3k0ikgaYapMcKBVA7K4nKWHjAka/3WC7DfXFoiy0vMdehsB1yApOfGdU7rO1btw0u
TbBhUeh2YSgFWOWXXRniBGxq2PYclxYd3biR3JtdMeZ5dSrwPC97YrRP9kkYkkAoM1R3wy3ethyY
qLnz4GoP+bQ0Y5NUb1NuxDHSVul7Qv1RDj5FmAbS6BGOtxrXX7EZQKoYVYbvAw4EgwJgKL9O0Bj/
6UQpeq3iJn5nI1MYoC5zIGfLJMkayMyRTW8J0xG8M54eDgoieqwy3bAghgsXIXiQTYONi07FG3c8
aPM328UyYgwoAz8pb1iGJOJqFkiIYTcleBRiMS/6hf7xZeNsQA8NyKuWG/bkghhoE8RO1Yijpx5V
OwjriBzeX/idU+nuiL/o8ohS5LL2piy5amnR0HspKS56nHMgqN0ioNuNTHWZifci1Vt/injz6cyo
piFh+AqQNVSFSoZjR9rhJE2sxh0+r58RelYHBqNtc8Kbv8iZOAOX/AnvBfvdrTl9EOe3PUoKF31g
JIQkyA1eDngGdAKExMYdWKpRuhCSQy/sUknihXoUjzwMDq0pKSCcMnzgYZIrJJrM+VNs7kW6hazV
a2xLTFs+LicvmHkbyvKV28C+q+NbGIs0CRChiSIERUibAZTyoO5s1XMSMXZq25KKNMMPLRWGYGxg
TY+TGRVA2v04ImJ/YucR3UqzsMTN7tw7nGWBZ06qmytbSmI/x63xAOa3vNRpT1DYw4ZS+9SfjuBY
bRZPPmJdi8e34JsQJDnLEOHvFlT487oRH8SQAG8AoceZTtr8mBqnMDKPmJNtHznM1gX9vmVMvN76
jB3srhyksW95iBUX/0cZI/fmjwiaP/CsTETDZMa60vcOtPGr1AwsSSkt+Rf8sAQZOOKeheXM5xHC
SN/1EN/fJtkPJX6xMv3q08SNqvS+W9tga46euSdHZ0EsF3S75b//H9pbIVdIAjDfiqowZthjWnKQ
6TUw4Iu8Bi7qTdCHkB1ZUuqtzHvCvFMLpdY/RuNaozGGRU5+7WmeBqvngIlGZDjOIZtWGBrq+wB+
bXRAUAYw06CBtwzsoc148G8CJcq6uF+VjpZapLXkbis3IrtsN+cxrqaSyHz/3qHGrqNvc5S8oxj1
i+U7qpkwxDHpr430LLBi/qWxQ/RNx1JtIT6HIDJ/QvUvbY5qx52uXQN84/lSlvaCfsYadMYxoZfq
91bbFG7AY8kLB9PDueGY0HtCo3gexfmZ+MwkvPYBwFB6qlCXGK1DitET84eD8KKjzGOTJZs/IHkX
kwfjJHpBvf/9XsINA803HYb934AeVSsXIdZvPZ5rEERmLuJyMVfh3UHd3jXdROW3Tl8IpVjqo1+M
0HmsGnyg2IYe2OevkhdQfHd2oMtZM2nCp/zBC1zSHEUqpn12rc64bVuzPEWQeZHKATjDYDQ4PgKx
cfi6SfGP6sWhR0M/blmqXeUtGYO4ZdjmsbBnOBsZyKVpESV4O3SX/67+r159f1WHJkWVxnuQ/XwA
O1fF45JCzfE/3eZo0jzzj3KttMdlZsM2og9vKonXAnvhWbArTEK49KafnFCdetNhBJCtTU91Hg0b
rOOUK25oneoxLNdrIGqEO66sGnvuIsER3PrdNr//xnO7yeVLLA9vTahvaMbT8ewuyRJicvQkL84v
9EYs8Ot4nhqN3Qwh6PhKhcGhv42ZsHIYAUFESJXRVnwpJAaDvKg9nvr2HtQFFMmwrXPaCfis+rGB
W6VlbIq/TFmgXz3fXBU27io6H7flngvA6dfZ/f9eaLeWhuHEf6WXzC6o2Cg9J9YUHtrjJ4mb1XwY
8QUhaWUbMzxHacB3ES2AdOQEAlXNoQmtGzMlXRFjdQuvc5XGR62H0ivMSsdhLkkAxYN3KsuvU3Xy
ZZKE3UzRN/r7DdlVr2LJGyf8TBUEbz/6npj8ZRO0DtorLTw2uCF8UtKSpFRbpJjGp7NEQVChNzKY
y+rkT3esgsoEUatCvhi8NNfm9wnfXnAeY4d1H2iy6hlm4Quzy1Su15MLdBeOb1Dr2H2oXGbQPLR0
edptzj8WKjPUAUX7HmlDt/Q0ceJ1eYdx4vPLuxHMIWO07986kJmb3s02buVPCDGabVt1/OD+7jbD
RJT6LVFgaxfi8etkHpO+K/l6jvAGlb16SUUYcSa0/lgMqmTY8o1al7352l9a6y3bSFYc0Cm+GvsP
1mqEJWb/8dMkDm217YHW8NhjxL/YwzHHZYINnokBgHcmEUH6EOz+DYwFYZYAjRMgeZrBySxEu2Kk
DKKT2HWe1GBu/DG/MFAXa7h6UKokbgm626Oo6POkQDMwJkEzcED3YiR3cVpf+GaRurSDaFjN7ych
HYOZCBC2ErjPOrwQG8hnpIIKNLsEyCD5FAOBo4RQ/BAA+Weq4FIV5sVwNJhgOpfrwwpNw0rarejt
QuYO0bIcKKQ7WA6LO/DSZYqmVplZ+h6D9eU08QQDQGbmk5CxjfQ4D5ZhRMsmyGSwYw4vJ2iAVL0P
BIfdMqwELokIT2k2l/NckAt1CG4MEVZeNtcwvw4v7EO8O+8VXrEQdNJn0lGN0EDLpySWVwblp7nK
xIxhsFaIgrueAIMzcvN8CltBi4CoJuPB9CWGErn2Nd4Au5cZRWvnzzDimaGfi8FR5ECNgc2FlSAt
i0ZTdstt+vyOLo+qk+ZV9va/5Rn4QhmbmFL+nof5nuw0JQR3OwOWMRjIfQ9qhL9WoY9RwLWAyRYG
lse6Cy2Hqw1hqM6UF7vNB/a3QdIqbW/bo6hZkjJmfA2fEJwndyUbpUhJ499fxAG0B5YTUTUq+8qe
ySkaDXR+uzkvLd8IStaF3IqcdHRB3UlLptavEyaFYlpgjCbbO4j/yrgavbkKGiaHdBVGTmZVeo7W
/UNWQ6AQGOlHYwFS56EaLbiEB5LbPjVqAPOxbnK1Isf6uusRI5H4RUjvQiBqxxPbwfmhhhHCHLqI
c5HGyDC58Sek9uhaHQ0PshFUu9iGKieBCTzRcwB+zJKGE3MDHYIwSWC+bcp3sJJZX4cq7NxTyzeX
iRvCNOpEtO8xotBm2E44dZSjUBkia36Snj2nY2AZD5UfyUHAXgSduF4FmT2iUAvZuEvG8mD4UHO/
ixxxbpiNwqMcix3pyXJOktyi7BxNVJ/cxZRBJeOqA1hdGZbMtHC9UE9OnaL/7DC1Wwkg6jBJrp2a
pDjcdpGHYw9JYcw71AjoIvZIoE6SSTYUJAHualS7kykHQRsZFg4PgIo1rZrBOAjw6LhcoGE6Og3v
ZMT/n2zdZyQGeqLHhQMIqWdzI+gmLF9uL/W9lvnv7wZXJeLYIS9BT1i8xSU7QlMekC7IR4QT7GOq
jAg/tjJfHvw8oXm2sP0VMDRk3/ZMI0Hq62vNO1yeEx9CrsSoAkdwBLDPO3YtlEwzP/tyNfMWuaOT
ePKi5rU4AvQ/2THSIcjJLMaptRw0AXc864tW58OsYJXxnSScdl8TkSvZHC1mPMBJmGVRz0I7T3wU
DWOpT8XZ/cZGie1zI6zX1SHpzXbHSZm/sI5nNisyWMzpkthIpFF8H0zhS8VG15woYOw158QXFQXf
Y9yHOdXRquLziGVXah3AVokmmN/N7kGL68pOcMrH3Z9uNna4O7MKLmrgOKcV0FmoT2gJP0H+BwKs
lL3CU8kgyeX7gkK93NkmG42J+aRVid3JIpexUWpAC9OlAKZRE4sjBWsHXZuX34904M/BNViRIswK
7IpeTSlxBbFsfEHT5RbEh4MkmG6ZM0aNGCnV4bUuHm6dLkl63Ce/aFqe8huM5gZtkynhmba+5lX8
hRF13ulUJ6dXKItrYRT+wtOn8Bb0sjpnlgoypcanQkn/iqZAEh/qxf/tivEL5xoy83r1KJtviDAv
Ae5qkgj73ATh8Adhg2e2ExUvhbKeRGgYQBcXc9ZuooGYCXD7XOS7wrKxM94+BZF0SovU2baN3EMr
+SThX+qdLpPBltlP1nN8hXsd4xiyMyg1bcDQq5PUOLDE5iyDpDgYW2341pbgnFIOmgg3dq6vjCB6
vnSjOEn/daLq6aV+RiqWv47c0GPNS/+tYi4b5m7vV+hhm3omn69ngnrfw3VX3BI9OKGkFIZSWehR
TwWDx0y94/2xt/DkOcoskt0br55v+RBjOUeDJAPPn+GgdmnnbPmlk1mdsF3r6lluaDwBD/l4D1aM
5x1QP4EDopVti/YOo+kXlK+lfCFmyQBGS1ImE8pwO7/X82X9YEv5Dj8UmlKhGOTAN0Sa1DjBZreD
8lOpvu/0Wh8Mch/ssW1STQyEQee8VMTe7Yxjm0KbWbIzSV3fq4rm3awHnsIVFUWD+UBT3+io/kP0
KE3JjkwIJQq4h/7Yu4H5OnF9crH8j7RaXj/SFoUTh7Y9bzwYHr/HzWG+ktW2c0ZkGSmgFiCYtV9m
B+7PUElzuT+e1rXy/OwOW+3xbMrmbaZTWzq0Ert/PGLoZC2FfEliTYZ+cFt3W2Ngn1FgdpT+eauB
YeAbBeZitmZ+Xy60/LeQu7T/wHgrbVIv9wYj/NcezV7ym8zTwtoyKPokTOdaL1JWhylTu/TzL2dV
GMdsZ15c7cuMaKD3N7qY9lO0/1qwjPTzUn5B3romyjPVe7WcmX//dcFENB1oLuBSVlozh7gU3Ajk
RGg9veXfSzofDZiVqyxRfAI2cJSq6xuTibYXurHn246Z6EnedYziOTlC/ewO2EvO62p2jItovpqL
yLU1gQjb2nsnLcgt0j734BywjDaelNResTQVOR/BV0B26oyk1lhhWCUFrBIcE2tb6RgQ8pP9oQqf
CauD33SXrRxmDN1MKaIU+21/LlwCrqsj5d4330BpRPJxE+rUcYU6LLDSPqRCVntfFYBNh2IBnMct
r3yk19Jdb8/grPT5z+T7Duc/KNbXR/Ib50xQpmE5kFUjMNKxLMw3J+WoKO3W5sjnxuSdM9AqOjHg
BNjzRAETL4YPb3dgHGjWyJOIlEfyjx5dJ3yhHlnGNB5geAlZ1RpElTe/wc2bD3Ursg2uc/Z9Klo5
n+S+ex4MIuleYaa/c1pZQgO82hCzYc5/xoX3ptHV7lwMz/JcUg4gMd5n8PZYBzUnunUfW2kcxF59
7OZ3a6ZUEPyye94WLi882stKLJYIuuV/ODfJ7pIQKwZ9RF+Y9XgPtlkaTqx8dC/iso1iTdeWCWDu
l3BNXLbsdq8yOBP9bto11Xrz9i0hcQMWN2qb5vtuppUzRuFe6cYvcfBSTjKR1Dh3jhgLOKy3cjF7
JxXxnlaSyhwsxxUDR2dLkZLv/cU5qSy5Pv0yE2fc4aYBKLmOgP/yzJRgsJgqYj0O0a9poloZ0fpy
DWpff74FHU+sleI0EhaOtZNvh4kM6MnYRy/slAAYk+8J1jcgmboDBLrhCyEFgQjX96Bm18sVSjb5
pTMLpOjcYbniDn6qL0Czst51knMp9/9HOJ5QT0fDlpuQPspG5/C1ba15chIxBv6DS97WC59/NKGm
Ywdy/fAoeTc2HJ4vWYggljMiVUgmoGEr+VokRD6qX8zwX6Xcd4VkRlPgHfUrmVZD8gwo5F64Sdjo
ulNtfCPzbJGSigFW/eKumOeP9WO/ff9CwGg9Tcl94R7fOJIvCU3H795uTOl0wn4n/5WoqbD0VLS4
+b7EuwKp+2QCSxrA0WxvpFYJbjqfZdeiDF9RLRkaX90RvTc/NLi6FtJUj8HWKNSjIswStYdJijeK
nY7SxROq75FJ90EsLj08TpEhr2jq0pPzCVSJZ6VNWKUFi5/Dv7HRcBrQ8EFNrMEp/HAxVTnlDhlT
LxYF/ImZf6S70AaFm23p+RGTcoQU6tgwS4WLWiVozDk1kbNEKwwI+zBQnCZMmS7oKLkLRqRK9lY5
ZiJpuwG/UIc2y+DhatqwIvyQz5i3vFrjLqhF7vYL9Ru8llVbYfSHJ8FHc42FGvDXTa57kYGgInfw
8vDKAtTGmQI8ZIY2PdC7AFGx8poSA3GFQvoJ7BoLyenPuP2wcgZCT+3pdBUOJlig6gFWnTgsx0tX
bo6E2kNjrpqRh1bLSd72Zyl0x3ApCzMczQg9avMJQ+INQlMmZlztx2KMQihLIoM4TjLX28dF4IQW
kr4e7bzmbgpLPSy2Rv7Ijcn31LyIKWaXB+GW+UNRYE1j5/KmqPJma3bhemjjYQGtOzN4aGAja5Jg
IgtQYDrX3m55nryvbKljXIN6wVq76l40t0Eh0J1yqsvbZ064MqdD638esUTkZEQwET6N6HjuWu6G
z06PUmSdbsoLaLqpHDNcsR3gF8IhlGpn9IkXsrUtDuxWKEHDFN7CIzbw7NLIqpx9EXZ34Sl5vloX
9yirOSYDiE+GDgiN5uD6nhmyNWa+G3paqaGJ0Ur/JXmqTMRybxThTNuRsxyUGDCX065s9SWmE+Kw
CR/JwxXFIU6fG2dxRsN/JM+43Y7QnBBnW5L+UdwwEdtK6+m2n04GaT+golbCTdhj1C6ayZNRDgG8
pp/QcGulq1cWVBg7uUzit+iqt1pfgawSJpfj37NG8fczRr8b7dDm2nxefb3Q5iyh00te5zP8Ks4z
UL5mL+VfvsZKv6fLRl1Ay9FsWl9QiT4YTZmMktFY7crXeU1JqT7O/ymnsyPpoyJB95+H9Pc0F4f5
GUNFaWh/Gqyvn0YFrLpAlHrx5RTRhR0DE1RGjkEJk5VRnLyXYbQZJ31LJbClGLXpZWNI/NqKic6j
zqzoqMXEGB+cY4dYKQkE51huGCpqjoia996F3EI6+MIJqFVFnAkdMBpUQ+zd62IF1qJYRHteSb8B
5GmX6vD6f+camDbqOx/tan6ZiogjsSqA60XIicxjv1p5srxeMpO6PFSCboW6pl80kfknbf47KfZF
glR7abfTi4kWy/ZFS90p8sjkgoy1mync2jLMZrZ65NrURpAp5urcTeNjKoES33xOSTY/PtSYr/ea
Jm6OmYd1gu9DNCmvWH0IEBTq8dStwllu3Mq8gqJYO644Hk6eD+5CpqQJiM2PH2AybfAKBYgYOpWM
qPQ7FCEX8uYpHo1bC1fGnoPTaQ6h9+miW/pbIcoBgHNW2P98K4OjkjG343yxgFNORPe07emEozNU
QKP5XZ3jM6heMAGSsA0o1ytUJqF1x5sWfuugldkgS/VmuhDIkOj8aLig7SGMiqPe0+ioXa6h3vSa
uuqcoQrMNM6s0VGV2L80F65YbW6agZp2zo39fdjgTauWlrSuDj2HzEPdo7CPLFgYTqJ2wdhP/Yns
o1gMaGQl0I5UqmFaLDjpKE5kcc5RP1PYzyVbZR5oT7/O909WGvGPx09eaAGZSX631HgpxIwIvZ+P
nup9bfL4oHf9paQdDku5lE9Zz0GjgWnPmxWcliL+Ai5PV1lKRDSEgcq2augWMnQRCQorAqE9Mb/e
ps61WDc5PLJ0WaOrsGFXxBWK4VCgRm3q1x4nG320ltDVWZSM7yRPeUaxlvHuvW+8bNYp5AEt2XoA
E3ULIdxfW6BdcMdNazHHoVgPs7S5bi438vPPPzjzRGNFc41puTtEyk2MLWcqHvxMw0eXFD7LBbyz
Y1Tvd04wIwcMryUcFGn1APr+C7JrsLS/RHwGQv1WzZi31KKYckahX4Pf2/L1WpQIkIVxH39B1dp4
XelSfK9uwfVGj2ko/2k/J2t+P9Yp2wIfWhZClKTK+RgWhPoSbqRSVG09IqXP5dZGW8NGBt7YlkvE
xMWryC1uC+4GTiY9qiyKkpze64ry2sdWNZepY0mh1jEl9Db5DWWhLMWWRYXWQXCG9xCDwR3mHhGM
8P4z/OELA1CGeZ039rUIWiAb+AANUH2m3iVAWQqqdFRgVQFb1AS0qub04fSbU61QlKJhm7uFA19K
b5658+E7nKoDlDr+mfZDXWMeVqpdOUBkcoWXFqsk6fh7Kl/Ys87Aljg9GCFADbbfVbOS/t+AB0oH
nMPKSdbYTpquOxbBbmU8JSzu74ZgB/PBgB1wbetz8urq2bUYaAR/tzLwE9HSMX1C1n+wWp7AEJ5/
ShDbUC5zZKDiipWFNszRiLmoE52IwPisZIOwkWVvWwjd/h5PUNxhIhFPczYRo11ToVGkpxbSu+cq
U/130wZiszvUL2KQVfPwfDEcKvlglRf9+0FCO2jHcvAeSHBjBgYupzQGw0Lnc+aJOgxIztdWXIF0
ihBhv4wd7CR21Z2ZmJUuG4+S/wf+ktrWb6o96Z/qLvyE/wbYsE8iWxlZIZ3dAdBXoVRibljCtjKU
K8/GmDP22ew9PQa1fMG51GdmEp5jY1QqPNkI0c5CHkw+GVQhlDFJXAMjUlmWlfuqQN74B0k3n7sR
GuH4WNr5b057484hA+vNiO1gYk9PTD15JXtwKYSLeXDPXZQ9Yvey35XCry2SerRMwtSOabMP7phq
zSuNf07IBCrWYyxLJgwTlevKxbCluukjmL3xM0S4p97ylkSAb7X/HzH3kXWgVOQW729Ko+jfgrd3
q4jSbclkcFbTXzOfcRy/K3PXlq8S/i09AL06/Q+MfUcTxxiISeDRzT0jkQwKGrlojD/qTT7kmU3R
3lHqkxJaMrcFK4OQxP3VYTM27B5jB+FskvkirXQjKyJlHvHoUQ1jXvq4snVRPivKMSohoinD7tL5
De2oKuFHycxMtUAIm1/RA7KSv3X0cqj31D8h/QIejEZ1zRW3v9AgDs0te+W/QJZtV+XIH+N3qwjz
TwFrn4cVoRKa4cau7a0aBcH2ugCYypakD4a87yTUWr78HBUB1o3SOas0LzLnqwBJRh/kw67uoeXH
teydSR85xemAL70jaYxAbCQg9hq3r/8pIa6Zl27zUe7tY4Jpe3UsCp5inGVcX0QfVTj9ZnBAoHLa
kdZ8T+wHMbEss5fbsMw2tgtLjE4oaYMjpnpQOkCi64IlkEPxswSpG/swuiJ64SeKS7QsaTe4ZUxJ
1xyVPwbVRWR6DStFsp0+Xc+JubBeKm4BYH6Zth0JBWDZvhWi6YU6G/ZGHyZGnoaj2Q397okfhImr
LtYPkhvvSIhPNf2HcH8RieQC/2aRXDWMmZQ5OV+LWIhux4QR7QtLOYRnCV2auM73NESNvTplJ8F/
8Ul0y6rU6c16PYumoC7vFCiu6wouVXLvn0DKJnKdStmM71I9IYK1nKVpT1Wj4FG+498DaaDUc33W
Barpky+R90ipfyjGzA7rbx1wNKHss/xic6/kB2a3ler4BwJ2P3vlWajEemugV17Qzh89+x7lc64c
xTr4NavOQkR18KVFtz+EBpSJ9yGdI3kixy324n8eiNc35ZQLL1hi5j5tNhjwu9ty8OMGByk/KcCu
xpPzHigDDTgNH7WFW5xOpDCny01b63EO4KDXPt1Mmlrgzk8CpqS+SoPYviT3ngaEJTZFl5nL1IDs
LSzwxiK3pMUBD78LnQOBSvkDezCACS4xWjOcx41kuA4Nu0P6l83Rt22S81FkY1QSx7JAOTSPwKQg
HShRFML1RKAYCoyYJ6YHT53JD3QY72/iyRTDSId9C235XG8BS+1d8ow93TcuUaqAhXPxbEJYDrOG
G3vHsBL03ZEfwytoRDIzXHKDbpkh83cKtoYJ/0XeZrZGIMAQyZ9eBCMiT/wAoNQuQQ5TTosptiI/
RN8Xgxmvzf6GR+SScvd4jP8PCVyJDHTcNBozzkG3RLw3aVrOCbTeJmxEOk5spCbi35XuEuQZraM6
ErjWgsxpk7zANWh6591NkHfXqA0o7idx5SI7jbDGFLehg5QaEd/wyNqBwwO18kN7rgrGIVYfJuhz
Z8QkXxyIJYp0BgHizNqwKl7MbvLAaawCvsf6QpZo5m7+YC1jJb1ySq1ROiSUKOpdR/jvSu3w1piN
G1U23M/OM1CuRKTwR1IzENd4ktOFRA0sA4J008f+q+avbthKbYcCVzcKBIZM14WhdM99J4EXmv4F
uquOmhEsmDGI+40PGZ5m5+ObYbfvPhgDgAb9w4L1u9PHbIxqLmCAldiYfj4pmr9d67b8cffw1ijD
T/278jP9JZsjCMNWK95h4Bj3moMy+5ZA/71cDddf5wfaOXcXPjRjgdxOSQ7DRxAo0O2e4u4TkQmr
BMI/ZuoTa6X7j+HvOVzHhkJM8w8RVyVlaQo8v2jrgwJapBOVeHQzAOUjaTj9xHy3VHvAqCiMzMXZ
pXlS7J5zKJrXRjQme6El8zYrW8syTSfvANwSm1f6Ln4kflgmYvg7b6Fxn+4pA5+Rlq6rQAcUF4Hp
Bw0yYsV7mu37MPcmHM3xP7KYBHzDz7V3R5rB+EEfJ5FAwGSVowqMsZx78zAltveVWnh+FyYNUxgB
mywJ7JEhSSXzHtjwsgBm7f73H8STqwoMcIi8t+yiS67xOgqe2Pm58Pzc94nyAolVkv7RIsr1xi2b
WRYfu4my0YKU+9dMK/qK1nQS/sjgwyVvUVKJhmce3pKvnUVBXZdgVe8DM1kk4h4HTQ0ox29Ngprc
u/FaRXqD4qov058DDsEF4C4xaa5fT7ZYXEaXP5SQaTsG+kj24U4Ou01qwXySBAanOz+Rv2HoSaAX
DIo83C/2VPOEdps84JYg65JFzEnnyqP0+ihhRdd/Pk2SqcQYPrXepEDkrSj8O91/+1OFEZzUaFh3
VzJBihOAxy2UaZZDqnSuKMY5qk8rc1d3j6Wu4yqokFBG3pMNoxPRO2GxpWjVu8pYJP+Vz2ywBd7P
e1DviYdCpS0mwqdo5kHBPZvb6TebILswkXTS6ateBmQlmi6u0gZMr+p+1mncjiii3ed5PioFiYFT
tL7gtRwOL6eV6GVFSzzbOl1eJQcI0BGjl+qF0OIzlCnIw2YxiuYTBFZlu5+GjlvvWWJxYXp9EPMS
OH5oUXR5iGDt5VDKxNxKmnE3/tfp2SDaWa9lJhioW+wog7CqsHKeznwT0fGJzIG8WWfbgXR0iv8K
MsjvNi3N2ncNAF/m0tuVebgRlJyQOZvNJu673eeXqB8D2SGfWi6fni4kBR3yOYdAY/uhjgWYYWLe
M2Xa//Gcfa71Ltd5VzqivmKm3ntg+HQypTzTieqvbda5nx5dpYP9qsPb2D3G7sMpzm1+Exn7VNXO
A+b4+dKvk6bFY9Sxp3Lni1iWaNVfPUGOGm7dDFCP9AD5AudkIOiy5IzlR8Lr00OUsDWsmt18OO54
gZ9rfnx/gPM930fPhNbFh+n11xn4zWL3lyg7X/UIE21+Tp4MJRjD8FxjKk8Fi/yI9XI85yeLKOpO
OgEbqr+eh1Q7Pk3U+lMlSAjlNT+4Pzc5Ian1211g8wj+Z7FTPCvjFIcAL5E0/ZhOeaoURgatkq2D
JbwGUwr+EagDyu6VWQY9zxqbzsiL/H1ZPxbB/oE6ipgULni+TkykjYERaW+RTGThooPdOK5cdxNq
45iz/gSbvJ8s9KJNTEXnuty0bBy3P8S7AECOjr1bteynPrTNdp8T2DpzhOjCy5qt6o0uAW1/cgg6
Q3DPYJ+OZiVyvdUSZVwO/a/SU6XesQ9aTZIn2yPuik8P0jBtSDy19C5wdDzEibRPjzzhYmhluH1S
ZxdzX6jdEBF4j0DW/7zfUTMrVwQY2Su2+f9psPJwCO7uw8Dgw9lpJopqMuy7LRoStAl2hVxMOqQJ
yNQ8ozNAyN2lSPYXzLxjUU8v9UnUUkmnGDXP3VytATcYLFUaoBwaOlbfJvV94jWZk5bwxon2ZmCL
lm/ITMNY+2AovCMTqwq7THOtGQK5AU6raWnVe/XrWx9YwTJx2Uy9NPyhue8fRMuMX+6Bxv8EglLu
+m8crr8PFRS2NcGyfeeskbMgU9GR3lImJtxjk2hGf+6Quobh5Q8bfq8peohi+LV3u64mcOfxXsiN
vPgBBXfjvjQgBOm0iIsdT3TBXrEawI6d8S1XwBoRDIr5K64+/uMQuN+34H64WOf46t3XU/jJATd/
pCsJkrZsweLQsGXOuLZHhFEeMosaz8Xum5zpiXTLHSU3Pz4MgvXWQxmYQ/64ErXmYH8jT1qsh5hD
TGMDlFCSulpL0F1QdxhEUU/Vqr+FIrkdiwa9bTbuTmOhgmg6DE1dcILqt46EtYUNKX50AiPsN0sq
8ykmxGIV8YaVyfYp5CzGx9okZ7ZGaXAzMcZZ3uLk46g5RQkT20gq133hyDG4furx0dmCKsM99wBQ
0c7T5iF+sigXkSYlEQU0C/CQvg4x493rhfGFzOsIMi1JLk5QACE+cihTdN7T4pefMoVDtvqXPtYx
bRgb8oO94Ha/HwuoHbhmBkqSl/voiexDM+bYweChPA2AlzS4tvoT+EiYOQiRsf12i8iU1HbDdsut
qpnDYHdJuArcrxjQGIVaait8nwc3g8psVSpZcbEjf6Swu56qiROgiDbHTkU8PhXehGoSEhvWmG1C
s34xMZ3V2h22K+mevOCz6IMnfjVFObMptGR3ChmOCKSK5hoDXdxVacIDKuAdw78zyOt/mu9FrHI/
E3ZzSl/dtCcJvgI2ZAjVQhK0eqdChT32nEruq042DCzFPePJxflREdTiow4X5XHymhkgWxCN90Dg
nIx8lIPA/MSDaJxMTSP+wPRn9F+Hc1b/luBCiB6+tXht4pauG6sHY69j2Oqarb1zEWyW4AB3oxKy
yin44bSgtLsMd1uThPPnQ+jqr2ubkfDUt4dSlCAS6oAtdG9aOahOgiSpimscAOkPz1zfkjSRZp3b
xtLn/e/iV7EO0xSdp5ENOuUwX4ssu/ndhGx8FkeaOPH7SJbbMy2f2K1eKuNbxr0lbK9zFKKPLF/X
4UrxxaMLWGUIpEGPZHw1rd+GQEP1FSH4ZxZZ8f6ybNS7guqNDJCJTu64LFBWBD3MfG/Nl121P6pA
wLoJjAIXvyXhlSbfTp4vFvuiAo+Mos9+q1zq4Gloixt89iNVaORSIkQpRmFkxcd7+FOuxWzrVt6k
5NVMGjtOjvDsDKu4zpZdjEr3NMD0ugNe7gD4NE1i3TrM4dYc1EyYeP+5kXxpGs3NaFEUbrvvGQ4B
0lBP0s238hQfVqaJ6Evs2KPyWnl2jRx+V35MC7mP2w3BStyyTKHOjzivwIEZxdZXWlUIY/+G0j2l
gFVks6Zkdr3hTvPftLjnVCmh72nEyF09lWItRSf9mv9Fp+SqF8pseq+Jf4DFYkuy2LrvWlQjkleE
ICGmGZxuyIL+aWsl1f7iZd74krV4cTC1t4nMqUasKCicGtG+0PVu68u8DM2/DSO5OREo4kHFCH1p
63CptmhfTcoWqMDNL/12dKv6uNHHxUma+WA1uYF4sh16n1pc88pVjeCYGr4k04TV8bpBSjoVxeMg
TAJj0RrOeYDiYE8GMe+AjW+l8YjuIrvJNWyyGGj/zEJVljutHZeNwe6lkoJLbTsnnVHs/AzTb37L
IyHt19XOnMEdl4TSNh48lAT7WfZQ9oiAbY8AyS0deOZFPPIOjkEd3aXBBJe+mOLhL/p+wM7ssBUW
NhPn/YE8o6Ar8mZE4/R12angFEvzXjIo5suoKVJwwixFARpiLe+5SAm3ndYD6fMVRf/W6qFaaT+G
eELYBPKn0fKfU9rEL91ikPAkkePZMSSCeCfUTJLIZrC2BF6N01wiZifBDYH7QHz7xymgTrdVRk9d
z8/fSCW9Rq85jMdQfbH9FL7n7xT90AQII1qSML1F8G9UYij2t3sNwNq3eaUilnFcOyMx7bn7Z049
FzAQ71bXx4r/qFWSyl0ayx13KzzQv5bKNa5AeXCj3uwwC8QGFh67xWy/fs1CDYbEYM89om5D6fm8
RtnQ3Bl0t07bk+lEEZ8/wQ8rKpmHAWRS21CFwXbwHJMVBOMvzbWADqQOp05Wx/CCI/bf3RPes9YA
/CaOBBk0VqFBLPP+rJjN/2q+XPdfl2gJ8zcrckXmoSnFzjJQ+WX2zThb1hmi+VST8uzrqaBr1sUl
SLNqf5K7M0ShxIPmPC6t6K6OTA0uEqHK3SNFN/ZiPom8vgl02zPJt4KJBMYcZRpZgKkh3hiGluFy
vPSAZfVCP2OlwHUJ0QOM4xpVHsyjZl/HMCSopzgTcVTcy3PUW614sLpNSffIY4i2SmlFC0+BZYZm
/aqZQTZzQZBsUqZBsu+OBdiAJil4hhXNDkQUw244i2sAP7y7SgNDc181WFfCXnVb3LeWtvBEjwyE
UjgTizfZy+dHMf5DFIRNf5mDQU42YMn1UOSbw7ZjsF9oFlPw7n9ARTiy69Xs7l8VR6IQzc3zc8z7
/QZ8JjK6FyV4GCh1SrBjnedxhWG2kzus0NNEYR4tBV6wijjkx7WixMfLGM9anLpoJEBIGGK1qL6i
vRJer6Aq++2Q/JZ2bbyycmPH++SE0M3JbT4FEtYZhBBUgboY4XtuYQs1/NeAyg7fDUiIwq/o098f
LLlQIC4PKv3/bKDIti8iFlVh7QLwUxDJeQgE6yB6djX7Xc6jx8JIA20mrLDMt1ukqouKpdbjCN77
5gWXkb1Y4xAKqHfWtW+pkmEJxR8ffAe6EDWTRz+3ppi30zcKeyxhbAY5XCUB3p52D1E3EAzSqOO6
mJbrb6OEgFsNFceBuybfG8plG+xav+fUwjr2ItExsdNJsA5PumeL2GJWLFC4qUUZYWRL/ta6kLqr
6k5LJ6VNdIdqJzr6foJLT7mXoSQYjRhR2tUOupvy+apjVAn3HVlAvLZMLijsVw51abgrukDqMegk
0XezN+dK69cX0YLGVuX2SzExIzOGNdN3TQHygU6DZpFExpduezMZqZoC3WQAvZczuRPsmWTN0Dk2
26emAqiJwiO99JbFtjI1I3wtyJF8BGdkVjo3os7krumW5u9MoAW5JlSXoOEz3+WmHIZ28+H6dzwp
1pAHzQbzq+fYKOTi7i2aSQ3PtCXg6T/hYQdXxapB713dbym82qhNySgjc0adGA232VlSj0JSkJuF
n89JSvKSNzP6YjbxdeEVrYwXat7vEMD+7RB0w/0kTa2wKB5eHNdiFu2psERqFlWRX3en8kTZ9UI8
dGCI6RFhvNKU15sLMFUAZwn8BMScQIH3J4XAgYuA8JqnNkoElWDRs1tC0jtkav+fndwkrw5Ge3uu
RwmwcJMt7T1J6Ab9RGcTHMgqceVB0Zq95Jpozu3QMs8CiuAPTvZncsg1CQJmKiwzeu4HVUyvkbY8
2obTwQbvucfyxKrHiFAg9nX+1aAbTKWelfYIU3Mr4QLL1a89xDVQ2S400G62v6g3NbW/GIhrlTpx
zVBMiPyb8fDtaG7XgvHQiiVjb8+otdKkP5XRN2yfvaepP8MsjCSjVIhJdZ/LZrWAHsF5fF1pGJMO
33NK/C5YZa9GFM+LqNcvBcDG+AokDb59d4Ru+lVXoXLwUN/d5qFmYjKbW4ixeofMbDxvFmMjp9Rd
RZy8kYd7tclIaugijj2Bg1Iy2wmfVliBf+oXb2GHgWaYCbcRzE6M0YFl7g0yv3QWae2JbulrCm5c
S/eAIkwQQfT0o/o6h0wwB2FI2CcwR/6PA1J+FzgvIGrcolRywUYj9HFiP1kxfRUO+TMmEICwBkuk
lT/YyAYVA1Y1wNC8LKBaooC/aiy5jgi4A9PYcEfYH6MgtOYfWdJ7CLh7XFJZpBtRARqkJtknjoQY
ENLr7CL7+AE79cXnlltVXaxU3uG0JkNXc7qMiLHbmuThERzhqRc8NwnZQt3EdRq6LL+tvt4BR4dz
IBjivq0YiS05I3FjQBNnQm+cakOZ7co11qlH1BkACOKbQJKFbRmFYpcvqBUwJ6idY3jGeqZiHwJv
DNhqJR3K3ixqf6ntEyCs73tv27vyPQnVT5i0d8rpPDjZgNiptGIobg0d2sFa11Rd0BNZgLlnJ9zl
ohm3/4LiN6DdSlS+IV8Q+IMwBxZ/MPL/+TUjyoS0iip12KIERLivKnEUYWopr0DC+gXJ0MaD7JEQ
34RpWm7bUmgBPUUelxfoisxQFLiU8+Y0q7sXwZ7o6RgOH1ZvhXN5s3umvLr2AGupITxVkNykffr9
9XaNpOtep4SxNPbecWjmu1vUFhra6onP5srCfe2z3LcUl1EqYOrEeWO9B0X056h+9OCz7ZGW3jO7
c8KKZAHDmI5U6mNA2+DYY1JH24VLcSScj0zqbF2TTN0friCBJcj5JLsxdkR963EB5pMAcH0vtxJ5
ndWSNoN+LAkgCAtt6v/WcLEYr/yY7GMJeGf9KwCG5PSX2V05XmDf/iiFL1/AXdQYWJa/ILSLRhiX
V+X7YhL/mNAd1LimvkLDa5XyQEEsO6WGKgpv9lpWvKeubFZUk24qvCfpjtzO96Abkv4FJzNdxuDu
Mef9XP1P8dBCZX7VHI3im89hszj8gLDf2jzDBlZmLBrFWcbRoTm7rCJkV3v3Y2INLUsIXueagAzV
uXzlXt20N7bn9j4dWsdwG4TJR2XV95oDxfGDTNW/fSF6UwBZtdt1wnHiqTFEgtKZcnCQARR/lCcN
TcrHTt7vgKDe2xppAxITe3dBezAjvyeAO0+0cZzVeNC9Y/yAlUQSkKDyEa2BtgYYljoWQ/b1yWAR
i07bVrHpuVDf8CLZMmn8RbhfMEA83mYUr9Wc0n/XOMbdWYv4FHBojFWJ6IpnrKuVyxP6VrJNI6xQ
Nbjbe+ElW7zvAqF3CnDsJahbGGqAkp0sUxe0BFTBqFzbvd+6F1LgIiHNvgIwMf3uPD9KcAjFESi2
KHKOUkCU1xAocqDvxCKpBTOv5ANpaDAkW38yeF/Cmy2gHW8hDM8je5ZTDaQA0j8YBvNVaXrRE9Yj
gtVg4hUAbCWSXE8LijWkZc4+2uyQYFeyXQvlEXD+4NHqrpOgVO40o4FcPlQwb0fB/0tBo2lNMUg/
jhhlbmnD1kbkTZOtiT3rOgzBs44KzHEE1OpO5CZ9jf8R0v4aIfLF9okfh/tgwvrG4LYyb2JMALVc
9YluesYx2LQ0FbLk0AuM/b5i7mtRrr1sAr6bKSWSUuL93g87IMeW59hnES9MnPCG1C7GbBqU3/TC
I67XAo8JEzafTYliaPGcCpJqjBNspsiD12/Lyxf0ShoUrX16DkRoXC1rpacpQ9NVrRW1OGA0zKoz
LNjJv9JqLZhKXQSUHvL1ZcoEpRMrxLyuYR8RNBUp14C+VykvqXloncYASc8SfSgkv9Jtjyl/JcK9
z3S7ZMxBya9OIOD67119zxBpc90o+noF+qtof8YbILSH/K4NHE4xS8JgIiRh5QMJHwZE3FcEudyy
Kb701Sy+Ln5xzshfzA4o3ZXoVQw3wHr6GOuIdx3IWpsshmrNj7sajb5NxJyfHIHPaLlxS6xXbnTe
WDv5KFU+3RbyLjsem7rkvZC7md673za+Vnx5zufReTjpFVdDUbbJSeJX1umNJlFYouKQYs/1dfF6
S3QRfakdEEEWDSZREp3prGEQQGqLlylGKaa44df0fH+ZvrEd5kSa8IY/9t8hZTzLgc4qSHBrL6g+
uxWvWgZGn1nhPpMZzmGJLYurL+hAlK4qK/LZ5DyFv0phGXCkowtjd1+BhVRb5aF+hC/vOyGGrywn
wr7dfzr6Q2xkYuvrrxKRwDKg0LPadL7enpuuPND2ZmBEz+Kpk9n0qlhnc4HHy450eHKYGZPB84mv
j0pgnyT/ptE4Y/kn1rH7t7/3flmMe4SqJM05RbVfLtJBzHxFSlIIUhNHUGJ17FKOVgTAGOz+WOgS
wCSBPjXmVR85cAwBjTEvjTLpDyxTHBXMTZBFLwQhJATxoUD9EIp1gHmoGFyVlxe4k/X2+ZVpfKdc
avakvIBfwISLHvyg4x8WejykDATiSJoiRihkNlAUSD95WU6gVP+oW/g3GKyKCB1L19XjI2yBZAif
eUF6tzo5vO8D+q8/5FdbixSOR3s97YxsxG+8Yny2vsw984Z3Io1pBvsqNZYrmWdjz95iZkQO7kim
fHb/Gj6rWNR+NuNdouE3vRrKeBKWo88ycj3fhmCgigjkd4E25SMG40xHB6tPt20XdrWa4yBeTcwl
5AgQN0lBv9zl4pmTTEQl0JGvGwdrA8/mWMjwHZybh3nxwVaxMnlIeQekjb0emCGcJfZsHwqf5t0N
qHXMvLwqmQb0ok2GEeSjlurvJZIMM82DFx2jZeg35LDz6O9w/9iaKBj5OEFSMinxki9IgYoPX52s
PcpoQ0ZdJMtXkr2hQNqy26U/sart7vHWIjlLvBP20c+AzK6/S4mMwHDIw2KNgCaZXjkPSMTlYJqv
2TYFE3U/OT0Gr++gAQlZMfNYSJKq7krNQhdDdleViQ6Bm+4bHFKx8NZS2rm2zbCbsbBgJh6sXWjL
JXWYNEF88hXE70SSQg3KlNb+gVygzfFWzDavHGYgGLeo3uGvRvLnQl+NmfOGwO0WPxAh3RIAf+DT
zLfpxhKiqE+hIcyoM5qgdK3oRkljfF9pwEk5uqVL4MhojAM9akTOKXzTuyM/XqmVOH1GAc7U3m0l
BkdZfrhMNEYuxmHqEnIrUBZfF5z8vXtJ2B35g+P3hfSYsVxpMuJvvEXZDbiSmRr73RlT+UXk7kA/
80OFBuVUzEyFK5ISgONrnAxZAb+DlcuxcTlug4/4K2Mg9Kkp0ryzInNe0r/9CMmd2ZBih3wEJVqU
kklFPW47bnleFPi8AKoL8TZ+EVBEa2jegA0IlEn1ieljP8QBEqk6hXR3v84+8qtbhTytb292NvP9
hhxHnys7vPj+9Lhxi0bOGtlHwk1u8kFvBWOv2m83m/OV8ynWHBfqWBdxZrJPFG6GXbdRM6PsZxdJ
lgLSKnyZlGK8cojmvwhWkTq/Uo+X+2oGdcJzz8SQ5Q62xpOkPltxII+kI48tmwx+tBnVFUXULVHU
nVFCqVMTIXcG49+GLqyD6hvPsmjb/8WukWfTxVqR5JVOwpWexTTyIAaLPm8jdSvZUt4PER5Pu8Wr
aBAClwjEk/mzWDbJ5qLBTUAqjcqA/iRN/aHFVRR9a92bEMASGoRWfbGxFoRzdiRxUdNCw9l0gm+Z
Hf9xIrfMq63Io+RoTAj5ASvPn2A1/lUnQhJjbRgSUAFoJhVLQvQnib+EnPCH5tdeG61SNel10qQa
a/EIK8phEoHV9VA9U3RS0+kU+fH6+3nheW+Tk7P88ocY9KXUiNUHAEYRaeJDP9kY2+EEdbbYn3I+
TBb9omLXJBOdkBmH69Op58JMWsYorNbKZcxC6H997xDygEjrbu3Jqm3Rd/+TAuze+yjdag5FVrU5
pW4nRvLq9ATFM9qt2+TEXDkbaSmlzcnSXiLzdxM/2ExH+doWV03chpoD7cb7NhXCgR1BpYomYmwR
HjkR0mvX4WqRMYytu/bplKUbbxKyrYxgvASMnRt3Ibm2RxCMB94bxJwa3m/IDQY8R33KMKJZ8wR+
0T6wK1vQr+I6PAsyMYuqDRqdF4xd2r29g9iC0ronmAvAoW+M4VydtAFnJcPXhsQ6DKJy04ZXCr0I
GPafiAwfq6i+0kKVy0fzssxQEszhhTlzxWumiB1npil8MHglg+l9+QWpnG8nzMC65b0OdIV/ytyB
PFAgEGuO+O1O97a4BjC/S6aly8iKz/3EsIFp0eAVT0m51fxbeO49SpQ4F669+HgrbabNWMqN2r9U
CgIvidE4jgcBn877/cDHyKjx5D9aMUEJ1+g5a0yFJLqZO7h6NrXu+xJ57zqteynKfDmGfBVn+/pC
RjFKFqs58l7hzQp/n0qroGywlPZ0Ch4mZ/PZ6wedtfE5wUkcifnaLUAmA7tqOQlTq4teqhqMwrID
Vn8QgrQF3ml1/SZZbvCrmOK1tUFgkhkHh6ykQtS0L9iyGHlvc+AaLyo+zHojrhnVsDvtWU5vfcEn
ctWl4PB5Mw1m74CGRxOeVJJrd8V4cjbfrGQ6/sTGFNJ5RRvL3jDKRjlLd8d736Lj+c6vP0BlCRkY
y0nB3NDCYoe4Qzh73uhoWsEzveIzL3tWi0tQ/LmMUfIr9NBokIi866++rSntFT/JVkX/ukAKiPv/
dhuEZo/PcUFoqqM2akxNdh8htY3dVhuE2RFo9FMuLrpTx7EEO/NaOPmqC3+Vr0y5C/d0WzIsnbke
JEs5LE0HkbUPDAaUcT7/FNiHBU7gtNra4ajq8ZtHC6xq+xNR3NhJPDKiHiTS8HsWZZBPiehw68KK
GXsHxKo5JM/7R/FrSJ2jcpHXm5/P33R2hD6mAY09tSjw4gB7XqYwVQM1gJQacU7f+Vw42XuP5I/u
pc8BKlp/ww82p5qEnUK7v8+Xs+cDSyZwwAwtU8+QwUFMYxWDUySLVXirWJjFbM2f/Blq+wkVPBxd
bJFLCGnaPPrGH677p4FbOb7cVwkmSuFNtMrNCx5SW9KliRatW+Fl/3hFanNdurW2kefG7hzhN5TU
0O7cQsbMXsvEAxEdesBpI8Epx+szjyVOTD+0HIfI9WB72YF+Tj4U8Hr/2/HdtNi3HDOMNzSX9YDv
+VEZlKRPUxiMUhtbadqmHYkppDixdPOfxZNUWbIxRBV0ys76sVeFV5deO2WbtEqcV7F+FrVAQfX1
JFp/+YkTYlMslm/Vc3mgnuStJhuttCMSYp6DX6Xh8XxAPONXrDdQp8s+8ifEaZZGraTiPiXcwIiT
hcrJjOc9h4GQDvXSGVEgQWpP1dKxWdi2znEglM9QqB2tfoRHlWeknwRfs6EW8xtlHFj3+X2WTFId
XIw0kFtBtb8VSsfSuBagzspVu/DmEqfbqhVlf1aYECivMup4yIzRHBVKrKcWB19VXjkMMW6zYpuS
lzxG33BPXKi3eb9p80fOKVLQbcY3DXhAoVloohkxU7IRK2AovwUhNwWta3ZYmC1hPG/9qf9luA0N
Z3fZW5XZAq63xAZ/RavoyWnF+JyIOBjaTJHUnPDqMlEwJpfiD7yTYqXAm7KVjLR+lpEFHj8DQT6N
eLirhtd81zOov7jU2+IzDlXgbAD2RhWrRqAORdNULVT/rHMblNdXnvjjSBVBNMFybP0qu+1M9qOv
81PodyQSWwlDBNHpUVwC1c0XJ1u3rJyXTfRAq2fGJui5I9M+6L4IZTBMrYuvuI6D27f1TJ2SN1aV
blh3M9ewoCDq36GJjaGdHQWci22EaKYRTt08CHVx0gXNdXc31V3CgN+bz3mTZ+QejzTtWF43Sq3U
LsQSeh5fzxgfv3NzLaTFK9Nb7rVMG/Yd+ds2eNoY3LLDej2MocQClQFnX2sfGBXqV8Ms0SsZpZ07
AOtZtpLpRk0dwPQ/T1QuHJCAqs6Ip3vk4tw2mAkf6Fid33lXN+4DhhFPm0bEyyPEj2onv4DFh5yF
pvU9/9RoYi0iAhrr84g9wrQrx60IUYInKGH3rFuKX7qyaPSy9V93+MphEE+3ln8hZ1DlNAHkQtYf
YDwJNkgPe3t/7qJc5XAiqCpzuSN6sQ17Isn6ybZYrfstuU6mggT+VWjM7VFu3XpJfI6tQljjJiKf
v6xAgU9Ns4FRJeRpsOOgTuy4GeBit9wxDDjNfsRhmgIi2tGlidtR023YdjI6z4iZUVOmfQ9qWaW4
vF5BvqJBQiBpkoQYCipat8ubZYnkn+D/lcPcvRkpIKlaEixsDLTY/1RJ20vbBTA17C9jh3IudL2u
WaSwPRNN8WblgpdnmLtewbkhK1PD0gqGkjFGStzYUULj3HewZMqfJcHzBxtW62vmPDfO1oqCdF4i
DW3mXbG9VK78OIQEpBlR30iBNvTb5ojUVedmwvnUJi56hbLFdwpMspYACjRFtho9DcFVH8s3hNIj
2JkW2Oh5+fMMW91O60EgBqXDlnkCWdU/K/g73o9BHbMK/wu9P2WYm0lBQvYe4zxeknZ/1R3jPnms
Nyt86Jq/OgHFHOPfa3/amAAueckSEAs74ySLx2kZ5SV61lVvJiZpZdJc4DO9EDFxbHHaeNqYO+Pm
JunA9gjneI4aGX2o6Z+yPWDAn0/GDjO6aVcqoYg/3e8CtJR3CaTdC6LodH4wuahwt8r+t+5WWEk8
d26gNZDyxq+meRVNW7KVqcmdSTzhdfIFb2ZImFb/1OvVCj/S0G7yrYP0IINAxcb3L5sG6FZALB8G
7tEctPrPUH+jnp4ufXZcgofVCXWpjM9+8AWULMuXwymVQrG94h8HFycqHCTilfSF9Yoo1IJULkCV
LhdXaZ4Fo/FGkvU9BCFvA719OWl9mCa1O+QEuFqtAEJzUucSR9ecY27k3cuGrQYSXH0IhF0HkZWy
vn1CJGKMQYfKrXcuAoy/fX50IHPhDswKGMJ7NkTGAB6aWPK6KiSQbCsocXLdjMDVj7l/tf8PPs16
b6EB54BEi2HFxN5pfRb1Rsp6AcJhc0arApH99Magi4XtoHfkc0its+bHJPOmSYaDkkK67WRURFqK
ePLRyGeElwmrfRan0Wyyi10gMO/U19hWwCh2IwaARyQsDNH+KSk+9yRz2d+6c5qN2nuE8GsH0Yjr
v84/R7eRhKjoKvdsS3mAxNfh5Zu1JvBNqOfHa1jArtWwzL3Vtd0xtEmxRei0CTB58kdSwHXi7jTl
Zntzv/91jmRko4F7BgiDaXG/khLoIcIbFtfn/IIpmASUbyU36xUOQACNPTOrP8G9UHUehGQhwE2C
8IhCIx3beOZB8m4ZMPZLKivVTUNwleNz9VV3bIjAlM88R8E4QI5zFvg+Q3ni9a9T6IwJuHRgyn+0
vjoUK0+vtJmT1UDHEvrSlKPYenYLTHa3lqdZYImNgOqgrPDA9s/tyXuIMB8jmGGdRZfpw+T2SbVN
K4B24cHZWm86fFmSTXn9+86NJ3j/911RPg8rRBB2cKOYJuIJjpP1uScS/2y1MRgJzXeMToytaKtc
lWQrkDsaVsL3gSK0s/Qh4FbCUMW3v48LyyX9uFAcES9RTgCeRCkefOhkR6A2FESD6l+yZ/Xj0eN9
GzSriBb493nziOdVlmYKFaR8Fmc+I/q6G8/pCPe6gDVtviJ26r/tlqS+eiO5vA92D80sviFxmyhc
B915FHZSDjLYBaV9g68LXK3bzsjftSnUqOntba35Uql9T+nS9JKGQwOGhOJTYiHKYU+wjiCCv1tK
VdNN0WbA3hUTRvZcJ6ixOMvXT/M/p7PRrYSs5H/WvO9PkMuDPD6R8dUfom8fR26XcrRBB8/oRcaY
v/xaDfS067AQzZjlPvkQznil7rCl7q/KY7epueoWUSa1yVdJ5hVMdXimecMYnaGBVNdNtWTwpeoA
MZ/nQBx93aXb+Z8RQvmbUgKg+rrMOyYc5BWzZILOrYioaWP9GK/WIsClU5VbZs0evB/aL/49/J5O
n+t78m+8jWcdLJmIYZYOyn0gnDmHW0W503yTJWiZRk/7cxT9qtLIp+EM1yPNcsZztoKyDzB/MId8
8/AgoLjrZoiJuy/1vtq0o5tHMQKIw8fO0o3bXWBnv0zZZ2u2LKtn54W750r32tIhg6APQqK2lvT8
mTw0S5J5G9zy+B0fgnf12pDvJzyDfT6uKFQzyUyYhbdPySgWxP7li0q7D7qBO1N4hd2kA9Sqt7bM
WySqu5qeWE6Q8QujWuBbtqEb0zvvzYhoIJ0jyEW0Vo7YCiz4ts02gQqMh5Qklyeca6LYTLjmJbzV
vuwm6AK1+eM4lUlf7kMsRhMrKmk7eV7DJdvRwbe3H+m/eLEJmyauWqmbIB5106Snnx0j2d2Igt1v
QkGCsExQZS1KvTyeyHh6c6Ew3umaZCHi8CjSrKsrHkGWld/0xV/NmupjrQ5Qwu4o2Lrgkg0+n+CZ
QXIe0gI+AAHKBTp2Vh+Eut29y/EbNv87DQczN46NgflZ7cs96iZwpjwx2iP3X00Q47NQZcKAs9HM
9VOPtCNX+glr98oyNCyTw0qrRTDkyqeel9T2lvzY3Xb2UqXwaN7s5k5MQkNKjGWXCKiA2X/na2RT
YkDqkWQk68oNfuJDiE/fCcXZxL8CNw3c+k2+FK08q4hsa39McEPu9dPVvXHkVCB+cl0tp6lNMRhp
V1+UPXJg0CgNWVQ8et/lISgo/XgNuOHep4ifWm2atCTIznNS8ZD+HSmL0qxr7KeGofMf4RNl1QXO
elv7pf2mKFKTYYHlpSDENxm1O9wufjj4gelQtVS263PFUuaRcKZUq3RHRVpQnhonrleGYspxYhpI
UyYVItnT9CeHMmAd49PfgpXFN59duhV3YxJx0Q7LH3tvpON7qslOHwUzeNxOwim7jwC3YHnZaq38
qGvluB5DUf4n+eeUNgdupxNCjosMXUVSsL1zUxpc3LZe+Dw3cWotQqeQ055i+Fo38N2w+kNp/MQ0
tdkt9L99FnTbQ3d7Dk7d0PXnhqGelXYl1I71zWKeCOGv7xcEvtpzglxUjAK3vCEyDXITR0L9YR6V
KaWT4NbtLBvpSmkR8jYeya3SQaybmcjdurnkP48UYu4UrruebQq3kzPkFm1tnYEQuT1jSk0lp4D1
WdvLhNtuapcyGZyGhdnSD/6ZXwEwPb+tHLb0eyzUVZIRULf7p4EffQ7lE3vQGtFY3vUYTpARpGmR
NU6vwvPjIJZm8SKodgc8k9ysEMUu9IBZY/tPS1KSmLD6IqMYq3w/lc8X/qZkohKrQsqp5MNBTrn5
RUbUJxm3vV7UaVkuk1P3mA9MNwmCHF6kv5jsICGaddC0cTyXgi64ZIyZGPc+TrPEQo5xB3SjQ8aW
WiQESbogsDLg7Wyw1Vn9Nvn192DFSGSNWspvl2AZohUUSwUxJWDttGZ0V6SBZydxcImuDXii0y+A
olqlJgi9kHmV7eQafJaBSgo8eXoS16AUZfgxcmMgGxM7DxHHQ4eOq/LJ9PB3wYEBy78/5mK6/qzq
o5FWIRVBe+N5HJopyLlNmWCK8vDyOqEnJJZ53ecSbyQFfr8Hj6fDfrgiDOKReKDBRfBSEgUXkQ5N
JIdfGi0Oq75lo60S0xbGAwR6+JWZ94WJrQ0qY8NKKCnJGzZ52H+cNC4LBbO60yeh1dUUkJB/qugP
xSFd9WvXT8g/o9dIBesvn5FGDRS4es8+WJal8TmqbIq12idOXr08PQwCu4bAay+a6N812Vgp/qRb
d9rtqFpvVoRseOAY4LX8MXzycpOjMCd+vjDF0REjAKcIgcl/qovC3sttCRpPkrSGEg+88w1eMZBh
XxW1FLMM1LUdUQD+96XrXGR5ltT4+A0EH4dLRxpVQ0/8H8XTMRN5CuBRcJmhaEEpFmkKFh+vCwW5
p/gLoq4kbGmhA1DXNhRkL7vTEahT58N10utH2fZFydzbhHhKoefL+fFgr41gQlvksNXneAFVZKCX
L9CEcoHojYEynipSIFsa35JlAKn4XRxZsTgkCNyfGxlx+zw2h85Z9kuGYqVxefYLD6R8hXJxMqOk
KcCDEkJh6yhHbfXuGo9gV21wdfPIF5cayhIYilfBWGA8+VRtZy1HHlE7KRRtvMqKsRBlbUwRURyN
qkGZ0n3YkIh4mqLKt+Ylw5gu3FZFkX08f4iXO2fnxDZkH5FLWYkNMqqkeW1j1Q/mmv95Kf2SDvjO
8xwBOcT+OgEYDgto1SSna8KEzfazvMNOqrC/lHZey617sM820lZeVnhNDgNkjLjbFNDUGiU8IFNP
mum32T8OGEzcKKBZtmQ/RaWi1B/ITM1OL+Bx7Hud6jvwiJhQCsehUVfGjjWZhMuX32RXIRW9K6Y5
32jAZPHFnljY8L+o72opG+usj3jP97YGuBehwtGZmyiE/nWgRlzs/N/lzhAtvV+Ij4jziZ+oNFKs
VP+NawNQudA0ynqpQvZC+7QpZakNL2ESUGrqsLIZu1PjMuSvd7mACY2IIeEpnfF21KKhabPz4ndv
pwwWlIvyen3YRAlkzE4O0fOfHLouVy92g+Hp7D/uIz7fTWmoiDQKycvirh547+XkJv50DOH1DeBn
kkGpHBd1yMz+nPfYQoVNtN/pwcEpvfG6g0RWAIq1dyAuVdQI6h24xk+EOQNFE/vBZMOVRYKvHSnk
X/oAFDWzrpPLAC+gbcW5FtgjE8X4BsBGnE4mlT0MdWjiWApXF1EBZG3XnuiFsmOSHtuNk0/BXM9v
BpeW1SDuEM4FubAjKs8vp0KXs02sruJOC6eym4kzeU+ec0PRTGUU0CUi9ezzKhrBktPYoePBFWgh
dsTost82KTz8gbU55Nigl73wVVGnNkpipWicuFhNfwfd9Hp7tfU0maEw2vC/JDZhcRcCNyWiipyu
6EjTlcOBOQ9TIpw6D14vBMnESv+DGme5fmHSbeERbA0/oJUkVNEJqXergv9UJLdqW7bT2rwt3o1U
R1d/uxoysJdteahF70Bf6hM7+FWAb4fAg83E1q0PsNOYoxqSBcBBepyIRLI+h8X1Vxi2wipU1G1K
h2aerX04vWMDFlNInUofEQInpbdVXCxOkQdNEk9DIx0IVwGD+WsSIyAkMY84kk8ehuvhme9ODiPl
YtBnKAX8XEjq8tq4M0Xs+ks2EoD01anZrAg8ydT1h095nsycv2KW8SJGDzU0MbXhEfLy9PPvjCFP
vta6OQTR5smA9LTSUdOXSu3pJm3nxvK3F99X3I5fEiTUdoa6SeAeEhn2aCTWrdLY9W+g1aw6KFxO
QM7d9blyzFDHkWcUT7gwdTy65FGsDtbiQv4cfhc9L1JFBHu3wZ2XQbjvoe3uOffw8pKThYYV8C7k
/8EzVGnnxT+O4ct7WhCJ81GuNb/BWQHoWkEg+tHjnyzFhB5JYErABXC846mGl+1vC3s/Aar8eDWi
mKsERAfhBw9Hu0bgpw54cnyUREAqUuicHyj5sreoqwrj2Dm9WLMCbPow+hh7py0nDGcCerWKEufO
ZkuPR/qF1ySdYaoW4IcgLeqdCzsrhDNiUDK/pgg7cdoKpnwaauYiopso6l6/WWmuwWe2Q4jxDptv
WIwIAzTTQmUUf3wKhaUrB6TZnNMlxAfrnJDZEoMLCxAVC4U59JC7IpEMIEgWO6XW3/VOiREhhECh
g8eFbfhytYQsVky71MYP9nJlJB2Qf/2u7Epd4PZf0A8ycAeekiu8xYSoxmlE4eBVhLfa16C1p0Ci
qnTLq/yG1NS58keehbhKqCTNcWX0UlSZu9MO1Flr+DPRdhJsprodwVmNx3ZMr4FZwEcHHcLmx0WC
dmj+Mf8sRyWglSgUS1cIZmTrCTbaj4UGSzPzDfKHE7FOqk1VBYSH7jGM7IhvmPKA0kyQ/zL+cP9F
Q8SSM4xS4EIyoS7XwfQRJKkJgNETKIZ81fT12O+DWSXxOpaIZu5t8ZbHAxdNbkfzLXUxdEu/q09O
YG7yMwlWA3cp/OuEFk7z4blLromwwpTgH6rPCxAwf8xNSddTJ3184mC+FYsJKDHJLgAoCNori/I9
KeW7KwS58XbQ2P/uzmEx9d/Ho+EOOWkOxSTkNNWTDSOr2fcTVCdFN3vQ+tI+yJfTlWnUBjfKfhIy
aY0wU1eZgAMOs1WvKzfmmfN5O44rjjfAiezERbNEGUnEd+Cdy6Y3G/BFVW9tLEM0zzAX3rG96lw5
xUNzrD4hkI+fP2/avaUNLxkGypD+ofcSPdzG17QL4aLHjbkpQdF7lbBkxTmHxOd5JA0BZ2fpgk8B
crlzU4n8MlCvSrk2wdg0A6n4DvMIuiws58F6w6CFo/Mffw0/KPU6s0pvH3CmuG/2IjFduwbQY3lC
CaT3dggMwry1mESWeCcIkAe4bivPGz5w74X6jD7+qp400FtIUOpd6zPJyNgURNtrsG3YVbw3XsSP
aLlw3FnJehS1IHMPZJB2Fz0603MEsB3Q9puFhoIJ0vxFWN1qNmAaIU1KSlLZZ5DSG5uEVGh5cQAj
quWmk7QxxtOXT6r00A7rjeQ8Q1WIAPbD5zJdc3F7DywctaYBcpi05wLznk0lmMxfK/dOPK2K41ui
5oSLoYgMDyaml5F7iy4DPj2kd3hvhdMKyONLAVvH+NNy+6fuhAoTdGiIjRqW9ziW8qP+AdOrzHsJ
djnJvBwohyqOqmVWdz66kWCHzhbS/Kw79GtRqn1CFNBh1jA68yqbNdpOESDvln540PSmn451DHrj
mS8dOQzN925K0lWHNTkFco/FxMUVUsPkfYKzwYeG4Vjg3zlDkfG3P2ooDUn3sniG2+tKGQqW+9GG
6oioz38/lCxMpE82ifg5JBU+iMZBcjwe3YEeD8Agefdk3DWoYQrvJX7Tv9mcdsr+Hk8E80umOBBO
hLhpR5UPDlcjowqyDLlu55KVHwm780jYayeA2qn5l8CQBy8EJTQlFzGY3vMoHIy8FEH+qN3PJPuz
CiaUCjTY3a/h0r8jv1HzN3aIxBlQtlJ5eN+01+1roVa1PxYNW13AUWNiXG+i0aKA6j0R6KWBB9ow
HBqCD6z0TIAl9/R6jFHjLQ0b/OKq7vcDkOgr6vNHWnGvj4qlVT98ISPUECcxxorL/RxFmUmCOubA
9ZgkZwlb/H3l5Tz2XyGxOA0tRs76cMgySZReip0qIubUK24NAB/Ev7dV3bJgpFmLJXYIulc1EMnO
zo4eyDaVUghttSfpmP3CnBTZKU8iRbCuCU5cN4ykxK0szAtYxIIlWEFZW0sbOkACfxAPCVrjhwfx
7MCkfF2V2a/CCEqcTPzAS/qTY7YPtxk5ETyoF1W4VI8f15exERiOCOugAaH9v+EZ2GcHiSFEvyyv
sFxwxGcygLP9+vFoj5BWT+TnJqe1wIuN3boG5ZyCut+SDAo/sMtLFnKPn6AwyWzWQ4JWkN0YZmX+
QZ7pJmvlqEpOIfQ9NH31NjDm9Kr8Imt7lwmVBqdFhY9u1dBFWE9Z3GKqhbQ6P+eUaksEHRqGhPkF
e5ygxom3VPUmT85rAGJAloBOA3cci1KmDh99+yMR9Pl0bRSSP/0YSfu6gT6RyJrjGZEq8nAxNfML
DfSYQ3eCL+c8xuqaBVppE4MLZJqF1yUDxH0mtmTq4kqnHEqqxmua1aAuv710OOetPeiBmlg7Gxv1
XLG/NVsGHGvCb+X9XIjto6yEj7RpM3Y/O0OmP5swrAqo50mh6BDyNnmD71K9m+DpzeMDcV2CDuyy
Kog624R7cGa0aWjuMNGvafGB3kAGf4I7Slr/KZVDilAMf039+OOfYXW3w+qQrYKXxwXqysVq3QXZ
54O4uk5rqjUpoiij8ZV9AHudG9yCACiJiP4hvz9M0a38Mh8gIYw8cL9de0zi/px7cdP2bUpWkMc0
QxVG83njR5soc8iN/4TjG8bSbtxGeW2RFUMVyHylV8uYGrgd9tZwnn+X/IppbC30vO/UiFIKAT71
DY8KVi74/zfm4kul15kPIS3fPRAoi4L3lEnM1IpRV974r4lVHcLoBJoWZ7WkOEHMsWq5lszOkTtS
Jt59b6ZnxDLZslKwkgZcqZh/361+h5UBQLJH1L5IHiKiFp+f0Gh1ot6JZPAqwCq0o5m6UNcfqx8L
hBrAL5XP0nFNOMTBf2ZNxrlR9VLSeMMlxmMLFq+dGIQDUs57+KRdTmi15xDbP2zo7C2E2QKCtRmY
szu+vvie4UJpjI4qOV0TPKbxzEUhZaJJ03mVvPlssllRFODgfkhLbsYMJ3HxrjxVRGx+Yc8D6Me0
lFwUeXNbhl/56OPt4b7R7VlXnEkjXUa3MDpdyqRe+4PBQPQHoTbnRWsahumF7388FemzQF/O391z
2ZDfzfmniyTthoa0VAXLTelEIlYtIJ0WAo/4yrNO/L9HUnRbwDmabqdHc+DApSFPDi4g3p2cQH3L
jdQaVSlkHypz1VoO5Y2Lcw7IIu1VYZwg2rSRPA7S+Csy47BVtimNDfm1uvs2OFxv4CGCF4iiwkM1
Ku9q5RuKfSJ3ftgKHS49ddmPeoDjHgzeZasu8MRHLYAE7XaFRZZr2UgIEEKt5Ib3p2+63Vk++Rd6
28jYlV8dF/sxZFiAwA7Be8PkwMTpb9/cfzjajmv5m14x1YK1ztbwCPOg3rrdh1QePAWO9EzY9siK
txMgiMEPYguPro/KpZS9Ljy6wCOSE/34Q+xtPaVuYDQmlrFIaJ35MvQ3qdCQXeMN6QR00MkMNkcR
V5LWKg1tU3ghz3W+kOZRwUIxBvpIUy9JbfkVnPwyUj2gOtVDF7q/uJi6M81M4Hpc8FEIZ6Wi50nd
gwvL/L437FqNcGK3aF+ZrVe9e9CLIRYpT2u2V0sk6jXBCOc51MqRjUrD2rhCLYqWh7kqJSc+4ycL
k8X8co/uRSWxhKSvkbJHhYjkePYZWX7mxMxyT6euYAiJk8IZZzrwt5uw7D3ic7Bcqehs9yHh98XL
1A205m9G+z4PqgA4S2jh7sv2nmUda7DbL+sVHXE4nMn7mk3fHb513csdI/7+ayN5eFlPpjwGxsNb
QFUtdlNsYnhQZJ8Y5JsSAaYYGgnSTPY3LdjnhAaMJamIz7u6GhrhjyaHnIclKvreX0OyWIEjwZ0M
9snc5Pn/gXFakjiOzlzI1ETp8cDjRroWBzSCSZgdkTP9rUZAoMReDZ0ne1ZlU/+aFxPBqeB42a/9
u3+V9/N0X4HV8hex+UhYppzPBLeUf5vIXDpgEI7+tY8n9F1gCNgsNVKhG21JE3Jr454B4ioCPROl
Lugeke0u1hz56tp5v+MMK0OJZGmAspn8TZK+pTleIYsa0saWJCNR3l546HGCmAmPBTpl02p1VYON
95KZBTGNEBcck0yd7cXE2Q6MCQvH3vAxkM2BFUOHWoCnOLvlPA6+ChfuJkm0LTTJDVryBk5GJRBt
EG/bUSJWO5aBskzdLd+p3IGB63G29oErlhADfA8WNDKQxqNb6yEYsHdijnUc7MZ8O6TL2balsvyV
rkeFshl0tWLi4/DgikBwx0szdD2gTs6pPy2QM9yYOLnDGL0DtOcosUuXSCeUXNGd5/Ndb8KqzGZY
aRQyK+j6Tdsz88UD4dFfxpkYHcex0dgabnxR2D7YJ2SpjJl1+4f3edfg9iSzIn1VlbnlPcU/odxW
q2zL5120Ec3A0FLIC1ZmJlw0zjPy/CAVB8fh8E1GJy5mHRBeBq4B60ZKHMLnnqWqQVkrHVB0zTdG
DiVJr0Oqkt5VQJTB06Xq5siC7/tnAOEqJJudYOYaFWSW+j/MdyosJ4N9qChhPQ50JtgnFAnlY3tb
YyMfsB4pmW2xgYBrgIF9Mzna0/BwauZgwzELX50hEEPUk8JEHceeV0F7N1VOUyfDjHAVyOR8OdKP
frb26xwZ9dtLwwvlaPELZeKQ+3SrKZv2siclaFcBzXu3PmgWPuiTHbGdhOnA5TVz78flqHoDIvs3
53fD+dxBUFBosvJ+cHQNONSU7azuErEHyQPlM/+J7BseGiTLFMdPtQk8rpTFnjak52pI2BBaceoO
KFP10/gJdmNGWWSZiq6mOt96JtYTKJQUx69HX39rnw5tZfY80pqvm5PivfPXaorBUGfV/TzMRh7+
58dAXClbAEnH13vQ7hH0NaxqX8G+/oQTiKvvFpwBqEx+IE99RzbSFj6EzVOFlUCAO7wxPSbfvu+1
rmYNCwIALmus6Ug2Eg2M+XZh6AqKYhZ8s/rjfTeCRiwTrq0mFau8uCQt4rEjyTXVNH0kxXlZ2sFz
3urRQ1VRGLfUHhH7FQixJvpfvKvflOsde7ezRe1rGn3VakroCI1WJ3/j0NYTHKJBjT/h7hbJolU6
FlPYTp0oyfre9RkV0zM742VIJbmPnx5mYD+qwbUXTuawmQEzhqGQ8udeGLYizoY0ccOvNlzJdrdr
BZDNuw/opn/UY5/roOwT31V++tidBBhQcS2/OiAKYbGaHWAxvTQrBj1rvPPgqh6ZFwTEanbK7K5W
B8CxPCqO7gloztldNGr+hcc2BLnoFPZnjY/S13Dw6DvYE3X51qzkfXrh2iWWzoDOMrfdaMSZSoXA
w5s8+2gJqTPcQNJZmSLrGuROf8EQeod1gudt5UxNvhSWTaPMwq9KROyJ2ud086ZcPpVkC9gGGoIB
hlkl9JGKE7xSvjOlVSR5CuzKsT5rlaVpQvMz/5YwiYpyagHXTzC06rIvumyT1Qq2+oQAblKD5ab1
Nl+/Js35c3nKp8ycNFuLx6VwLv0rBlSSkdA+ZBhZdhQaHLqG0SnlcUGwcXoFVHBTaa5vJXPDF/rB
yX4ASiNVBJEnGMuOn/97zUmcZ4G6x/6OlO3WrkLIEw9yxbY8k8PBsK0MkAxW/XIIPvdG8yNuTogz
tE2iUSYHf9beNBdL9ggnOBIuAIRjvVkKgEwK+gBJ+lQ3J7vRcehdpn0a1UkSC2re+zaU6SDv5Rwp
Hm79S9QeM8ChoQC0FRW9llacbXmwpR1+v/ATCdr0JZBBVlclkHsEa38S/Ku9UOWg0MCtZktnviYQ
k0m1Wb/Ct74iNKcEhanRBNcO1bfJXEUIhobksJipb7jKu6mw8bDYriUc/322cpaPqt6KCILz9p4i
wfX9C4AUj+0l3zcRb4LQCy+ROlOIV7O21d4i3NHk7Bkk0YjIS7OWt5MsSDYYuO7D1jOvq7UCWmTG
ws2Ek6J5nLy02Gw71mZh5c2pL9pxUBjUCvwtfyQvt7U38vcwYBr3gEJmuY+1l5b/jOtUU3ZaW0mB
WYNdsuDUduuqv2p8uz6IkaVs53uo2yjVWa0EuWuvTX4iLzrmiDAQDZbLwiornwBTlXN9vTOakTvZ
GS/CUiqOV3bdtyhyRzpIUusRPeTS+8EvXflwoRTxzTLVOboArULuBs04JRPy/8QY3t17InzHfCsx
ZndVQ/Lw3SYaUwqFOeN4gp1d5DiBdOj2dVclZAhiO33eSvOrd0HFWPiLJaQN26qwkuQwrtMt86DL
ivP5NbbZ0NoAXhILQfbKUIpljZBLYO3KeiM9VajsAVml81x6evEJ6cunze5kzN8oca++MaHPrjKS
bEaGSlb2sdIJgw0I2YEBz39TEwyddgivVxUvKeqBBv0orp0jQ0IDrCl9q7RALZUzh9qLZKblfEF4
fN81si+KAb8xnzJbNPngd4glG++bFVZXivcgYYe/2h8EBdVHXHznY8iH+GCvauka9Z8Eq8xsRyze
st1ikHVCHkZ1tV88Xzmibp26cj4fWyvQ9aqP7HjV7yId//jPLI5oQ+9rxv995FeSNF5Se3mpx8ee
SdlMVxbPr4JLrrdQvlYsJ+ih8OGWCiWlQWA7m90AvbWKErrcrCRkAYjOQJdyU0k8Sfym00+6oaYK
QnSGN4rOekyAJWI3L2jO2q1h3rV8Hem5oRwmkwKUUki2PbBTLkfh9PqKeXXQInVOm2cWZsSoeZTo
vpwoTI/Fr5Py+v/wz5Ur2lc5uop/kW4Bjjcd6QzZ9+rZ/CcHov2Jo0D9Kzk4srqyiNiMQq44V+ve
3eCdiqvXX0TqrwuwgKr7rN6IUBRL8g7ZOp7LklEUrDZXI9/EsFI9lrur5yXLrind/hnbj0035xXh
C8Qov7j2HZKIr6ntKXKXAak8nFCZbmeBMoNWz6AdfdOZaJvPZAFltVAz3XS6hf/ncWPhWH7i7Af2
kgyU0pvwP+DEcaodcJ6Nw0aKChIeXs8tHDdimrgoDo2PcwhnC2Xml09HHd/nCbvwAGhVsp8wzq5G
tlgyoMlLbTeM8kjgPzSmxMUnPBecZmejvTlAjzEMWyLG3Vv51u2CAfBttMhLyLTjjpV14nCigy1X
wh689LI/waR3jexdRlF62n4e1qz2hMfcSMvNrrykK9ehW32bPGooDN7w+nLhtNbcnl+3ta0/Ua95
asib8sZ7Rt4YTRPxNr/0Ea/dW8w3kn408489YCtRR6sa5Z6y8Xxnz+KmGTNDM7UMfaWJqPleWWqW
TibnpqyBJEK7UJM5FNETTvxIVKVy0bUrwgu1v+8hWP31j5jSIMVjEHGSThqseJ4Wep8QRIUVrqt3
o22DtfKt5Pg0ePaN+s0qV+LpQgjIUToxQY0bkFSMygklnvZqcv1YMUAwrrh0B4PE9oBQaKpSjEDa
b95mVmjlOBaOQuoPdsnkU2FUUVKXw7/r/lemOMj/p7cRMQsXZ5shZ6kjqx+PpiD68lmjdjG6uNWb
7EaWwC2wsqf1COgPdaqcZFRKOqUdWWONugjZr8O7AOXVDuCfN11p2or/wA+k6pRtrw0FpghALgrt
umm2sYcfqlE/am/xekDXVRohFrJ1R2VPi7UYgfxSqum9bABvl1tmM8nc3F9KLm6YgpYwKZ5MV4UT
ACYCYrL/Miuw4n/rY62JHc/Xjk1gfc1aINYMwKx+Ol+tAZ0gl9jIstCKtS2cbxnxhBbDroB/Z/Pu
FlBkjQzfIJNR03UwZqNJwCc4SuHJC7nH55iodUOb0lHX6KhdYIUk+DJXs80vNRfv0Jerw32zSL1n
ByPJrLLdIX6EUPlTt04/Q6HfpuYWpMWJT/TtStzWD8Z3nR/+mTcP0giNOSylX9lQlmGL2asdp4US
HpacB4xftdzMrnjYdZ23ipYCBRn3Eln+5JaIrD4RpHa3mARehqhGod/5Yeu2vWBABZRqspbgZV8+
VbncUUE5eul2jOg4mLAsUjfA4gQiicOBUwcaY3hyPC8eKAlX6kQPwdGl+TwR5GRVF/CLdHlcF7a3
YdQo/M4mMdjKfVp6LqvBd/nCumZ5zH+/Tocy+iTvNDE+XdyaodIH04Bb3wOTViaACL/yilDtq2se
4g0L86c4gp/PpNL4eriTZ4EkOySXjnwo24CxSAiles1zdVxEjVCrIWZIAG3aH26mlgIQ2AjwmmuE
7GV2jCn7Bfd1SeNbv2/aRh9K9HNy+hV5z6OYDhS1abenTmmc3dW2fpIPN9ER9RrVo6PsmwhlDrja
fKTPXsd3+2BIRFMLAxyx1/JiFG9DlXV5VABHgta4CRIbfkJp+uOtmUa1DvZG2Af/Hh5kB+q1/+EX
2TPxfCzsWa71zcCZW3tIqX/V8mfJVsqlmnGcppLLniKlUMgrjKdL6kS3RUQit9UqWXCtE+Oc2b/5
QqIq0fcTrmM/yF62ztE52XN7owM9LxVCQO7wUdoFbosCr7xo0+x7EDDFh11qlxNLt4gzbg8Z5C96
FVNsLtcp6Bv8+Pnr+0YYuu56050Hz8JGdAI7EQXwUWrZnTJTl0PN0M+Ngnjqo6Hbs+9E/rdsPdQx
HCpwLXdz39Nco+HL4xROSlhLBLktFWIiIbAuc0dnL2FkQG4jhc+ktQDo30DEG0sN4r23Xw3Cbfad
vXy4qKwUFyvffD0CGaUfvYrs5TyYf4q671iNSVqddeO3zyND4HbH+0vyc42xFLDjx2ChARi/PrfT
7UUylOsKX7em/qFwzSUJ+iSN2ncCGiSSWrKL3cs1FGMxHhBccfEhseP0G23wdKcaoKgwQrDL4w5N
CVXwzvsUr34Ihhs0shg1Wn5fhvgDLIBGrIolR2ZLMttEpVY0D53j8IJ7ht9ZV62l0u0wEYngriyR
QuXXW6/WPFZeSYBFbCiXJeFJ7boYDOTEtUtV1dHHdzTEnmZjoV/M5+JyeJxSyL9k4T0McdTCgdUM
RDRd30/gSM7hRiOzWit1x2jmWeHFkjgo7TjsEwao1RSrt7h8NEGGV7Q+SZAxnTiVNV2JLj5yhvbM
Vd6TO//ZPwKIxLcRkiTHhSqDxqp+3XFAmBp/GiAsVzNOGhrN1K3wNoP+/DHFV+4jxGXncowRdzH7
sfGKH7YFwLts9mZgClsVru+pUSm/PLGrroI8VIwOhrg995c46zsl5iT8B1h8/u1i0JCVAyMLg09u
unAtQqUFyND5ExIN8yBfNoUzaPtLkfSgouVEiEOUAPHvTjyaIGpZMhsoVtMy4Zx0mtL1we2Dsngo
+a9tk30k+oaBjUoFu4/KDJ81qssN7aK0jE7eAi/TpAt50XXlQ0rP39i9WhXvBCGcPABe7rnEw5ut
CbOH0KEyaH9hXdkJpzsuDHQAAngrSaUumiTK9FuEiYMgq4tc1Aqa3djhowrh+5KV5nsfThrzofIQ
J21zVFiUk8ciTGGkCBK3KkFChFjhWXcc8NTBdrrTOBHAZcEGldPH8bSyrKQIV4/0Q5dkZRUG4GJE
tS1lwURkB+nn3zqjUsXrfEtBCJoSr4j+5MOBeYW132jsCF/6ZVSubdaY0KrNmBmpUMv374tcnwf9
/L/0kkcNhi+eyEoJGyEpVKqIo8/oKZAsn+hxWnpcsMRbyymAvL4T8zHrMMOxGvPvmPsA3ov4l36x
alIGBWcpWjLfWn9248njmEm1ooGjBqNS21htf4bNQ0+9ZQ08b0dIFN7KuMg0WzNz5lBFBBvikLmw
aGI2wjJTtVGVy2xcOKc7MkFoz5cooz2jY/PGlw9nFt5KPHU99TACn3GLeJHPdg5Xatdfu0zLxeYj
sTyI76kv/j3tuxrzB/4DXFBgFU/g1y5ygom6EWEcvMtLNTpDemOm/elvv1L8Q1jIXJkfCTM9y/0m
65qEl7dliUM7n3q5NOv+x+9ak2ijJgzgA+mlZXL5qM+Ec+MTWauAA6ODk74HkySdXRH28eg2MosI
BtUdYpti+jnUOPC+TtnPwRQx4UWPw0Fm4yeIIQkM7tSb1x/koHqCajl+d1sUg+jO9Bs83WgA99t2
jW4BKKTelhcQkBVk1EZrKyvGLaZI4nTTA7XzYNBmZyHWQE2QZiCtkLYwC8byKgcOPq4HumZTU5+k
s7Kp2txHvGgIb2vKk+V53rfgZ6x+ua0BENYLYGwO0FV0r+D1zqww2TPAQ6T/QkIHnijGTlri5ayL
6zQjn9mAQUeSEi/wJV5tXZcor92C4LGNlPRjSAtp16QUz+K6JjoTuLMBAMVdgsFoxMtQgshF9u10
wjtZttcl/DFVywG2DHqzCEWmdbHXHX3gjDxcVTLp9mXOzShCTH3Oo9wBjjo5QE45CoY36F8Og0/B
hu4hfiq+LvvCZee3Zyeb6szbSZQhtKYlvFxHhb09lvaDNdwdEBZvPabRFw3D1HIzuLMQbUd220cR
9hJ27zFcx9b8AxssfzqUtzeDwUtUqz4qaWrR4qa2cxMkpgAkaK2OA3CZ9HGnMKPMBmVoWIxN8D6P
S6KD6fTnwck3ckkOqwTjv+i0RzxsLFNbbZ9/HuXUzW1C+Vf5JW5ur5BHgzEo1IUFUOMPxrayv4RE
JpJyp4wp3VZPs+zQFRfo243lj+r7KCSY+veug+xFp0HPjnGSlyuvgLlwzn0JWqYD+L4oP188XjNm
0q6xAThyJ4mMQ2bgh0qXmj8rUizEgLiAPgOQ0ZJAUacy+0yJIq6aU2W3AkLYbxfHalG4RlJkFC1C
wrhImBq2ajcF5ffsK0GLPb39YlVoEa13RI+LQeSR/BefaiqFqmjPlZ+WdcxPltvfzRZ/k9mjHtN9
+lgYYv8N0KUVlgi6IoKXSx3r+b16XcEv2UpYwkgrwRJzNYQ8TlJhFGuYmJy3djFBkYhKV9vuh9uY
k/Wxw5NIn9grvUc+GHNs7pVo7brjUyTnBBbZ710ozQegIqZsSAd3VHvleVY16A5CAlY/+EDdH3xo
/dLygE3ymMQNvbp/94w3GpPwApyRsly3JHJ46viF8quDvlafo9nljbMgNYzsfWQF9zX+LyLN9twU
0kM6UQa2hcyUiOc26P8BG1HXBhE51ddtxTAdnkHowhG86v83VS1CvaZrI0k4W+bOjaUc86CPqOt4
14jjKr1dO3/fjAzRabIfhXT5bp9wDRizPH6HWeBswK9g443dtt/sLsiNtG4KO+8E/aNDQMVQckCR
5ew3227HYU6dDSiy7frhcYm8QmElBd0zzvDHTCIQR37/rfkCooo75pKmr0RfXnDyQzq2+f7HSPSX
3a+9KComTZxq+6elktHW/phVxRqSBPYjfkqy5PCKRIiGVzc6D1LIi66mZYK2VrcEjAoopac9ZiUG
78eHHIZrRapKG+zJK4fFl/WgW+oC7XnsfGuNIkKY5GfT6IaeHkfBwmzCWzk7P5JPgWBdylb+fWEV
Lw8vqgk2gHiI30xV14QtrnAWR9AKsqWIDVosdyFFpbyub65VYY3yMc8p3bODkhIL/nWeRopM5rw6
zagRbcUa9rl18AoPBgYafAfCZfzb3FJkyayWYGLuaPB+XwumwlT31kaMuezxX80uv+B3Fdy1abyw
fPSB/xzuxXUDR+RX+Yy8TF/affmiTHNMkRPgKoRILQLD0LGsvyvSINnP+e5UuDKs1sXDrkSg3QHN
1UdHaaghP2ISObEJS3kWRbmy4NvxtAtNMkzcfRoasqJNd8j0jlfv++c0oAMRAto+Y8FoqLnrTdqW
V/EJZ6/p4T/umUIG6GAeHchxD309vUscVaaS2Gcaf/0jQ9HatR/1u9+lD7aCPiuzLPS7w6NaF17G
jgOFshlGJdTY2sug6VEqTd/cl6R51RPti6L5HhBJzmKHStwqj+iFBg11YVn3Q/WNo2yyWGc0ZZ47
mT38Xzh4EEHyPGw56/MbNMdnwdKPJ29nS22PROejBVByBvL9lttZUHh0w2SS0ZbWjmQ1ZCQ3QjBr
yAfmUV90ZClWoj0SRNDmAh4yojqqpcPfpJli/FVa4D5/Xxga8SFvkObK7p+dvyWt/q0mZwY4mENf
nWFQ8CjWKMKQ4iUDhluQYlGKhdEO53+XsU6onjbyLpq+eEBU54mbQp3uQjSwkFUWKYgExGjHItEE
G/hqqjsNfgG7idZBkzBVGV1WVK4nIZqTkXYcjFwqzgnnC+R+EIyL3n+ZVJnAqSv1lCHUjOG3mmxp
P+ULawIeu8+KLAuy3svgXAuQsbZuOMM2wxmSwCevHJsI4X7oCJloTDmiPbVqcv8xkiRkF+6Xj+vW
BA4v3lfVl+sNiyAoxefigSZ3Lq785nr9l0VyCcOC+b3b1MUW0PZhKkSpjhvySoNKIK32sdbuikZC
hOCvhg3oJL/I64HCtN61ED4j4YNn2pzBDI5j8n05BevtYcw4+3SF0DRkEOYE4JT+uhzFmE4CVVp0
KpsCLjbZXieLnBIuJKDsfifWSG7shJ0hDcY53sqV1KFKpIlSbhOeFPtJqUUw8cymPxa2vN5G2nO6
Lx8i+ko8WfH3sNhjc47Gnyglj5IFBCCBrtv49ilRD/cor0bd1v/LqsL4K+y+5P6jk5ZZm4jF9FBc
ToLREIR9K8CVL91FFQLl2HVD0wvreSntPA5WagnMoMfKgBYWZu0gaOHuOOQW0nveiFxs1tvD/ejE
wisoQKsN48xF7KEtkgocApMG98yMt5+pOL1zHgwL+sZjPvzw6ipfPbmloz5jcY+l16SBypAuHuiY
HTMROnSWFQ66WeJsJvpLuQTnJLb3rBM2xxTPPi56ZMlTIbC5Y4d3iMsZF0gtqr2h7dYE74uUSvPX
gKdZHCl74owLb1/rwzVtXERObTdUwBtp6Wh0TkWTJ1X1UORnNzbE0WXAJIlZRxruySpQqRrQ/VMv
8PIoKpPdkSBM39ETh3Qrmr4oaqmVZrM61RtciTfLa3v+VDocVF7vOdDWuHcsacwNbMwffXKVPw0G
8eiEF+qMg0V01oLVVD/OHe2e9BMmkcnVggr6iBLySSOIseLJYrVOfsaR58r7jdnmxdpwW89bgywk
U4SfY+c7GJFXwArl3cFlj8EVf7xhoK+t6Zc19KXO/TxynypFR3KBglMgaRLoCzhWAFRORcEU8CZs
ZcP3t13dXigohDkFCmcwBhdnP40THFhFBdXeX4n+U0yr0tbw9CcjRhkapuowIvvpt+eoLFGKimCn
2emK3yJBBSuCdDkRRKnJEKCStiGAHv67IjoXR8VxJ1qwUz+RB6yTFQACTtt0jeE/pBwAtownY+MO
JB8bJCjc5BJxzU5orOBnLu8GXHcqv3VsnpdN9wtynfljHJ7MuQzsKyLp/v0lg/Jt1pKSZ6hGhEtW
eQWi4d1xZIIJS8bMnGAg/1jRIGmyvUHpx7i4/C6govfUhP+ktSwYP+Q0BOE7kAP1l1x2XqhOqKaL
5kAZ4UUAQvV8Z9NwignnbodwDmFURc/7Tp4dq82axuHe6EdasJ0DE6Q35T/o+DWG5+CP7DYXysni
MzlMR8Ar5oErd6hd58oQHfHv05lNpa1cEfs12Q6klifE/Yzu1Tt4cjbPAAWbYh/r3hXSpxNzbd/K
7sAysINxghMVEWk+qUR6K5ygX+J3aEaein0vUz2H16USv1IZazKmFM+4CwIL4hEKcJyyrztFVDZV
i0OgdPqM/xB1cWMQ5Y/1JoNcjCWHEChmQDXAfmU9HIRtbFTK2vy3rWg+cLjF2XoeRS3RaEr4Qp0/
Y2MVzeiaDy0lS0mfh3Rtcvhsl/xO4VfH2w27yuCMAz1FU0VbAmk3WJ6wlG+T6GQNLiXaB99vYmAj
1OuYmX7IUFWyhWYSjKFJzUw1da/ikwNy5K368BduTnRb9YGy85VNSwvo7OCEQnx1f8fhb7PeeIVw
ENC6Z3wuWcsIvtUfQSZUUygfS3XUJqfL4AK12S/PkGCOzuN8tFt3+mbYCNmgf5BUu3NkUH9c0Pik
sLe7UPbCUIlMtGrnPdcArb6ax5JbpHKbFO+8SzzIvFyzfL5Hz+KffHVh7Xn+O88LDQ9DMCJztw4j
tMGM59U2PeXMWvGpKesO9j+ggVhcwukNUsar1i9lPqOYArLJ6b59hhZ9UbRJi1t2NXjfxfxtwish
4gnVcX+xMLmSOT0CKzmH1GB48TIjQx9geBsd+W/cuTxOhgAyymi6Dfzq35j5PHWJCpjowgtN0Q+J
d5ahWFNeuxDhrTk6a4UH1oh3bYw39eJ0kCMo8OocSXQFA0Abuquu3DBul6A2CA4hR4Y83yBM1iS3
qBOD0ZTAJqH8PaTMZvwUc+Xe2LfjDNn7cw9J/JmegEC7Lm7NfRxOwxm52t2ei4qL2MQablUZgj44
o6qL02YcQ1luq6qYmglFXCkfdkfKY/OxBsaEyvzjXcMIiRbBjl2QwSjIdFF7JCqe5c5iZb11s2gH
Fi362v8uTVimhEZnoxEfaEqWWxivaLvcVJmjRnXc5R3KnyjznymY/QELrwy+CC+RKlEQ4lW71T3n
5jSlfNCq6b9OreWynZasx82Z0IEHW1JaUb5vpqmdIh1LLVRa2UsIrfkacXDFzcyldDfHUDiiOs5Q
ua3sdMKjI9cx3PgZ1hVt4xOy34tRh1wyfDG0zZGIabstZvRxMBI0zrY456CQJzNkkd0zs/AuLqmy
96dTfH08OFhXbwCNERWcjLa9rWpQRj7EAM+pGLDlLkg4qHG8w14XEvNgzgc+9L2tkVeOCgpNZyzY
vORfo1KnY2SkLoc7/9mJKKnB+XXqp/JZQl0M7S+lDDlhX8+EW/kggvPxXytAjqGcwoBoX4vXW3V4
1m2Ld6fb/kVu080OBuLcMbJNd0Oyb22BdGMTVgJ1f69QkxHr4XfndqUazFUxf5VeEI13ZJs/7okY
us1L+pqifrO1PrjsTVXsS9n9+iBAaWmtrg3zQ/fhq+hppkXe/79xtkYU2uPBg8p/vJaF63DtYoWL
18QobbpXG9j6/88QOouqrPIQnO3nfIsnLKjTkyUyAkAzgBJNu7xfelIPDRJyfK4WfnlgoatmxEbK
b/JDY9pGXng0wdNflSs3kROmEGCy9+QCcJcjxGhsfyQwuPr6SIHE69BYD8uR665BZWiDb6ktLKLg
IQ4UvJNtdM6VVXRUQMpHVokc+7TNTsoqaTnsZPAIfBjcaeVuLOhWdjbFVJPdmzF5TvldIyTeuWqn
30XtYMGcK/tYUNhf90gc5JPy+fVtmTFKALgyZ6UCNJL5yeWfLkFEm1dO+avNqwLqMFwEBhO7hLlL
SQv6GEBdAbHp1qxI8dh+afsFJk5xUdvq0Qa0k9tomqvK9WlCLHW/i1wUSrBLhMOgDHb4En1CNLBy
h2JY0rJ1jtynShLKF6OK/aG0d8lH7iLQaKHzlzoaLzbh1N9GgmKkHoDXRGffIwdAc8JujLDFg18D
qB80gU3yrke77YY1M56Ycl70CbxvKwAesxFiieqKLs0Zody7mXklmHOMgPCmtPqiscNn9zIptcJx
vfNlJPb3+jEKG0drOCEvQkr2f0wumURmXUCyt3EExYsK69CBL2U9GvtUwk/sbiEDnO0fwgOKOE1f
3c4+oBtsci/3RCByTFb18Of2Gjdt+UNJsj48XSZEQWx06RXu+OxMR+O3jFBN+kAiVmbi68OjjPy2
df4MsASrk+mlSM/GeIllAl3UeaRG83Ky4Wjx9U5V93pzh2GLZm5SF5N23VtS/a5IYZ/NSxOWFPAE
D7zF2dM6gsWyBn8g0kULgX8Q0i15VFP7TMYu2PESNq9UwT2KDlwlrCR8Zl+vi6Q+ynC2IshRWk9Y
igdlRCXuKmtr1Tqs6/mZD/8rrg6Rq+AitfHkniHfpZAUE4ZfHJP+6C4EefPgXyqg5hKMIwI4rjN9
L5hJfPM3Fwa7JyVR0pvxdkrU8AxVg/5ROZ322qg7oyVhg3GX1fcRis1FKSO61CpAMSY1MAPhT66n
VNbnYPhePtWXv7s/kjV1b3VqoDQ0X+dlVWz8yrD/X5gFRSA9Ia60yHuDKAwwDuhUtId2yngbQbLJ
vFj0JASzU713Bfz+75fSYuVyMaX5F+WtQOpyBioaf95p4/wbHi3gicLPgXQP8D9YU5DE1DkIr7CT
C5s4RQhvLC5CPTboSp78op3Z5ZbG1mL8ZgfF1X6ibFmNLPAKch9BUQ5gUZMwnvxUJ7DbajL5lX9y
H6Hy2XwpikopT78V4LAg3YXOGGaRpQFdZ5TWXyrsjRaYA1TlZnNVm5IsfmJoH/ff+lYfVwGtTsjH
RmbljYdeauHXoZyc8eVWzdg9ZHeyLQVxpGpAE00pV03OLrXhRX2q5Djz8bJw+x5CmN9kIMdYJIQB
NErWoa60piEL2Gn6eLvqiCbmL209NwnWJyA+JAvceEt3Cuv6t7uAMmU90Bbv39ZtrhBDTSbZIQc6
IsoCL7nAjisUgZSXT7V3Ph72a1ijWCa/K55tXScW6FktHqyrRCO0Sxw+pA1TfeB6caLRJ62j6Hcc
HxqI+Q5ZoP9ks2AtEspMQwKR+WIqnP67F9vlhAz5OUJs4TBUnz55Rug/BGs1N05varcOskfEQiwz
sBdfAS083LWDNVqkCxsvXyLBBpKyQPOeR5KicIA217r145I6vCfuV46N4I4WsmLs+xVq7RPU+RVL
TETH61GFu9mOBVS8WGY54NltJI3iVznof4P8UrNmbnHKmREK6psoWaRkGUDttu3obvmR5YJkaWq9
za4ct2nA15Bsh1JMKQlp7skNspZrEPw4uX9GT3Wvq5aZrCMJ9TW3tFJtj0NUroEG3iV1lBcjcK3e
ZB+RFeLEcXHyvJoe4JJaZZ1R7jkSBwsyGBCbibNwSdKe1a2vQs2GVvn+uVctPjpDnKmXHhy1crJ1
AsflfpGmhMyTUwAc7YnCi/aFpPqdqBqiB6i6oTBAetMJib3to4aGf6PAwjjtSHKG3ou8SHfcs/MA
Lufn82Zb2uOpHtMm44xEbKcKF9ZYhAGCx7KtDvCXxHOKdsbTOt0VjG2hgeMVFb5nj5XmnXiGubTQ
4XHZrV+Z2ja5yLyi+QKZr5/TssxO7txZe4gGM/2x/6SB7bsKUuK5L0t2sKqHdL31a1yqYSF0Tvmk
R8pdW66xBTuMnjzR1oEqGoZLIFFm0IiklDyuU65GnKYFtgMCvvYURlRLNVOjC34TcS4za5I6aldL
7+fEW7yHiEIUfASCewVX5opKV+mOFr08uWNE6EeKuNqaiSQvBXU51trHSCIo8KuwnOBkjx8d248Q
qeiXZxQdQ7PNR9Wx79gUGw+2wgt7wkWy9rWbtJIQttd4GxgckxXeklrDlSDgrrLbWy6B8nYy9o4M
Mb/5Yg1TNx9YpWD6AudTYzshE4vjaEp+xRXqDfgXVhgJXO6FozHGxewR5P0sLlkr56d33dPcmvgf
OSLzTbXiC65rr6yzCANDPjo8tWURpotmo+u/ol7g6BwqQRvubMkIFtGRGbEBcD0ldx7y2wg+L2nN
SKaujVWl0dBj1c0ikHOjWviK4WlcsiZChGLkluq9JGxUCnOI6CR2muxeM+gKe5wPZBLQvKixp8dL
L4UK6890dnOQWlwYu5uUrPaBE0e6dkHNCN5/dljYWGeZMWOcpQX3/wfK/6OWTm0SjEm3dNeFbBhj
Vq6cdoIkoJVmyHZbe6SD/yVcWLYsIlAcKLQ+cT438mLiC0aYJvyDsZyRZYtuPpYmxINvM2mnTRQC
5/BKTsi0r/j3kUPKzG06FJ3RJWt3SzREQPdrWZJ08r8CkUqxVCgz2PLX0hbrwkdyX3nYf5EgredD
jmct3wTSGyVV6bb0bMVnf6EGPUa4fYfbm2J+rDqpDt8fF+P+DAOP4SJCbHfnkzA7VlR4rejVh86U
LHo/KoETmpch24iedZuPCIFejcijXmpOXtJYcG23rWM/68j0FVtNi2fip3NSpMBpQE43gVcTBkPw
RsD46Q2JouEpmBKKiWjCPwmHwiYRAJwlrR5UjFmDaxeH4yGdc6ElfMCyXEar3yxXleyAolGE/4Vs
MqSNydI2IiOSLL9ttGCtnPripRB40YhRUZBVLCGhUrKPJxIbaY5guWBGwmafliilayQpjuKBhOm1
fJbxPI4dqztSUmMlBClTUIQruArv5y2Trja59o6j7wRrvpsqtYI79twhkZJqn/XYQxsatqTVUqJ4
mnXH5XvTdZkT/IHqrz+WIv6tUgxSXXhksK6uomuKBltMSvXRjzmXypwGPAxSOXcpt/RTIfPDJQ5E
VUjqMww1KODlO/p9b7Tvbft8IVuEf3RrNGM2LgZktbRrQ9Pbr1xK4hbAn8N9C6j+yWGLYxZFFxzV
zjztHuT3pu7wuMo4SdZU4ZyBUzCHkmm/Qg6/5G99EVgQoWUqkiBDQAdlgxyvkkDiysWLvk6xcd47
I97Rf/9it/Pv98oJReKEVc0pTvs1QQkwStt3tAn/T99OxbdaDdedUPZjxSRiPme7RxVA/mWdNTYX
U9jAmo+I8pq5Hilwh3v+qHMbFDqQSD++j5RF09PPW18VXkp0QcId4qaxONQf6gKIOxLQ+D+cgNUB
MHQAwRzDYSqYrOQact7YmYbXSniFk+nhvPxNcfUXmhoIq2l88RTY5N4hiJVZ7MHCuPDecDAHdPNq
Vo/bPepNS2tLURg/xDGsuyC1YJFrYANWcjcZ9MsRB7Sch5xHE41GtFmIRnXJj1LPvjPc0Zk6qu9/
HaadWoncKMjKvR3V4SW8D0i8ArjGSp+6zRpubCtZ9G7JiF2FG09f/tUMlvsL18HWna0HM5w+u8xA
+eVRnOfMCdPiU2D6EfGIqiWCFvj+f80RzMwwBINKePhd9UorColNmypTXkgUSy7vgSER07Zl1tzV
LWU8gKsS1X1Z8rum+/Rf3hkI/j6tgZaa/Ror1904/SzCB8EmofYkSbvX8zQ5QsvnoD8WHZGdBmTn
K2y5amVur/J7AY3urneVqdbsRZomDobXm+rlSKaDLP0vVWw7KuH7+p2P+4kmF5TLGuQPN5QjvlxP
sd/Ub7Qpb3R3VLxz42haBFRLk+Q7xFGUWxQK7Jgs+bDk2W9iPwUjbxKKEK7OjMotWw5xMiCMOKtb
6MREfDWVRASQZVJwKUu6pdtqO9RBiEHNaYqIhFu1Yw7NraLKUC/JVxKWZ328I3mi8NHy07x1OjDa
l6G42sPoB0AMXG/fVLRteirpt2LDW8kY0xp0xrXx3wrJzjVq+B3DGLtvVYlg7Cb+LLAU4Uva5qt8
+DoEs/cRg/q/xh0OzVmyShpxWXAs4HNkgXsXs2hKnGIEAVnUQkkhVspHOTDcn72RHByRhdH+Yb2B
L4M2CJ50dXBLzsjfBl6M0KJ77ZNodQ8pxgZ43IekjBSwHmgnsUkA5hsPZMO2iXNJ/j/X0qWyUT7F
oTIS3I4ngrCqEkf0UGsej6FnRkMq1BloKm/ugGJVvxBaBOpkTmLpHCI3X92RKMdJ2lOARPjrpSlU
fa6PNzdFZuoY9ATuud+xLvFo7VU2K0xqpQnDlYvftyWoZbE3djPu35I9FMd4ZufWpaPvIktF+cMW
/8+AsBlOx9tM1RzxNrxufpbvzFXg3/bx6v8yvynHTMl5lWN2fomaMdMUGqlZxqXo/+lUBhZFEkFX
MvvMY6Gh9dBvAJKHXYjPB47SSUbjHhBTzUqbr1B0TzscEDT1a/da61H7hbFkYjjpK6CZekDs4XQy
yffR0IRqT1iCG1ZuLjxswglFHaN2LBLoaEQN3DuB78MG0gvFs2J0ub3MJ9igmS9b0f2QC6mj9U+H
y5zePXJmmNgn4wLUdbI6dLRAcar2wgR8Xr1DGgyrrBHCQEXNxV/bmrydV67EQ/ZK+krmXiEyvBfu
ulGfo18cOZ30P28P7IkCYjEHJj/BG8JRYaXSGC+m+kqJMKCz6JOAUl/DR2k1MjjL2mROXmcuqXja
7XduOxbeHUANMhyKuamRBTWWBLnSsAVYKKCGpnu28ed/46ImoIvdwEsHyFKNwYmnfJMscx9koZhU
RiNss+PeMwNy1mbgGQ02jFEmmH/R2quoL5YAqwkWOFvP8OF1kW156kZSeu+FHz3F/R0E0jht0jBp
2+5gYJg4s/hXA/B4kHvLtu0WM96+K0CFyLMySq42hjrmqsEvSPB2q/AmJm1DdcwYrknf7F4b4hrN
9F6p3S9/4PtixDk80pWaOMTm+eJ90z1ZQVSNYkQ//HjBDVpf8geD6yITlRcShtPg+dhzl1MKinqA
5SXJwdTHhpf1hxkZh29uYuyCkeYWL53xJzu780rsm/vGu125cLU6DBaFWO6aj+IBBhfZTOUiTC0C
NOmP/2YxgZi6Nl5qqM8sMuHBUaBU1JayiSFPJZCei5lVmTXmFo8EuCbFZCZjH28XOXeviXi30V82
/0hRvy6NdhUYNnw2ll05FdMuJAdVZN5TgloNtQyjBuIinGHJ23+jGtfMgSHse8XycCCZCMb1ZS3/
TwTtA2PVd/GPC9mupOb/aU3oXz4sB149RUgoM7PzxMDgh9vQ/atCAXnhqAElW4yHm+qleB8D7EMl
Vg9N+FWr9Ig2U0Z4wgk++R9gxlJJs8M/Gg2qOPXPt6mDsuKX08UGA+ovPrioa9M7K96Yc5ylMHee
zSYgyADw8MHPApNMyxy+sBQ7HjpTlcPD8vjVkQa9DwflkltX6+RfhyDnRI1d1dmQNVwlyVkUdinb
gE1NrG6dwL1pIUo4DFO+qa1VivFd395RyRJKqQoLejrcEIdBq14QjNcKOghQSOKOa8jK7bX4eMne
sLnEpFfY81v9LfAjxshi76Ex+68R60olb6aUJbaeFumKhOUp/EFNA9SKIa6DoYlQPZQ4uH+aHI2+
p6HG5RUr7XDcqUv0yCGJXfDx62jm+e7427SU4KcYAsP997NlBeLT3AKoxoP4FVqcn4giB9PrmVGR
Bmc7+782+ZxkYvVkWWOtYkhu+PWXddXnl49QWqf2BcNKhQ88K2d2uikwyGYAzm9WLLe8NkOXyu+5
VnONQImOOmPr4Lv8rbXUJnHNhOOwF66Rpnb4g59/ritnX7hg4bvAmy/1llLEnUE5I8ySORiVyBoW
7wzzBhqOZIbKFvhv+4EcHOu8b4SNhyRNohPXSbfpMwMza6dRcryXE7ByPOhOKRI0XZRbFTZpuGlP
WwsNxZ9RwMd+0sHUaoD5GHfImoc4fEFw8uImvrwsKxK1AbCW48GYEWVUQ4NCrYXlOgOL9xB1cuXh
aEHIjEVYJZm0qXkFNKd1P858RL+OGFFRg/MynsHM530qFQVNaSnpliG82w63zCezehymGVU93jA9
Tl153IuHTNXZHPJZB02Guvc4etq9wmr88fPTmdJHtP5GMomfArXWYoiTls1STS/s7iO8uEb5agE3
C2uM5sMVz1hg+fnU9sdfQNNr41L8wSxpwiuWB19ci2yhxRmn7TglRrEVBfmCPB35aSeBMCjeANDG
RC6UXs3f3/o7MHIsyw+Dg+FIMBZAjzoaGfkSYI5yLkX8CDHyesA/QwucWcuqRnBYy+TFuyHKTmZY
ODzzgUek+AYRCxFHXVHAzAtDTEA5JO6wfUX0sGUXhIUqjFiUmVnB1W3LYOoKmADVQnc9VAUYrQEq
piH5wCLYqWY2UXdD8UW1IAwSvkI47JVTpGIgTcE/K/8pEh93LTekoXt9rAZ8iz/s0tr1CPHUqWF6
54/SejfhZg/miIA2NxzeBXz5k7LcHqkkqlfiofxYmKf56krmiqQEtHk2gD1svZ92oahipXFzHasJ
dEvmpo+ThARwLCVCz4CNnldCWxrHC+NqvQkfzT3knt5IQw5ST2+vIzHTtaL6P1ek16SFsR840CmN
PQggmJzn0f3y2gUSSe2wplBKljq89qhTNQbOx6faBIZ2fLAFj3uLoIERORFj5UqJrc0lNYky7Zov
lO7/3P0cd+d+K/lbFSFTAch3YUbANA0Hn4DJ2RZk9eRjkx2MgcVKdwcvsBZ85XnJhuWr3r7VSWeR
LLTnHONgYYWm6MJMNrYkZBNt0uuw1TIVhiFHNmwIBPXUu3kOFVZcTYy31ojz4NBSi8+jjHN/n+Uv
OQk+ly7Wsu6tVHpHfCsaJehw5LP5A7717ucCMSqQcldIf9ZcZ27rHFYHNgjtLSy+bxFDlZxzVmM0
33u/HpUPSH3R+ofEFazOybgojv2waJaPixcrA7Il9X+G7wRCx4oaosXqdHvR3UvmyJ/cg7Tzs9b1
Ys/PjgBs8muNPnNcWwyc+NkVShaKUgam0zNTYzUyRG2H6dUJlnA/ctQanYhT70aYjykmPpQeVDzc
jIVUe9mhBCdHSctqhz9GHmFamxkDbIHLKyDRuosNqxYTphaXP3iX1m7dOwWOLsJXQ6R+3QugxhjZ
Q4iAuXju3Kh1/lB+eZAA8NAy31yg0LvSedLjCsqXzwtxBvEzpaUt+8cjDcIYs+kN0lcRB8D7mTPO
MDwkfwqeq8H6XBCFifWa5N7QsIBhbfAWHpIr0u2u1JpOIboXCfpaSKVxdmZVaLhVdIoXsfyzjgjc
QClVzBjvb4FX4szp2w221WYdlT2DEeWaNX9klW9YCAWH21YnLAqRYhV6bpK51W3PpDccn93VF+sN
PoWFD+o8sFoICGjUY3IrGXRdr6cWEvWPBnOZj6onIseYjprRJ+zvVmI9onXAB03051OEeFxbeFUS
w/n1NNDlUDwRkSAVifE32uG1aIRd8Nr7pS9R0CKlJxEYgvn1Cin3WhbnqkQnFE87Qb96arxbE2KI
nxuvNYBwxgKwX4chC3KgnCVavZPzVoZbFFfnYpDj5lXJ67SEXP97xZogdto/BsuckQytEPxVNPHt
KCWTljEAAP2a2PwsAvLEADD4Y8r668/B4NK9gnVY5fIGgR6yljqol0M2tSLwOz28lprpXRdgoAaQ
BHn0G5A853nGvhUiSwoAPxM6mGe3MS9wODSklB6C7hX5RBpLEhg9t4bMfBd4AS1Boy1LrKmO/apf
A1A0Lp4l0L0LrLZxOJ4LE52jFYJsmiyYKWmoosiVrPGLcqPQea6BDosxCwdxOgfAyFBGChazdaoM
t8hvi8jC0980MXcSzvvcAStQtDcZYY+LL+Ln3802PNiEVftkdVmo6RnV5LvLC/WTQXND99AmgXMR
5BMgqsWgA4Guf2bw0g5BPzQuPgof0zCXmmwSI8kC8VDj+ycrcvwj/ll7SQrs3jizDBk1QURb+iz8
ccyYXcW0jWK0vdnfMp2jLqM+6mYDt/ha9YrB4XYrQYgpF9FyGTqG3hbKuJhqOFnEW91Qae2tbArE
R21alY/9pF6zG4/5zmYHIK6dMl4nFG/NwIapAGKNT5boGj/Sx0vkoXYRf085bS/hhy0WGq0GiHec
6UCi2gjO5OShEp9u1a22QosZKqUynstH/pbKqnEQfVaanTR0uNsjNnfO28zjwVyjHKBUH3MHwc8J
TcavOfYMfwbVTE2ecdxslfxLcFKiy3FFFicwKg3g+KoKjDhUfX+VbKJ00p6vieGMZ8eGYoQZ652h
m/FOP8///BOvzwwDQW5Na46PHhe4kd0jTG2X3TP9rzOEkUw00bv5N/7k3sf7E5CHky9yYOsBgSIA
fmquRbXtR3YdnO+gFxywLdITQFPKckEIg5Nt11v5x9zYNY/EmUgXLGwfudHyEY0LR91+8D+lenqj
e6PLMnlyRre4MLfwxXD0B3V0nEd7Ffxdu21HCUm1OZNiV/qdwCGQ3ffMtkBbVamJYHKiV2FnXarM
i3KDLFLLnGKDMmpDZDyzu2zucR0gwrY36zH/D59PwVmtFvjQD/uTV/H1oe0+XkYvp+4mYioRhAab
OMxbOPqAjv10fcbF2+J7VdNRCUvX/3PPxyq0gevFDVCnu/e5UP9/zSOtmccKJ0JQMKhYFfjqeL2S
9cpgYjl0g0CMqb3PmwSAoBSaJa3/f2FTFksyJWo6ILDhkbhUBDYv35+7vWHedulMXaVZEn55sEn0
n2lWzSFf21mOOsIUBX/gBa+2zm87vrpK/XA4P+NUx/+r7tGaF6GkoQbNiZoOGUAD6gc5HwqLTTVj
k8FuvBrLh8GnA5wfNGaDnkK9aAkD8y5pjYTDTSEXZD/IYQBhXKESSQy1Lb0MZ/5nYuQOcB7+aA1b
V0dhrkW66eY06DzYLa5GlOz0M/IxfPuiXFddr62GxFnUxO9PZqe8Dzo0H1Oa7zjCVXtm3a4xA5Z6
37+L0XxSH2UFINwSqxCK54lCITbYKz5lx7GRe50SH981n/Kh8kFW9cMPEerY4eRbutJzM6nJJ+f3
kLASFSvf4witEq9HlaCAsxFalQvFjnXFOWoXib7q10XU5WLBApk528lxwLWSKjI5Okm6yItjz84K
u9YQ3Hu7LVvbOsAIwT+CSrijSeG/AWFDqtWaq8TRx5WBniFBhm3GXeDWefSNktqbglG+x31bOaFu
xkwM0YosIZiDSiccXaKgjWdk7ozbLfdSO78l8uOvKGMVj4d+K7HWl0ZY8+7s1RQ31iak6qUX/6nN
bHeynsR+IBWa8d6OlUxNiUjgC0tLAjKDbgC9w1MDXg9CfKR5TSuKq/y9ERWcJ54WBvg/u434Bf0m
XbjMtsVK5D1iMHeK0UAVgPntgEvRO9li2XwKw1pg42uhS3o8lu1WHo6POKzhIH5FyAtIR4vpAlDu
fWJGuQ/nRYVRH3KIzpnuDMhk74VKyvUpbSeZP06Xg2ft6+FVlvqHUGzxk2UTbvELnJZQPl1nYSn0
hXGtLaQGK6TBdqam3+MKxKEOkvSWqfx/NkHYA2taoC4t+n0FhPP6qgPvpnGtKMvv6QmiDzxEHq+m
6o4w3KjHhZJU3CWpLaz8ZzoxBv/w7LEU/OdZrGv2me3H4mITRbwcKqBo/DcdPnmjhEdKX6scozle
biX5Vau+sxjm+Bg137yIRCQ9jKKfw+2FodktcEfYiepzm4vgMEBKTSEFB5D0yuS3/Y5E+e+ALi7o
mQH/Kwi1hNTFekTL58wHTcGenbZWguImwJSKYRxVDgteyGuXaegTpGndUwKGKrjLg7IrYSi87M/G
Y1wWlnxvFSC71BlWOrK/9jh4IbMoBJ2q4ys7kOuUYkXHxDtqwd6QQVZFWGBDSLIxEfw2K6LOmWAl
KL7gMoJHZSFhkLkqJYr+Zzeeo7vFdH5zotj8RpNBQu0yp8u3nocPeArnD6ROCjK7D5GUgYYauHBV
tYZkIChxeQ6COStF6u5OI528si92MGlBZ1EujZbD7bhL0tWXiC1MqtT8KjW3WwazlceKgeMoFDT9
CcNeh+x/H4lEgKyciZvM5x2DYmfiqojC8zyYEQkji1g2Kf8hnSQn2JqiZfQHESKzgAX4XSHp9+Hx
zW6bRoDizEiKZ1nsujldhopmIDte8IfSQMuMGA0ztF8nnXlMpYuElny2a87IvIsdPfpnHAlosiDl
H3bGI/HIFhYPiR/NUQu8+6ea7O0Ew1b5DiJSxdQDvGcBlX4AuAlfl4G+I5NaH+iJ3aPjPIzc1074
JsI3v/cwHX/d6TMS+2HahKH40O3bjvnRGHmoTASjEwkSJGR6cL0KcYtrU9PSy9TkT+Ln7+koILod
hxNtTiOiSAUGe2VqnvjUV2WZOdufGOGGIymSFVEOVws3rtYzZHq9OAKIcl+uODTS8dpRMGhWKKdA
00fHB+CnqTb6SDZ5ZBTOT8H4jELgU0WIOTjP59Rgt7rmoEZ655IvoMAyKIDXSI6ZROkTH2J19OUO
gVzFr1j+JIpQ+I5mZemgZE30bv1z1LdqqSafLJQhDsrX94Z+ju1x46I4iCByOeG9TgCVhbyXMUqn
msIDgih5OdMO0B/LgQiXPSgqaT+0BCZTlok+cWOgKoxulI3RiBatz1AvikkwcFl5UkEQTKYVF7io
wu0G98+vJ+Y31r+11M6GseHGPot/x16OcdhVJky1zlmZVtIvLc6f7EEug99n4LZhAFOIlDUPlp7p
hf399uLOZF/Ys9SErUegygadPkHZvgatG4LA6pmkQWDD1BmMyNLmVQiBGfNpZY/gzNyB/hcdADZc
d9+7ccS3nSnHP026Rjg0NNaJFPmhp6NG4zjXFfaT80dJ5jjAX3VVLzMz7HEdeNcVUZSH2W2xOLXj
XI+RdPLkmQPT16oM3qftyt7+16RAQadAtdE4l0no0PPuduo3U4bEwWsfylJ/fwZbL3LZkFPa54ay
LTr55nryHrWcPBKCNPJxKZTrfah/OFH766IVbw6yphkqsOrldU7RyIQ/+yVOZWq19jocsCswFkSs
qeGBHQeZFEAy3yFHGjJVnAvEOjJuoG3kuLHRQ6FlP++mquW7rAJyIcxSfq0v60SjCH1J61D9cZyC
agB8s/Oy93fivG7Qbl0083XVXvy+c3eujAKOgkUVqEi9bmypwW38SWgSwCos/gbKGU8FuzyMJXAF
O6lD6ahR4b7REWV8x0Tc5LFQfH8vM76AFSxpqmtbccDkllobK76FjPpi0Wv17TOu8SaKcHvW4+97
ygPpdfGcsPTQ77vxEZHVoUAx0+XHDUpr2yvMfNamZcVA7TtIqKaajaOnHQku0hkf0YTpelVFg+2V
xtC3h6J9yHNSmBAHe//XPITuMXxBBU4V3vGDLTjJOqYHX2xPPEuikL+UPNXC8XOSHy8yuC2BKD9S
i0iqaLzumOmbegfCe03EPiWl1YNNUH45Gkdiih36go2IJWgvsWdDcdlwQ7FK24WlE0whWi5wH0rY
5MjSZmQn8HLmpYlRRqP70PFKMJA+QZq9tegvOTFJDfBxA6OTOYGgFAF0k42zHi1bH2Ka3BCMpv7h
B+Lv9demNSIvgulSjJxVgJQKuSZ6eQdfp2pwu8pYn7OnfIufFeUlsgiJ/Z2ec4dGlJEmOrSkv+De
uELIW1RPzXZgSWWxatgPYugXrKghwfahfY5Cc89TCrixIQbMW7f4SuBrTksGsSoHO77i+s8yy16g
fenpGK9sW3Ahb/NTjdDYPuAyZCLSjH9SCebyf0eASLyl1SVFm5VEdD9yT+R7GzQgxmSkxji4P382
8SGK8UJaoPTMUXEmQZKSR6DelRndqnC6ACib5yrzv4zZPxCC/Mh97KOKZMXy2YbrvrRJLwuhnqz7
VQsugNSBjIfWWVzs5nebBpoZUw4BBByS0vX05WtD+PHaPIyBf2VJ8KzeEtukZI7GD8R0qAAHJVMo
gfFnZzL7hKlEys3FL2kwaYKYvVKZpTltn+lMu56O7ysdB68N5JcsSq2wjOq7O6SQCi8e+Ikmp5lY
mIsVIBTCPN224U4VIFDehJBgLgdDou3TP1TUNr9p0pIzPXyX5LeV5HNXfWHMZ5Xfs7t0hkuOKYIC
a0CD1PUEp2RAQqD5Bq4Ak+ChN9GKZ44rhIqtxu4kz/9HxvJIdtudaSQ2tewWacdlMUt7HSeZflMU
UysRY3Y9eH6J7AzV9gsdCkPHajZMyRePCBK75yA1UgDGScVGpjwVqiuhTd+tK+JaV7EHtT53PPqU
/wRMOtK3N+ZN3K68WtpnXAdaDbKvUNxNNfZXoo6KHzVtvIO4Qu2s8hJvd8EovT6feZ98VLA/i4H/
+FIDEgck/0IaJDnMqMQWp/MOHvYNl8l9+h4qPG6qndNdIAsFFMOy4Rvf/XMFwrJ5mLsxhCHbxseO
+Izarl1OLozgYKugp4k+bjOL2XFUaaWjAAO0auGbqs14r3J8poWyRhW2SSQnVJXoZr9KvwsHIcFV
p0gMjt1hXXb9v+3BNa431PZBdJZqGEOo4Jqx2d0w2soM1OT0tAgKz9XrdeYgMlmA/ljuEE5EpCo/
UNsPR0E5K1aEORj1PdjDr9VxhzD+4sxgNMAnpsoGgXk7307yFofaWOH6uaGWnPPNcD3fMtx9JjKg
9OTaDt+Xp1Z4phMdhCu4cAYZyEwMCARlzIrBQ7HAREdArUszWhzoMZmyF/Jb1CImUV6jcNNksiFy
lwlUkDJvCpJzF4/ch3D8iJrW0RV4K1KR2vZLT7hjpWdTJlmxQb06ewjvhbZOD+zpOSkJSIkD5AqB
mpcotDEmuLBlMdbiQbJtxVjLibsv5KUl4d27vRiTmb+Cldst/IePK/y783OMYsYB/Eevq4E5RMHd
isz9sAvmlhYqtXiuVxhhpN+T3UE0ds3v7AsyY3ackvgeJtiv5r+sxqCwj0o3mn6PZOliFJqqUJgY
8e0HM4lLf2T2DKBb6n+mOxrLN9Pbg6YAPcr7vuK7XnX8Y+5Nvw1oFEztI+f30CnWZXK2qGL7bR4l
bEat25FYmOoW536BTo/O6w4O4/MsommQNtVu+38iDzu0PLWwNKLk46fJbFcE5MOp0U0pXmzg0DLc
v3cx03RgWbLfXSdJbsQSceVq6kjqikXUgEnynpUgnrU3gZPltoaZ6b4XE+d9haxJC5E2uuPCNZ+t
c6XWHR5jL/UpnonxSXlmvx7cadKygu2uB/WUKOUjM+RKwzhl7owOS7SMdcCwaiZcgVfAvCOh0sKY
Jw4UMfz4fNfC08XjH2CH6FkurwjXyXxKWbbMzOXx73P/X2ghPmF9QV2rnCovJLLbdWmBKRqZfGZx
b/SPtGe/jY1UCfLs+FHYSFeK6vHbD4f7uccBp00t2u6m10ULpdweEzG7XjY26QspkoLiwu2OxCQh
xTqCxtmUxG4iPZxc4RM+H5MnN3SLPOlOtSJDWi/i6sR8GmN7iH2Av8YAGZszF0omctXFdSQbmOaw
eSQj6mpFl7d4SteasDm4ZS/JBxmOR160D+Urck3TDAXnN9E6p3LvIKGliMrMejKR6he9e4aDaVgN
Ny6bAOms/2YdJVxEtsuSfR4J/YZsMjOMmt1Z1DX0doixf9ZfaRkjKU79g+mCWihNQOrouDDzIgSp
lUa5zAT6xeoXuuPvd6hk3IEOlTbc8I/8vJE34seHtsZbHkAMAbLNc1+lJXZsdwHNwpAi2upRNWbM
PhHaGdCTkIlsyKuf2k/WckEKaj1We18W0LquiyHD9qW8xH3bVEi6Nna0/Nx0yWf5jSB3/FnUTQCI
e02U1dGQgdtUeopb6+d2HfJoFqVKY1gqjB6sIN4OfpBONjZWDGCUqxBwT7QfQtmZ2EQAdBG6lz86
2vx/C6Fsm+xEOfsKaLH3zqRbRb/DKW56XOdk7FiNcTjicCLlFlTu46mGOiGs+dBm3AYLd0XuN085
OXzmcpB1IbrGjwSgtT8vDEI41W9Kfvnn7XxB+UxKEez5ffhcqOT6IgRQD3MQlgP/uq5nxRXc1Hwg
1UHTTgGwPe7jkaKJZwtD/O9DueCIurLVUlZIZFD3RPCB1SA5/K78OTCF4OvadlNayaLIj+YIQ/p4
w4zEdjhYHVz4TVZ9iP/2w5pe3Y4ahLEwAipEEuO79egKEcfdwx4akBJ7C9MkXN63JPIMpI1l8L5n
r0RzL06ThppDLERh1u60mzXPU9wY18V/3nOtfcDKNHIOGNzGWf92NRgMA8KezFzaG5Yk4sLS+QMS
ho0tgLWFIS+LEkukelFGEI41WD3rL+9QxLhidv/J3HOVp/kLrzgsZEZu86557ovreuM4c/Ns9xWF
zfp7i/5JcycwhogbeUFmiWXSLLBaFvG5bHbeOCNts65jSDK0JUtkb27W3pA2bkcrhP3AQ4cgQhlN
NfI8XgoDZ5VgRmXKCBEQ4fB5ISLiDVcHqUFk5WuWjKH1DHkyQ6o+rAV6ZWC6mxhVvwCNTxTuerOO
7jqLqs53CSb1w1fMz70wmPxOkn4GVPl3fpvzR1nmYd/6HCWzDeSqmRGAjG76pvSvIWMWAVAHDGeZ
FpHHfjnONIykomPBLRdSfugIiO+bgs5VTLbLlGe3/LSs0UulYes1CvcB/qmZU880iFqUC6az+w2E
4eHvt0k7+6kQ9pNt/0Y6rrITyg+foY0ELKM75LZshYt0pUrr2GiASvx2kUX5mjvuzDpiFEsVhG86
qNXRZIco+GuYnQ4BRpQMOUTmwJRyu576jutqnhtXKa8Np4O/btL7DO45oxFeKFTUmF9+LcORSalb
tRWZPodKLqo9x6ocD+3pqRSJbblUjmJOEOldbALh6xatTUMRayv6Hb4a/MaB4hqyvad/IUbvNlaJ
rQZIMRkGVhcNMBy6YU3AHj74sooun8ZvdZvtmEEaHv08x61tgECyTwBpLefmXr+90/1/eMAl8KAS
4Pr0nvyVWauFFzrsoQqYddH2Vqml4wpY7RQBmYN34Zxy73er826c3+wUJumRBKBf5qWZSktHYENa
cx6e6YB+B4xDoDHWc6OoJnO1giAzMo7L5ozIUxF4mzJq9pvmTDxBfzoSsbNnE49fADb/UYtv/N64
zeStS0y/mCZ5ouaS+8PdOObezFschh4MlQTvKtJvssRxVSUYp2ZaQscO2+qzBOVw3bq0Mh3X+OmS
fib5YE0BTQb8EvdMccf09mx3Ktd4o2zBD36QFYA3TMlYW9kuMt9q3hIy9q6rcHEBNkQwnwlhpqsr
pagwCW1eDL+EYU1HYX+FF6funCJnEwFfCrLKABUfkUqAaO5++Q3mKqO8tQ8PchPkfux0nRHXG5lq
8O6r/9Jx0One5DHFixagShMfc2nU+NfAvuvtHXEP8xo4m1JaYlEHMMQePPX/WVqzolGeeHfkbOhW
5bHY46aggrvFB7Y2vQSvqomPuGuJm+WC17gsph6P/HIEnsshAZdt30cXvn+soM/vhLKBcKe3P3VL
/yBNxtszwXPh7QTNlNt57wMJHC4Gqx+dxSXMpS+jz9DO1VbFZn2qSDx3cKw5yeKY8Rgdqex8jA5K
675/DpG/SqXh7paBVO9G31jncoyk37hdQLN/nVyiGXea7myRiuoTHiPawstqo2MXw+b3+M30c9wX
Wij0GIO5NgnU558+UD8zv4GLJN1qIcqFGAgnc+CefDty8AasOjyfKpg7ShSZfp2uf9jwmgHd3BbY
eTPCt6lv2rhdtEmVOaEYDIikaRACKKa5PxN8sSRv8RZgmO0LiVlI+LGxWvNIR4rn/MaNfaZvT0wJ
Si96zIfw0EheP82J/ub90wN5w9rcaZX+7EtMahZepUX4s+KLi0VX9npETlNIzOfWdWkVwxfFsiAT
TMZtORN5jBIpckuHHDi95xZDBK2Aj5lF6ksGZvKSylxXst3pELCo4JAu0lYf3cqhPauxxxsuU3vC
Dbf81aWxtydfmAAVHsM+a/A0BbfuKD7US2vBgjylsLcnM6unu49VxpLJW52GFWRNkEdYuEXDOG55
jZESohRDFvtdTsR2EnYqrq0zItDP3+OMMaNZtxGysObN4weiJ8gxnIZy6JlDdVq74mdpF7Dqfe4b
PsRaM/GNB5tKqECIzmUQav0R625RfB4eyv0zq1fyJayz+sz5HdYwjvcxzlApe7zxnoO8imxfiXWv
Kvjbt20KrWNi8kv17TTN+6T6RZCGBPtlCCXPqYmAGtspmrTTUcHwNO801Tmu8mDui7h04eRyjP22
UfpuVBLBp7xI1avWVRQax4EIj6nsNR5Zx7Ax5JchQ0P9ASLWK5Jt78snPo0TavFIE2L9CITMA3B3
0UnZhLH2uTBSPspGG0dlHVpxBMIV5h79g7iodbj0Tmij9rNqg2izLHamrexgni7EXnzD65mhy7Oe
Fe2+5sMd5zfOyHzqe1nUkkLii9AeqqCi8YdsXdb5yEgptGSeKDQarsShYFMkezqgKqNvrfGpIVab
YRn6X6+9yVMmHxHbdRlirr0C85uX4LMlhPvC72khKvAFJfwb9s563scazAydZ7/zkdEcWcB0uOmk
kRmGH28xcBIe0EuX1TlnbuaTn5icl6DE25NvyvQAciRSSPoGpUfd6/etiBvNL4F91NZytrH1TdWx
WSfetnNyUQW0HwehcVi+KHNDG2TmMs98/xZfE6soAQo/ovJFsXlVHz167EdvSuEMKVOww7Avggys
gt3UB4LbBQkQ1lk5+1gOI2HyOJprm2jmjd7PiGnr3m6ffzKlkCqkQ7ljX2niEJyW8t6DWyYiwTxk
7wVZUcQpMmcedNCeb+zZ14XPKcs1yulSx6xqjETh8SdHetYd2t7B6dYbm7qPnw5bQ1K+butqBchq
UFakNBeYfGq0Og/hygm33hSv1qDwjW5xfmbourJmBNHNLMCr3uLG/mtYzMv8EOypj/H6nM4k/C01
B/60gjBv+LOmtm0UEPjgcNkJMpDXHgH2wTGWB/yZ1qxIP/IvJo7AfRGOdSRCd53W5G43T71oG8+N
L6c8M0QP56vMjcrJDtA1gXDBYXrerj98i/imV/Dh3ka2s15arJm8UVz5zqPXgpvjHMAW3ztbF/+e
SV0BGEShVpS3YcGOXyb93kJI+Ntv1Ma78B929Kz0GtcH3qynZ0ieqlLLoA3a9WJ+TbRGMOGasi/v
8txCmEed6sCj7ISgHt61WY7VFHjdiAPhbpEbiGoFTnrF5SCsh0yZhchSH2b2ox65+YrEsr+GplSx
d7cfCZF4CqqErbR8WX65/fnjc6QiHS+Tuc0CTkmgv2kCm0TBTxRzoCYNLYq9T9rlS+No/kAXEWJf
Ux3mmc+83YvNeL8ws/VRHA850yDBZ+9IbnPyQhh9ex5RfTru4Dr0tJ2c4GpYd0KC6tKBHF1RFoK3
t5yeBgOHI04extZkoOz9qBH8wU8OxxsHyKPo/0LJ/luQeLkY4m11cL1Fht4rTGsnFnVCoeT+NYjN
aleqBuLeXAN+4FaW5XyaVjg9ZlHXg9W5Hc9hLvlnuVGp9t54jXV7A3QECTszEkP3YvWpBjHbKMxr
I94wdS6IIu/wsVZDueDh9kfa9gjjF8lpZhNIXBfjiC9IddgKBuGF7orVZmM+Opnp+gmP0qI2Z6pu
/mzoIs+0xzzGLQYJXGMJbmXYCIK7wLtODM2mNQ6Ty83QvkEf8GiQrWgrAYff33Thqa198iRsoeeQ
iCGPhElqz/3PNNFL8X1K83BnozWwB5btvDdOBf9yFiZIBUq3TacyTW+RjXsNhhpWxUWVE7KphWke
pfyjkawnbg2DH0VjtF982QLLS+tvxtJBT/lJMyFd1oiey9DfEQ7oe2mlT+5wD/Qmohq+3rDjLp9r
K5FkjoG8mQ7HxEguQwZUy4EzqRngwtVXYzqTrdXwCayRBkWKLMif4uPGguSq5I9lTRLJ/1KHd1Qj
7BGvHaSC0wt+G52R2LjG/gDR5JqUVQ/gvxYg5ksB8Er3qC7eVIwBC1Or3GZaK3pAKDEF274Wzo77
2edvpRdJbG5hlVxMFzpYmEWxAHOiiSi3gdfEFUiDxcC4CCzFoGgmIoBKrD9Qe14gE9YLBd75LJSa
RWs0B0rQ+I0gPwMcfjef3f0iAWy7imBIWFp2kyrwcWF3JxHWKf1iONG3kkh4oamwgTXtYtTKEMM+
I6wSAJav9oK2C1mYK7QhwEn4IVv0j7DUd0KsswN3twlssvr+Z2O1v6DEjd7JzemeUAdC0IS9scdg
1bMRx4JO0gNznKFUY+JWvQeZ7M2SUP5YUHTM1vPKOJbBVuypHv2NdZpbul17+4caFzUDYkmDlTQQ
XlAcrBzST1AGYhd+509J/7evXMl7CRWJm8Unxc5oNHZxWUbaL8jttyF1IBCp/EuSdiTVZ9Z3pV9e
46acdcwu7zy39l9CFYO5yW70fX/qKi5vR8T+3kt0pCmSapvusdpYDRgIV+/Tee8YKzzOdPY4DwDH
CIwORtVz34tX6541OZ/qXW81hVpJU0L5cRqJROpV2ABTS0f5Vtps1TqhLBFmq/4vsfZ+68039vU2
KMRvOJanJ6XbxDJg2c69pTCvmtHHk+EB4jsG/3RX5v1DAaPJRIFcbVxV/k2wxEMNlTOxjfuYJ91z
rlNxOzkaNAPn6avkwkVPim5cZjcZ02HAPlWchKs+/bkWela0MbCUb3IWWhdn/nGoEaL2GdqEZ0NY
WVr8bQ6RrOQ7z0hHgrtzr8KG/vTcaxMnsekFVsz18KV2fk/W9j3kgS5QAaXjJAmDYSxDpT3R6O6V
Bb0O3SRf7OleZA+0oK0OfuMfe35y0eJu1cxtpnfdk5jg53RGNhXjSqbG3aX7YFEMN7vx3J3QXgbP
HxsChRGn9cZvHbiJBgebmDBrs9uqO2TX+ObRBQs0o7wWD+yiNgQd0SKT+ZZbZhhWz1UQmcb2HM6A
honTDQBDCUsLo2bAoo4OsJ+A8TOKXcn70tjVHzkjHy8tg9bIbWZE1gfCZQz1rJBWDCF6o27EcpBb
PPBmKOpjbaIFWxRGDfBWoz49foNm5i+gRmZtoL4G1PaqNEj8wOWObV2bRBk8SRL+60+NJLdL+cCT
U2sQgXgV7fz6J0PuTaIg8umPYDPCqq6Ay3XxxrLF+v3OEaP/iqUzjoLVgCi0WSn6Anm622Nua0Y3
LF4EBeZSG9HJyKBHQH/3DcylOlXNWPCYJYCWirbkBR+jw3GO/LCQ//89acktQ9sDRAQBCm5+kjDt
uPilfcZVXnwIaZ1MTOaBnWSVatt0Ivj1xHJir7ErOhr90BvBExI/QDMbWKEsfc73AaxOIzRdpVCI
fwvHddu9qYnVwLizWl+vwudrknFY1aFAB3S2JlmFs6LO2lpDwDb7iC67YhmTKDiKVGf3FCLcrbFb
hUJ1V/LQXN02RTPu13YJTlUcXaMKn6yI+NXFk7Ox+KYF1UrOV3+fHAa3k8AmT5Tyf/iDXWNLb3vg
BPNF4MhxVDVwu8pA4rCgGrAFeIdoWPg8/2Ly2au0TQRZKkREimIv7OSUwBdFAkcJHoaV0vcn1YAl
isWbXTO0P0qiYZwwnPUEM1dR10sw9EQ+zCf+jKoGXl3WP6sDCm2OhfDpeFrNgCllvI2A+/7b2pRC
h/mv8/rSB8gyuPEoJBO46UrA+NfMaJknxsSl/Ly5UfGF2KLB1L2mvAh4LY9sFTwae387Gee8r0Qr
kRDGiTr2gjzg0AV+qm6s4tedF5VZ1CwbkILgwlHPmBLFxhyDIEdLbXmtw6Xngg3amXGxtIMrUeuY
MfFbm7CK0dz3R9SdBQ3slMp9PftNKU4DzwApHTDnGkx6O6kWKh+WAHKBSHaSkMHn80RqUW4LB6Qn
ZoEu2DRR5/eEaRW6Z6ExH3+YzIw4b8+MTvAFYaod5D7SnX3WjiplP2r/c3hl89Bs0JkPKzz2EhQL
HRTSVbkgdVxclb4j7//gRv0+3e1s3BpSK5ydjrqqf6heUCdBtaIEtivYuogQwNIPQz4DG/ce0zjK
K2pfLwRriJclv61a7JTJr4nZc8elX9LN9DWkvdiD6ZBnDdm6M+qe3Pg3g7T7UAkGZ4JmPGhHoPrW
DvYGGgIX87lXpz9twUZ0lo6N+HkSd5PsCiQE7KkYb8sKXB4qKpVToODP9G0diRViaZZhtcl/2tDf
DRNt3/OW0gPkRNYMM3jXFyCnEk8Mai8CGxeK1A5B3E9FfUbwQI2UVu8UGFs8imhegazqtzibOBFN
ZLtP0WgnM3+/L8EZPcJ5OO+edZ/uULXlKbOlDnAmZt06rpc193jSsAUK7Ht62RssUCyTDqEl84zK
8sOyW6CTkhl0TYqMRxMS/dfDeASyTJDlB4XYSq778vv24AYztZwds7dO/sV49dh2Vqhj1AIwaPpZ
ISaMCGwKgb2IxZdmvgTqoe2CUCjrUtPOZycQD+ciNvzeTkYM7jmF0ktqIzw9X8/uYPnm86HLxkOA
EBWKYCEoQepw9fiXe2BeiTrdu5ul4uFyWGqhngTdBPwmwQLvD4JxpM/V3LXaaeGLKPlUfoUeeL3F
DqXVbB/CD7xpYASQ6qZdufZ+i7jEX+uGunF82FOiQa6j9+sRfDWYSO4YhX4qlzLEKVjc/PSTEhIk
FMZLRYYAzuvCS0VadGxAqTQbLBMHu0fJ34tWz0vqn9VS0v2qHkroOQKAj7eiPkTUmaLaOx+P8K6o
T4fr3rjFkdgHEooXv2ZANp7DP0w+CnCae6rs6bwU1Q6QO0ZnJ1Teun9g7lAJ6hsTCMzgMeCkvwYr
11Eb6G6kBRVgOD6TIF05i9dZSa1UrtD0hI2s9UODDhuUhd7aHn9b97e79IhbfcJKuGST7sFaO9e9
a7FsB6+7L+LkPebymBOf1B5RiYnt5ydaBWl9szRs8vgrObKSq5iJ3/j8bHumzcB/Ak8frEdy5RpE
D3fksxZpI2nLFCqReo3wX381xftonIwYQdd+MyzSvgmxxFxS04hXLi96adpsQXWsLJEPYQksgkdm
t8vLIp04oWIHShvMbx0B+pnppcaj2qoPKIOCAtlV7AKxt4m+wey8OLzfyu5T2Q5q9kxjAMwDSaxO
i1bbQTSjTm4Okb9YlHvYHtRtCCvrxj9KJ2PDnXKstKTzR5hQzS5NMNWS8JBJmH2vxFUftmjII4LM
ZvnDIic498J92WswgV1jS9dhe0rLfZ8OQv6msETy9EWSNww85nSkz1OfTVCaYHD35N2Tw2f9lLUN
lcmlAO7Rnj85KQi+D3uYUJpsmeL2AwaMA3q3TclGMZ4lrp8HVmj/4ev3Frby3MSeKNL8kCi+C5sh
gynjZfvACrtkL4afmEYVFkA0g+bxH1u3YM74zcUbSfDDtl3axhcHflzkgwuv/lldaJPKaxMC08g3
bO3z/SpyCrhvwyLkXPhCQg+Bd6J5zzu7DxT05HsZmF3HzKG5qYLqOSck3BECWA8qFJpeqG27PDs1
od7frNabjrAgDpd1QWDOPu6kE3Op/xz8Djuoahbmk9AJ1AoY/AuskhWZRjXMwE6Z0kNQnllVhl3X
jEmAIuHYREeYhTVVB3QCd5UiVOeRMInB7sVwLkWAr+bSpy5GBDUjj/zhwF3AKU+nHG1/EjGOMJk5
dXZ1oDEfiM2+4evPHJ4glwflkOXULhkgxNAJ9A0vkieZlaHDfy1CdYNXhkkiYtwXntHs3pg6hqFQ
j3KaTD5elUrjSBwuY23UMB81k9eXFmlALAImfB/jG56UWTlOYiZbnb8qM6LEbzz5Mm+0xvyAjjpf
faUeAkshkVB/0TJBHCY64rhL3a6l/i6uWe6/DAmvOtrA2zsGJS64hJ5nfrMkKz5e6tCKKZ17Z/ev
PNsMigDh0hMckaWwZsv++7ApQLP0vRxvlsQY6bS9H6q97zlaq4PZagw6rJyCyyXSEWjvVLman876
siloJq1hvgbaWlF1mbj+DzqtYrQ7TZ3kHezZEyQ2EF41VrnOF9vJr7sf1Yf3NLWKOv6EHUymjd2O
ZEslHkOJKf2GPa1abo0Eu7efS8iMI0Rr1/2+r+Ni5VwLYrJA4vd77BUZmbaVBRRgfQ5sKTzWSmLX
cvK83fcNQWZpzU/CC7SBGmIo4P4xZp28E02Odu5l+bX+56OTGScDy/VpcVJEbP3CO/y3Us1b55D5
lGsOanUZwZEd+Amz/d/wBoXtGDu8moyeIqZHpku2MFTAXPdUqEklXKa96mIJzjHf2kqNen1eYCIo
xsOqMNCdwLRaRAYKQ49mE3kfaN8DDJT8jbEZOTtFDogWUPJJ4xFk8fdAxexv8huLvIG2q4YeEKjz
jMlv0D058FjP1UX9g0beRLQuQlSLT2apBRj8m16Ut3A8OAL9u7JTQ0Bpz8AUsZAt5rJzJ0/kicQQ
i8lSp7bftl8DIffLvFZwBmoOFr3gSSHNB1BdupYuGX4abOb4GXKEBIs9BV815lm8dK4IuCVZwlyQ
URKR5GcKkApbI5zk1UCH/WKqvl0Qe3a29EnhCKHhPoCFdBdqkZ+ghVyqKg+5bpNWK3USnbVIZe67
79X1FEWdiIN3ZwVDeE/9WynOEPoY1ud9euP/ONsoMOlYG/Iz84s6rwge9LcY1QQFDPWCdwh1Nlsa
xTTG1QCKctnVuWy04LCnRZ+35PYtm/yw5vBnD56DIdKhizm28ITIj6vUY3WW0g8nlQQfFgvWyq/2
IOEDrfAQpO5mWvB+HLcTsuTbmqnARnlSgklRcR4h0p03lDLqUxpfJvzb0yR4/GeCGA3hRe7STreS
KBfS0qhaZOuQuURdy5g3Db8qpBbujhG2p+w4I+46qYAYayw7dOT+uSHlLIgs6bQZ7N/1dwElVcSb
cl2pLrmttHYM/tD8tDYR5XCuLDASWMFFvIPqMoVuS8EyqZD8WP4BNz2u/kfTDIS8IOp9MgSpn4Kx
mz+L9svLDl7BOHGzgHYFO4/7c8EeSogxGsRQ37LqAI5cmLHdiaJLgUjxhPVvrJcltUWySDbnWTYj
fzV7itanbtvZfEVYjsNU3v0G+F9jHvCKW2Zjh5z39yZx7iMFpLjHo1/MV1Mbned8Tl9oHTMjIj/d
shvY9puXT8VlXgd9Nrxv8yRfR7MWSo8kpEPlT0IvxXRmDEFRe8TS7cxvVEhuaGulUX5uO+7YadJX
ovrv/GrOCCDtcRzmj62RIhARlITQQE4YvGcLSA/pFaWDvSgN5GFXzF3Zm18vGtNdLzLHFKE+WrSv
2bWx9hhXkfQYkUP9yatRXCDMB4EptDicO+vHf3ES4HSDALDx8iK/PUMQBwOS+lBEeVDCFszeIP4G
0nN9RwxmDkKyxQsVn/j1Nl0cZnOvZzw8QQM3d+3+HvhUVveH40Gkw+nyhXTWfEqtIt8+qPhTob9r
3qYKfbmhMtjDGIii+npME39toxyuYwKuVI8WjXNJTXWwREnuJYz6HljxLLkg1/WT7evQzTFphndU
rv7LQyLKfnimBIahl5/hoRjYPo3j41W+KLsOgQyKEDKw/efPpD3lEenR0HqRaQgGk5Ozeou7qmz/
6MwydbBVXxQyL1mkRxV9sq2QpKSLIbot0GNOhpsujpUnGyTaJCjfCqU/Ahc+HOvBEYagWu0VXZVm
sBav5fWf3XMZLI8lPtzSjjOt69/z1FH5ETbUs4FHXO7kdjPk7CyUffW5fXaWqqeiW4sI0Yofup9f
PRIjOQMaZGbp3tm91d6UPW6IihfdNwKOKMogwK0pq8GjMw6K8UQycWTIvLKFY+G838ko7/a7+WaN
oMkIgoMsOhyHsCMm4XtXOZOywBBnF2kdyJEQnNJtdbd11RUxFi8L/rdWpTOwmcVvKd8UBjm5KmCz
41aV/XaacxSQ7BvlcsTls2KBG/7n9m8f6nLbR6UuKdNaEeBf3Us3F0d6EzO3Em2maNRlprbQPynD
zkYUcl8vV3C4NH7SwnUM+Jjjc7WdB/2dxAsvrClpkvGXEzgobnpqlN/3YEaMvAVNxA9icASrgLIj
t4/8egxQpapkTjs1J3HXF+AHjpbUp2vgo5c/8VB5NCErkqhcVofAWOW4diEpbtiPq7l+h6t3eUVc
FxT0RcZ+ZZy7JavotY3Rukh8EtydbKtYOhXGGFPX5ycaxvQQIijchJ1BJR++2x73GfaFSwRC/gq2
8c2msU5iXv+Cib8UuR6mdd2WxmrRZetRfSUcV0LvZIllOePZULwXE4/qJtHFmX78jrUQEtskEpag
UaluKnG2EnjsFqekIFUBG66h8JoInV0ai8zf+cMAPDNxwN/KdBx4+cBmOcZko9n3C3jeR26kjr+o
SVDu9XqQgsk5ovvBPgWsqjCfYAiUR4Ihx3ZP6W9TEtO3DjQLe3l7K8q7nQkYRZcZAyPD72x4tVrU
oSp52B/C1/qQcArJYt+saVJZbEzT3ARa4S9ER1+BCFDACJ0WlZ7LeJZTel1AchIjA3UdDIjGRWvt
EDK/b0RjN9TgcXbt6jX2Jgzk/tw0sYTLlCAYFMWXkqikHra08JlceE2n83JlpolvjpehnieCw4cR
7CDVWyG5QKvkpw4v82akzbiDum6oBnTJXtCfEKZMxXdRzQJo1Yv9aNu3IayP6PzOLRNFqHZ36KM2
FCIMKAO3CZaiwU+2Nbzmbc0yVmLtToMsTC6Zfr/S9XWGQjik/uHRE17eDEgK65N/PyyzOF7alwil
TshNv2tIgzC7nX3ztXTg/z3UBkwJv2UOnni+LM7tLdH48B7vc035YcVfL3HWLS6coJYBZTWb6iCT
I7jYoeiEcU7W06m6500tOSLdek7QtIbgLeFZE4NECb04uGfMGhzP5n8z/d5WmpOM1ZIQRG1maQCH
VCw+Fktqwn/T5DgVbtc6hDxxlIqQE4E53qHqODOtfGv9ra/EFATU/4t0acTwcmPNQtgki5zEs5un
geZ52kStwGrUSKxxz2lQwiOKpDic7ouuIdEJKOlUOuGMaKVHg6Yz/fIo8euUbljMFisTD1irB/GX
CpB7d7fZcJjxK98LlrloKDLeTLSaKLtGsuz5mxf95gBRzCNc3+Gpaxwkyv07UEUQrkN/czbdL50T
uyKY/AKVBNQ4aU3HBOzHiarXea5aKRravVs9mj3TAz2CO+mizo43NgYMb9fs/A5cY4ojrKTMpDyL
op8wDATC9EdVX4Npfq+HpsAgz44+jPY/BQZDnIlhpY9gSjpVY/V+dXalRJKtpPy/8b0VGU+7hVTS
mXQhOxHeXU6TRghWoIj+JMqwmUxGc4v7snODUuc+HkS/Kovztxah7QWnTcRrj50EUyyrqkf8RJuU
CJPP0O/zJGTaZQMiAKzQQWd7ZiG8SieAElHpQsKIEJhafSDhfBz5n43lgJTg0zoyQQWmvghIZWQf
57xgwiBXJ7mJeGa++xQTdfHb1BVYwiYfVYUJjfEYbhD2CQGH8n4MbNhXY+RXsLSDJaedaS4NQA8g
YGfJ9jG65xw3IrA6jraueSpNdKLGMgpqfdy8tG6djA/CuaO/m9dLQr8ysFxwkzu2Nn53SSu88lUh
8tQJatTDamGEBdCr3N/NK6S54Ye28v4H/rfX3fBtVkIQnm75pU7dWweuMNoYIwol2G57i5VP8Y84
3DFICs19f6Z7LOjt1HZy6E4Djck0D4tlxDtl64+Zfu5kH5jvsEBuK1zCoGXyEOLKhmOtGk7bWtlW
1QspsRxKOaAkzAJzYifnIg0wOQC4b0sqv4Owc9ol6Af+PTymWq3CVGROFeJKq8gC2uBbuVuijdo3
Q21minFA6+nu2868dUSiujZGTSfPqRz3D3NYCsL0p+LlYyl1RRo395vTnzrJqY4bxjprZnEe3oUh
D4Jk2Vllnix753x2vCk9pxEP8TXIv69o3kO/H4JgaK7X7/wkND/Xd4Ine947NLdLFgMxiIKmTYDH
AH1cUfjtMPr3hSnJYhpfthdaBp8YJHg6DQJG8umYXV08mhJIRade9fq8z1OCNFks8fR1xZPmfPHs
ux77G6ALHY5PtiW8qI3FrTdWcmYIRZlXr93vyX8GzVgv5xUrwZobhCZKapB8PKrxKoywelMCnYK9
l0nWz53iSU49ZmTsguspCnRB5Q6HZOO2zoObol4B6uPK5474jzJinp0L/TqM3gBxbebkvNFb5osC
4Fg90o+XkLihSm8mnEXTVzyOHxsU1w2dp5xfbXn4nvrD59f+Y449Ao/302plHTA7tE8Qri3tmP5K
/CVRIwlzvDi8BioZy8Y2qmxuHyJ92+QPPM0NJLbR7BfqDQaymVBnG/MPa+4gBqcf8CC3hopPsbe6
AESSh7jkxX5diQZA51cOHwCG7YsyQ3psQ/JaUfSSq+5vQ4UtosKbObsPrKW6Bb4IbdnQtxeR80CY
vR2p9OjCWVSHxzNYevZoY9H/RmLD1AOaA4ANOGWMzY5zD5Qa3K28DTJ0iMZjX/5Lj2JrWvfn+Xe6
NubZYz/KibRO9u/nJH+nPVT8tI8PkcZVFbPbgDKMDX8DbL334jENRhJDbmfzrWJF2ILQxAd9YDhX
L/A8zOx2uxBfDIQN0p2MJu8dICp9R4ZrkIPkH3mZWXMtakEvslPCuEgHbvTWgyMLWeRXtiNIihsP
fsh/pVApWwlkqDjTtConiCWumSzfvQMl6mSvALiDfbMOdBCaPRBdNlVHsH8XkJUsn3GxcVe8wtAL
K6a8ASwp7AV8OkRMYOJPW+7+NrS2HrZ8K9/nRrTN6x1qj5Madj+WGwjb9fNH+4yU0yY4SIHOllVY
R7vLuj/XGVg+cSyli5hP4Xq6KTVglLtQmsn4A6NkEJMt8DlJFl9jGG1EGm/6oI7QPJXfyGi9qWIa
dFSaQumICNR8dolp43/PXYtCj+uhyHDp9W6CiXqW1WsQheCL+GB0mRE18wjArl07Qn4Js/ukDhj+
Lw8VDOQNJQxCSskm+8SPTqVArN7pM0q5OERjgJGCf+1fJAEdI8j48LMrRWpDUTRRQNzIj8RH9fkF
y3XRVR3MuxYDE92VBuCijkbWW/qMq444zShuLt1bCITvHgGiZf2ODPQqnYQx21wtq2XTK9IZV91e
/GaGzwQPGtuhYoz+VilbgAI9A9Aujzs/tWtFFOd8GlqkLnd+1AVEHdivVT1MjcMal7Q67M/QUksZ
0Cx+C3/kTgIcXfntFO4bvIjCWfT1wL13t2rzdLr17QQ1Ls8faoorUH8f1SbM15IFkvWtMZyZho6c
m3xP5OHYeACGHgoYM3ij6MUXj6w2DZVjGxy2owBifMldIy3/NcLeYCv+e3SHPhOOBcGMi5NeYh3S
5tmiQVoPpStZcxJPiBtBvk5u/Iop6jXqc5Ocn9g1t0IaO6xYcVCBtXVMmlBGODRADKpzM36FjoKq
tU7X6Z7l9tqu/5jjvWWkqh/GVqzGR3R9ySm6ExgnNi9/Vf/wgIK1MI3zVeIL9lQVs/mCH6Ej3Rya
Sbzr2rGr24KJMBiVuylvueMk/9eJXhVVHjVYNPlOBIeu3TUh9hLn2jO2fQiKraANzYk/hisX1D3g
rUoGzqCfMqsczd5DkexbTVs8UcEFrZ2ACMP7JfeVc+V86BOdq9KGRf3u5hxRJMRvfdi4Ip63wSah
WtOfDIGvqJeXRe5dCeBkzgwDxU4BbYzs5Mc5kVqdjaj07x3ftNQ0Oxo3L4BlepWF+xloUg5ZSoD2
i0/Tdc40Xr2tToSMIEO9c1zkQsxzW7M5jzEYjRbgcqZ3+vUZOpcC1nRCcSLw37D2hppggiocysig
4f+XU2kEVlHZZ2AmlwbHo+Ktch2rt9q/8PXSevyB2DPhLbHEYNamFC2kHBiYzQXNCK53dd8wNKF0
54VDIGA3dYeVKqmHwbUYwDK7qUGmKtM9u2ZIjj3Z6CqN5V9jcy7Utir6ICboKcSQZWU4jYoxYE+c
jKpD6C9LTVxo3rLCmeWGbHzkN5f6LJwfh5H7ZgnzwHHoDu+M2oEVehWtqyEZU/4xSMd9ZVLVbk+O
4DRYjVBH8nprIHtciBD0yLJVT4O97XqBxca40K3wVVkE3GD/8gopo0Y2+y/0UUQ1soE/WH8A4qdF
OzHNagXnxxde4tCbD2f4pgZVUS+BPL0UkGCqZ/1MzFAVw+DeyFyvgnHgvGKf/LdOFOvarSHCknTX
AxEhXyLKmKbKo+9Qanr6bWji5rNugEc3NF9tLm0bpCBlxSBHJy88dJ5BftXaf8x0rbEDqIQ1LUOg
tX0QEwBtEXH1k8ol8dn7ago2R+af7vvtGl9LNnRw5+JJJR71cGLw/5fOyObBSFUEmlxNNIWR2Oyd
QKT2SeTRv+bn7FXDJeApJ0lThDIceJuDhSiPAEuMudeV9QbbBk3aUIKUDliFOL8FdsPEvCig88hU
u/7wR8MkdMZ0psX2j+mkXt3m0xvyNnZvvlOBvlHOpmaSkqd4ZQdIiwNq/+V3GHBIpMMhqF4tCTL/
R2RXjxFKn7djrF67XHrZcNkWaVBJMdyyLBDsac5i85QLfJXOtXDkJVw/rkGmkMW3gSUkK7BeaZKL
qkF8IR1KZYJhGHaOip+3zpzqnBw9h3HMY+kunGpmLpb9fWZSgKBNtpNFtKQDCv9rFzTRvMrl62s5
w6VIlEHDqetuALPuylIj1Cdr+r7/egFtTbUROKKnGj1sE/9C+95RIwd4d1vakOjhZ9XHv083naaY
VNv4vznLC27yTZGGlTsrHv44Z4ChPIu7R5kRsJnJLtuiIJMfUH8KkJgCrBjiniNpvp//WHCCDpN5
qqx4CwtmMcZVmLXy/BVzl0rBz+o9Ug/y3RjwQh8qy4Esj8HT1WyJ4HXmgvwylPYvDge1vCScIsg3
mn351mk+4Oj8jlxRoWyX2waIPqr6WA+O0k6diXpp3MHh6RZNvPBl9H589diVUZzKNOrL/gOcFtGA
0Jtv/ulzVcFpXF0zzd8OwvBfPmPiMoK3Wgei1as6nOfP0RqDqPewtTH5vxlRsbg4yudzjnKdL7il
d7hCCCx34PHjVM+WK0t8c7ilScK6cn0ivsKO1WTNHbwS/X2ijI35keG56TcoQwwPWs/8qwirIQLu
iSdMLVmjuVoznVRxPVJkpIVmQL9lkitiXJVuF5wYolVrCqyp5mbaCZQXN9gYnC/633Uk92g4tRdM
Db3rc4UY55AkVeWEzttViBi4TNlDSds4fBr8enrURj/RXyzp7qhVyMdqr8PWgJ870xX13qKNtYqm
kuZAmp9AOYLOzuRN0aGVGpVDDQbkBk+I/N32fjVDzVOTIABc87NN5N3c75gtlKgRopj7jiWoPT8U
IzhI7JhZra62olIdJfFCN0bsb1VFaqhj9mbpunwIpdw+5oBz1RmUChleytk+re0wdMB5LTJtG5P8
TWMXZYWT8Zjkrygp2fklA3j2PSgTSpNw2ienwMh2h1QCFu/RJ6IpL7lrq7IExw90rgMWcTiUjaKL
0o+57B9HWFdX83HWymTSAIc3brghUvGMRuRW7JHY1OFmPtHP6eK67FZPZxQSBewqfXpvFzrCO4fA
XymrqXTnkqQ3QmNTJRD13yppsYeadCXRN7xwTwvbFZY7kZJxj4JMxxSC2nzhrJ734F/tZtrJaeqj
uH5CFnPFEU6gwWAGDRA47e+02EiZoeGWKB9G8vOUW1NfB5LXlqH1YVqjWLjd/YOJcgcHJjzqDF9W
i6JbNUSTY+UgRSkol+NKxf55pm+vKmogoGElR7MU5ppVjayBnNy14RcCBTJLay2nwsZiV6blB8kC
QjadB8/gpS48pzfYPGcv3Tw8iRSVtq24IqtZKnhDjTEQZLRfBiH0NP0i0ohVev2M5MdTWu3Ryrtl
djsNBq8BCBGeb3Q5o/+wDPH0qTPVBAqTZQtOvnwh2/NtoQEPMgZoh7D9KG9/sU1GkxDmbpl4g3iW
UutCrEpVFhw5mlQrXAzgETYqQPHyM4kVIrLsW/OcSOn3kcjIPAcj3O+LNO5jfm3KZO56G33fd233
/TxaRFn7wiCuV0wwyFv6g1CgyIILaSqJtMWwZz50SLRdeGEbGKQUIxuZDtARakReFaOewtVG1pBl
v37IHJNkUPpanDTEU8ZolNnfDtRBAZkx8qcdPGRIuqvIajdcl6jqO5rGPqIxSW9waA0hRXIfWBqX
GLpdx8ZPTtwQkUjMuDUIIQI9L0MV+IrIFWscSE/uh0nD084HYvWdVKiAwB2jYJpgrvgBoBxlCdSk
J69CTiuraQcqdb0KTgMMPZVIug/g4DKdUrgit2RL1Mf926lPUbd1LeRLD3HFIvRo27Tzah6BPtQ/
HHzS0OB6h7wnGc2avgVgja7bu6W0tJAIsSlVuOhlpUKy2PWwn7q/eH9PmyS2GS0bFxA8eUO8G5mJ
mlP5sFXZkKreatHo9g2Ge0AA4WpnKy00UGhNS2+0FsGH96EojdssoXLHBwneFJvgkFB7mazrJBgQ
ORKL/AWm/bA/bM/+Flpgf01YtA/s6FFpwFR/a0Ta4x/Dg3Nmehhp/A3/5kp70Mr/DiE3qguNmgpq
ozo9GvRAK3j3whcg+pQUOWQ1QLNGohtnKrxW9uMjArNHtPyOS6bZCqedof6J3eSf7XHQEwW9/6SN
/tULz8yougRoDRoRxXXHJmpJuDaOU/yQ3HnX4fu2S2BD8dCvZgOB5BkqAjZMNTrBUqQUp3/AUiu4
AEGVI1rhSjolzYk55PUZTQHOuwJGq2TaXwc/WmyYS/x8mfmG/5K1lNfqcrTfgjIGEYZVfMs8Pwzm
p0MM1isVqWcUVrEvbQlmpKhnUj/LQ7zWhbsR8nOXXaLSc92m04SI1IYAs/NttQrV8LLR43aUTsmO
4qbOLhVPm33EuG7x4ZwawPt8nYXzUz2yGdj/hX6UPs7mQW2JjzlAR0vHspx+Y7wLA7O33yF4zZCx
f7LW9C2bEGqd9ep8beSU3Rn6IUZd8JbkZqZwSvYBvfZp5GaqAZVCAL8e5cCuc4N+24Q79j2+2199
nszvpEPpSdmrJloL+CHAQEzbNVmNWpnp5HZrcgUKnbOweLDGS1Jxj4n2DVjyXtYxRAJYqHg0p6tx
j7CDGlk0L1j/EwUM4xEDE0xRvxk3LRz3x4uKIRcDjnQtn9FLU/AqWhkgw+aCSHi/Ib70N9ZCABg/
/jFzcT7K/QK8EmeAefmsGcvQldwRJbj0JgNb7RwL04xiAB0JS5GJkM4dbCq9XtQr/cL2GasTqPuM
hQsGf7W4RulPYP5nzwbTBVqJbLPpn05GFHWPw/qBnvaOKRVpgqYD8CyqIZ7wtLHGZo4q5VbYphq5
hfJflWnh/brzfPydr4t3V+8yCIuXJgaeZSxWJJwUempcxcBA7zWteFmX8AN0f1RcZ8/w3m4yyffc
femkKjy52V8e0Avve/j/1BO6Zcs7xHJWrrkY7VoJdwa+mddMtn0D8smJDceeWryv4lGRNawd9pJ4
H1GpqJXehxMo4v1ZYVvOxIZYDaznh/nQeClG5zdG6oVBrBpxgXvkiF9Gn5nX7+TFl6AaJAjZowAW
oWEZjA7VdC2kNZwmMDj6svcDwyzsZ+7Hpfa/ij8S7lQ6c/CzqhsqsM8v0X/2wVRAa27z0eVGlN1i
uFFkqKxi3myyI8B+WZEhUyX8OVYoFQNOdIfnTRfedFeWGtc0zoffx7ZjaYzmAUXvwBb+pTuhT6aw
xSAAmfMnB2jdPEqIhDqDC5ukcVXJ+Lb+RBxDW6Jo8idSebEMGMNxwaHSS7bK6jNSHibFRmHZkPey
R+nOkbVctEIuS71imMYoF8h0NCM9C2w7EC5m51XFi6ZNNIFmDImOwWZCLDPXBvpMukFAdNHDLDMm
T4ofq3YdwejgHXUCawsp2MuahZqhC5UnMGTfUemaIr0DoBGyIGX0UhwyV+wMu9zZCKXrgmzTk/WG
x1NhmOEamvFh4+lPwiaDuImmCbPQuoe0JNpmychuvNH2j0j52WSngRv7YfJBPw40ZGm427Dkyzbi
J0tb/1AzGlTgmeuAIvl8IuQZAjt7guo7autF+k4FOd1V82WZ6atM2p1Yfb/kU7A+6dIvI5bdlHSq
AK7UJMlycBOs1yPmTCSip/kQkktGMk1F1aA5BCjuiLZNkeHTd4j88tpqxXaFYBGqj65N/iFk7ugS
oKPEkyj/+UyFk9qCYoXacsByBCmdbi6derz5nBylFnhVQaTSd3LR6b74CE+zoWAqj6/W21W/8WwX
NefzE7T+lruKw0fIZKzK5add9rmfVr8XlwEwYfOpNUF3mqBPIDD9g97tCQFLU/tM4orBPwkAjTR1
bXgr9zmr1DdtwmChNjdUqmiyXMa0j/iiGD5J90AMhpM75VkSCmcF5lexo13XO0+y0HRO9TQShczx
JSjm/wGdqbS7BvgC+Qi+9Y2yD/qKlv8W+tnxk/pD0meG3o8ZCKjIINi1z7VzIVuQNQ/sVW3/viOK
xxxqUkld8uI+FSaLEUwzwYe/H8kc0wN7xh0iY0TYww4HNaUKKi9zMKq7UID2pRWu9TngAIjwP9PN
iNOmEOOi4t3CGqMGAEY9hDAuSEdpJOIZUFlj3S2RLKwagLiBxsQRVbw6GPn10TUTmZcXnQlxCqhj
+OnnlEhyNxh0mJU2GF1R/2kZx3nKb586zITLWRSFfgCNFOGsS+JSEpebnhfJmExwN4JgPJ8urmkL
iWO1jiQ2qiIPmPa6K5RaMhWektAVA6MSr35sEJzY5QaEprimkgK0fjL9KPuuW1uOKDtM2vkUSTc7
YfOwQ30GHuAHOZomZYKIflEoaKw097CW9v88fWVrSMGgQyyuPGLuWzZlsOMMmgkKWaPseN7f75ar
xZLOCWm7kw8RU5kSElpZX7GnBtU+3qCf2GXixQyFizkiZVjVHe6NvBbSrDi89zE0wvHa6EA1oi9j
93zQdPSe0wNYm/0Ne5NRa8KMuXTe/XNJlI4mx2wnJNcsbespvRtLwvOUwLL/71SV42YWdLam2JB4
/Lb8gQcdnmaaQqK+uP+l7TpEI6FtQEAajpLYsyuDdBRZ4kN90FOfP+rscQ/GRv72gAEFgI/8ScpV
QNX7EoUsmlbWDo1KSI0hV6NiCiDlu1jfXUL2rtO31CPQxM03aDaek5FdlvR4Vh/Ca3ZRdF2w8CtL
qEAxC8vbF8QfjPZrPxTV5URAaeYXx5LGnuCQAphxqRh8vA5SQqWzKtEgIyX45Qvk8ivpfs2RtZxg
fDVLXrZ6Xil607j4Ck47Twzu7GjrFJzK6cqj649/qfoy0n9dgB61bSPz/r2xUxubScKuYYVf9jYP
Gb9ZxU7T03Vqx0GNv6Hh07X26Wwjvwg+gERQqoQENd9hhA126VdAD8x7sR93jdvV9IldO5t0I9wJ
cWMzh1oA6HBPEj+xs5bkI+yALDRdsZ5JidEr3ck/g6SBajAcdqdupzBCf7CX8KEcWRuIr/LIe2az
T7/GFxHGTf53Q0iY4zhcdiMIXT8fLBMiAfsbnWY9fMUWVz2psnEZc6/xm9p9c7AzKWIlFzccijjJ
H7ENxirW2UISQKK8AhoC5h3M0PNk9aaV8yVlHiWp5HS9CFdJDRX73vm3nEAIq9rCtFq7x2qpGL8q
P5F/T2t4nAyv9yqfTut5mfrQgL2bpu96s/QimA9klyEMlkU2XPwiGOywY9AXsqY7wCNSCg0kjzHh
qDEzyRNpRyqCHTuRkgwzAZsP1S2rMtHsajb5TXm9CZWD+74nK7sndk21pKJMRXFdrLwu0UHbx2lH
/MFYuRBLSHlaRUrtaoghE6Q5R0zwySvm4p5pwujgZakg/KTj+IsLoZI92ZQD+9kwuWqGcgnkEioL
dHCKntW4SJi3q3oZYHEd17gzimJDF7Srk6NWKbBPHe9MUs5aEkpVUs8j9zl4z7YpO41pj4+gkswv
VItr3EkQWwWYwUiQPHCCe1g29wFz6Rm4JR+VWQ4e5cJZ7PEk0MffZkGIRHnSErOpbxblffW6n/PA
Fo2lkaEzrbkRdhwyqakhhg4X/v+38tPGSbd8kiNZ2bkk9Qqf8icwvFY73fbX0SyDT04LrJ0Pf6i8
mHOBYU4/sPuC3OcL8Te87IdbHh2Q5r8fhBmwB6utNAsPzb+wb0Pz8enYgh60nr7ZtdJMTyITUK1d
b3rBBpTomRdBtDRCrke32xavOp91gcMdtBJy1gWM3ZFdsNNAXjivyXQt8/I1UQVys3mcxORGeQ/g
zDjUy776uZ2nsbGq9e3N+tcG+zA8qG6/AI9l3qRBfdrBiiZI76K2FuLG5CGaIFa7vTwHGjZPsYAF
2kEfS0VUZHu7VhF74Iwxl+XItptAxKnyM8kN7elv8DIE13xYg1niLklX84VIQA+kWgtZUEuoiKZ3
4NH0W7eXcF7xDEcH4z9XEYtwVyqIx81YG+St+Iy54UHQKfcFt2u3lR+jWDJDa7wBkaFFJIGvl00N
UKxDHZZdIYlghibO0p2ZmNxy61JyKELCBe3l7LctVBzxk8NlFU0YJXvryU2hIUgFneAXxP4sLFQj
gawuh8OYMIznUsyLundGDsWGKyedF8haGepgdEmDBTVVqN5v4piThWLDA1/YuKtAxxi1Y++NsW7V
NAt8xLcwp7YOIkN3hER+klRE26zJ0g4h7H665Fsm0T4EPUZHblUa0aXCxH1zphAJ0yPb01IshUdj
08pLRsPLDneYqbDzCiGCxSWZdnNkX6Tb+sEnwdaNIShrFO7fnIAiUdR8mrDf5/1buTP3ahvUz25y
9EhH5hV7hPJn+zvnZu8AFWlyTgFz3tHznkBNy17efjU5vwAyNMpycvmecQeaB7VTPBJNPemUxBLB
G/nik2bHxZjl5G4GS/kf0WDq8ZK/Yrh2EUZmHCRKL1W4/I9KKOvdiZViutu91tZ2hqq723TVTfyS
dD/w3NNxP3YTgadrLFi2OeP7sqxF4u2Ky+3ICJTklkBLWdCniuj6qe4MdzFXgSEI7jk7xqWU7S/3
QGv1gseZ9Yy5l8MP5FIsgzPXCD6aJ9dsqWdPHrb3mhAsw7kIJAMOQ6e7JHZzrjHaaZOwlbzMYie/
NSao9HW7I25iD8IEFhF2mBjwOlE+PJeZE6UsmbW9dy0QEi/9R/o0ZRx2x7hmtSHFyAqz3/y29kSK
2YZANp1Kre0fOtAZpIr6fP6saeU0W65uhXbXlGtFjhmQzJuvL/8ruITibPeOrqm4skCqfdXkG7T+
7KC4AXWLvfHxM4oEusKjIoo0F2sGojdiaO7/oyVIq+cGVMaSGu7ROh3YImcXw3BnQYtbUm1l5nvl
E/SHYL2I5Op2nO9rxP2J7KJH38/6fZpzcANfssq2S1IGCBfR5wLD/BLcR40MOJDliM0N9BTBCYLq
Y4gPQIifk/sCywvbsmKDQTtbr9tiMvkZyj2FwUd526+ZKUbY/USlOWqZW5dnFdX/N0nl6pfaK0LZ
DMQfIo+Lx4o4kWTTLUYj+LIfx90LYpRXqz8eJ0Nj4GsfXuppLZFbK61L8T29pOgULF2LDPooNu20
8BRyBnRreXHrzkq/YCbrMksOSaRL6n4PhwI+ab4n14dh0EueVdpGW+6MWwb2sfHvXu8dC77uoUAe
e4lt/Uc9HLIj271onAhYLXbq2hgsBaY+2d6fKhne07Wrpf4pgaADQl1xFMCVoJ63gxE3btvoUuFP
+t8JUSFpEXsiH5tvPjwY5kcpJ/VSARQiuAiKvL+FEZqTbefRGbGr9cJ3g6K9fr/2KZlHR3DihF6U
ClN2JEgdZ9cjDB6TjpaVyU34csF3s5ooSz1S4XsHxLQsdsstI32znoWwPEph9T/pk2TQ3kE02weF
zmUdtGEZ7CqDoja1bbBGOZDZEL8ZJFlf/bHJwjWfauIiooNnHlJ1Is6FuhUUGc2R2DoTaQqnvaEr
ik4uiUrG+zkWIbaLL0fMnYrdl259KCs08WASHRSz9TeiGWrvmLyrJqXcontGk7z1DDR8fiwfqYo8
u9YXHJogiGewV9K6GabUcqQvXwZxHRXMRjJGqB5zY1yO2nLjljfkNoFJjuV+naTX0D2t5uk2VEqT
uoCRO1NiqRqxMYvJuYQkujViqTU0nvr4VqVp7gOuxl9/Myvn9bJou4mrbPKkauwyw75ph94dVKgK
Iw+FHi2fJuCZOXDtMHXAsTJnNTv+/FrebXlsxmjPoBK4aiv5PUmrUNPNAb/Kg4qmIxlkQbVmocJz
+OtNdujjWl3e0ZuRg6bxmKUvhYcVxXZBWzXNmP3ZN4lWxG5OkQ6dzh/n/uqX/mvMJOMr5HRgR5Qk
NBKewmXr1zIaYfA+hjSvEZOXnC1rnZFYOO4gXxrP5+P7xIW0uQQRM8Vf8yGT/D09C1oZa32RGTY+
JlgZgEoKkp8RBFmX4fKxk03mAmiVsxuoaDHHAztAW/QwL1/KGjgP/JwlIt1fRqoyoGgLNFXS3CgG
I4OMZKhBctf16zepM8ZQ/hDVRvBfwLBeMaLXMiZ2O5XBWMZfNtap4q8LtyrKI6qqvZrT8s91LRlt
Zh5822QD7uogf2+RDBs53KkUrT9XAKlHP4KJf6d5fEKAusNTG9oLIl9uXp/234nokUrdZTOaoPk4
1kcdGqKhAwDPrnPxOuAOIBZqQBxzTqDTR/0JgDxH0TnYQkWp3ImpO7NhOVXiT77I2Yzs2/vh52sm
AfSqIult6mrx1893OqnvMYBLW+yWGDNaiM6g6NZLKFDxufVOVFj1YLGXhf/+FEeFIm+hNj7Amljo
0UVStG0k46KcQHOv5ruuaNidEoCzP9neuZrTyRvY+sjfRf4EgIiYMZQnwg2SB6q8EO1q3G4yIz3m
wmWw4Wv4ePSqNq+3SSFtBJqnD1KIFonLEQmvEiYXIgtTT6UOQ209TfpUhe7GyOYLvKpmMufjr7h7
NgTDPsUG7Dkr8IJx1TZjpL6MifL+S5dKAyXTUtrVRoqR+/BFB3HmbP/tG4Au6F7J2A0U/SBASiYK
3HrcLk7QuQgpmAyi1eF9b5Z5qTd21tq+GZl066IBUykbTRbkcHV3wYYLISBKLnnF+ZiL4J3cDOGc
C1kGyDoSXK/yREUVwCcUwcvp0x5ZMkzRt/qLD7QgceYDUhYZhfh41aLUalHt+Y1ZIi69Z6qn1LzM
yoiEyGo333HlXcr5SXpN1ackTjEcBirmW5RTcYtI9n9+mSav1LTmlxfVlAw15VYAek41B05OitdL
Y69HzLOKyOZIPw8Nx2HY8oE3GjenvgNcIyU8k+0uNeEii3VeGIWZQ4Y2kaG76GoX9B5Mwx6oWc9K
VKsX5o9ualwJJZkzMWq+eBpDV7nM/JF8725lQ/2IJNJh34gJPoddpOEbKmWDJNTxMlaRSAnureAO
wOm66X48fT8X86yf61vrvE4JFjcMuoG1jgAZl6+AREkaShnC/2mSg2NoNCiw1qDrAiA8Q99LHGQx
jEyz7Ji11wx6DigH/jKa7VyhgGQcnH9AYdpU1IEpDoJp1zN4Q2V8/Be1a2TYLd68+3o9iVx1HQvu
Ah7w+beQKcwq4gCm7pjHnO+DPem7n811zsDvZcRXb8Hrh88+JWMSP12wpIA+BBYuaW98hW4S8+Ge
9HBnBlzzENchsX6sOmJz7foAhDuc6qJHz1OoDzA1eHNIZhCoV19o+7b+aNP6KHiK7/+Lu5GsLK85
2IFXVcTT1zo8j70xqZq/UD9tVnsz821gI2m4F6GMp7aQPkw6x8ay/61wsrngTyWFYCAEWydvb9Hn
2ro47dcyQmxKerI3x5BT1frmC2IqDdtW0l8x8TxqztrswXiTbVaApgCoiZzKsD89V/pZuuynRb4i
X0pr35J0eS/g7IcREdyN6McVCaew31EXWUKWOdHGAFTcWpI6Tf4/mmMGttAfDk/EccGO6i/Y2014
m7LywkC2Jau9P2oSCj3bxIoJFnP6+GQhN4eYrji0i1V7lycNvmCKiQfTm8dkKU9Xt5ccBz/Ngp8w
nGBMPSRbZq5pQMVPwlOlHvSmnXJpR8SJaHnXg3VSuEgQvZ4xHluSQ/9uG+L/TUwrYn1YJxH/zPf1
A6EOvP2GGLm+21ZqvomIk17Rw0Tq0+XbYCNpN/JN93Fm9XKdfkMSdL7CJpDtZMJFkDpbfhSIPo4v
J/h+go6RPc2KfywC16+fMJnqV6o7ZsxxMXkEp7OGjTeltM9tIbD6PMxnkILwl5WAEw9SoTmanv9W
cgXxIdUHx+hKfHEfY9NnkIn19ps/jD6QETZJ2CbgKxkAKgyzicAWslJXRUH7/p/L6rMWUDF3k+Uc
k79GQQnChExUuhbvTHjoxjpKHZqSlDDtgKsmYOFVb1qwR786z22Dx5JoG0WWwt1cPETS7AjJr6pe
seLFebUxj6TV4Fh5YO4B9kG1nDk/URnVK35HGgNzUDW/yGSZVDOgrG5io3HlroV7xySRDYkfamyK
HWHnFMhy6yKKxYF4J8MP0HPmIy1dHHJPZkpezEcA7uBQ5jvWKlVxB2Lxs3Qxj6CWg5C9PtuBESIl
9tJuISaxdJAmbD+9StvKkioRPdSBqDlsqKJgLSxcySUjQYknO8llVelBF5GnNUXR26cV1H5bJhDZ
h45MnwUwHResPSfVdsYy5V39qmMY5pU21mMFz+/4VoaMyaCihdlONlKP1OFmylLbxnDeMNlIG5KC
8WH3iu5SKVJBM/Xiph9S/t9Iw9QGXUSWxWb5wdb8f1ihRaB2Unu5JqLaAWr1rogjKc0A2sVjhNYL
VXosv0xQb8tpRMSKjNvf7S+0y8cj+cZEXCX8DPFYKkilXtiiZzY/GN40m7n2Zz4p4QspTDm/p7mG
WXJXNDg6SRF6hhlsZFC1vMRmC2UdnUbfLC359D3mezn8Yo4cKumd+ag7P6fkataft6/nZm6/ySWo
1RxYHZuiGTt+GcFSeamz78XsaPPLXuvt2JR8R0M+OIjOe4Y8pkKbHj7lTLcx3NJi5insEUUsk6K8
rMs3dKCaN/1WixZ6IJeC7qzpc/5NSIRpygK99MdnxYtEBB2L+2/6rxHdBK8X/PObECxEsnJLo/8i
Jjn8GIquRkAsW7hcT5DSS+R+U9KRQLjh89ClO84F+OxUILnPkOdY4iwmrYKlQmtut6sRnsbQF6Qm
yQbUIYghtL8aBT0vAXJlWYIrnrqp+dyzW0mFnwTArd+bhr23EwjBGtbPKkvBBkwXUJxrAMGefjTm
gxClzG+QyAQvouyZuIlO4qYoJ55+JQyZs/jCqejhA5XSdlGnVoKD1HvS7/iTt3Fa1Fc3FdwQ3+TL
K0apeciHJvI9oaJHhVvYUdzQVGKn2doCxsS+d77Yk/TKLCHCly62p3WG35WqwufNasT6GenlGmlw
PE8krdIDO5DJXfdh6vjMjxaKgzb6sUQDuoq1jEobu13uuWVHZzOQQ/mDq/B0LdEL0NwYu0IASm+2
JdqoKan1gdk54t0K0es0VtZ/nEMMmflK5Z8ISYA5/OhH+nCD/7v2pxGwvmEEQ6IfwCHpxfy4Shz0
M7ehtaTRZv9D0ShsBZ43qkvw3OQA+ifEv7noH10OWQxnjQHmXt9pHJoN3DC9jL+GEKAZnLBci382
T9l9jdj9BdT3JXvtJ8lBfPY0fBOSXZ8GWlwJAmCtz7bP+8tjG3wXxXAAyoZdC+6wwYGmZBHeVjCs
5tnVbwXUwljdgZ6sZOecH7P+Ajs6SOj+5Y9lBr2rx9QRf+TN5ze+pgyYtnEhNMim9WVaZVdSc1y7
n0JGQleITGnBgi1I911ipRv6xFByAdvnz+OoSQPR+w3065f0EUBNqLKG4EPVQASMEC4Cy0BAzmx3
Iwy8VJN/hqT1dkMETDb+/h1PjWfuh4iVaVqS0pTUq01nOsn4gJR3k2RQpihfZJNfgt2b8QplQ7mk
+8MwGgbxL+2a+3kLHQq89ySJa7wz5LeXlvzCTb8UqVTTBtyJGaqaNIcf8Xq0+ifo1l/U0hlEZ5rC
JqKY58laC4vqjFDZ1UPRO17VYgq3uH9NomYVuRZsaHMDaVE9xKQVs7075sKvdnAYj/2L2ut8pICe
5572pwmn1la8eZc0RYhrEosU8Ytmq1OMLPpH74QM6W5TYPWpDxr+rOQs1ttiXNUn2rP3DWzXIhFA
O+9S9HnJ0PV+vR0IpUgENpLC/3UZ91vQBMnmc0G8//6Dj5ba6Q7jvWT71W1/aKLqHozu152cp8bl
aTeW1Ohu2eUpf8RM/lu3QkD+T1MKPMiLrHW3cwEZTBAYiIrwUAM+XLgG9AtajWF+Sz0tDPwrucpW
GRkZqJegYABh3NJHEEqvWwYeL98cKeRG3iK29GNsyIi+zd92mdhg3TYT8NuA6W4zrj3PIXWu88q/
ZUp5pakW4Ezi3rRYVC1QuOmf76S8C/QT6e1jCgfc5uMSHC6BZQ72bbC5Yyh0cNAXbiiKVUKatJtK
bexgcm6dV5rPRyesbvTq67rSIhGwfErThpeJYi9sXfJpj5qH3sBAFX/j1bvD0afyDrv+G9pkL5GJ
ZdEVOIsaGGFGiWuwufRpdjrNgCtYoOHEXWokwRL0XsjeBvQzWYXsRvD8pg/iiN8sXWn6HoSbP5TP
lgfPTmwVbliEYFgtZ2NZ0X7k8XTs9OQAaTTnM7V75yn4UXs9Wjyt+Mj2tO4EdfOLkplOf2zepQq4
JJayNR/yuUxG5ohkknDBfPi82iM3s4pExVOaCq99iBX1PzfnFLuqasK8FD5gQMUyjvYntqL9viww
DbsQTDcWpnyQCgk/LBjEpBiUF4Uj0IabjJ4RT15KhbgYdES7CeKUUx8Uko7aR2wCJJKINZVblUta
/ySiPmJzLQ9C9z8Yyv6k15Z9T1ShfF58UU6APL9Dj9pHEaIiJUZa1NXJkj707WFc6Sw3FeH3EfEn
g9T1ZSmC6dtq0vBUEBJpr5Lm0ip3b3pTUzEQNKMcIl7VLOlrAV/Ya9OrIT2I1PBUECFsjFOkp610
kgjmZyNahu+ipecTY4XoJCpcmc/uk6BeBWas7LUVuW702wgUG2o8Vw2d5bjIqd6lR4aMmCQJBdom
+X1ntYH2SKdFHsrp6M1KMOxRg3/HwnVLMQ00uLt8YRaRiIq76skD/toP969cuWDroQwWxFx9HtBr
KaBVmPwsnhEZyzkeX/xFnIjU+tcONzSy4D1uOQWSAHiIZV0Tr5ltRmJxPHpZOfaMXX65YNxpxDdY
//WLMS7rhR7Y+CESjQLPFSwvNzIdz8sMpZnQraCmME6qA9jpeHYNpOVmt5b7T4992m19u9BnXNoK
qJwDw9DxR0eryyo8v5gm+WfpQ1X/eEvJFAM/U0X3MtI9bFym1fulktwFkpI41KBnEE2gm6qPpKrO
FT00rnFYmp799BfxDms+iBA7xxzFd9gk1nJg6UXOblQjk2Un5hl9KokuaKSYy5O3Z9iPwvbbopid
IYdLUJdeX2QF2zCfrBwZOekFi6XMrNf/tIuyZjG5sYieqYs7Y9iAOXJ9+PXc8MSfkCEGwxlfZTVG
z+8KmvKYWM73nXunEKqtGgQWyw3AxyyHjl9FdfE/TeCo8/ScTlEMfZeseoGPQDMDYeZlSYb20aMc
13YTscpXjKqhbAttiR4tWes5+xfZBItwfzP4KGsSZ8PeenTx6AweLJaskQzXbTsh6hn2EyiE0SWx
/CinwTTRCHLTI3x9otwKLvSY2ghcrrbHY9cZnJF2DgPMMFFA/8OKmwFTp+8sMO8nTzHj3g0sIVyY
fg8NLhwmejdeR+v9lTMXenmavSMetZQrSBg0za06GbNvK14kYxBh6QAUfULyg2WovzEmkpMpd4LE
2FHHpQBQtpZiC7J7aKmzQh151Kq5dfGModsUUalH3S0BIqTyMEf6xbmLEgRUmJctFOXB95kDMBKW
Km6Q07BT1e9GU0BqulxcwkVcQrYc9o3kIAOHsr89o4twAJzqvd5hqiHcuvc6qpne85qLPz9F3b2C
XqNMge64XqpX5DEY2pNrsrWUqStFlVwIfXyqgjmBRjt6C/6SWYKEaZaXOkRnOvaOhC+rZAsnaeHK
154p30wkoIk89/CjY2JDfvfE/TWgOPS2uQbQepvd3gPQ+xfCyriIcJ2ZjANT+r+SiWq4GxFLh9nb
/kJERwD8B1LaySZDatm3rKpVQd5atAglZTcytWTepUzTZ5ZcrafVf/EZGx8XBjD5AfQ65cSRN4As
dXXqoa3oOpgFFFB5hrjOYy6L008Sg5mYQt+oZFigSEJlSUZkyhfIEurhNXICiNRXYlOOk4fSgA6c
0VnGvaZMwT8WPphWCWbId0Zrrru72XPHTwqT0+pTwLnLIAzYpweMeKS6X+oXmsO1dELFTboWEivI
P16SMNIXjBFuznX4eS3KBVTfniteUlCdWvjVQQaP3Q6a1LDjjgTcESZu38NXO/Fm0DKmMdSuIYIQ
7qcISouVrw/nwMespiHlD1Dmj4aVDFflFTrXFSe8C6J+8lYduILY7BThwLpIIb/IUYVP0JceRHqh
r+vMRLCdRR9i3efRLBxmmrLCSdKutrT3kwKgkXO9fnII/3OVfwloVLYvQJ+McyOSYJicCfyFdeHH
Qwm/ISCu8WJLJYm2i3A6s+h3fr5vshNT5IpdtAKnbOBDQXe+nQXTAf1klcxoHdrxY3Mdw2w8R/jR
GyB04ZAdpjQ6XlEk0V/lghWdSWOAW0HCXDTBK5jKmdqGwQRVEJqLABpOAMcyXncz/HtVxilarzn0
2Rphxr077AEGaK3k8sQ0X7z39DOFCVePuOhSmt5i62/nMZL0kXewrLG3mqlP0y+wmboWeGlsCA1+
UbAnB6ABi3syTlBmDNZwS9OJ0QtOlex+yeh9lvRbo91+9mJ6gY89jAOdHo38iN9b57AcjfaWJShj
Ce+6LXbSn1COcTXkN/xgBGvh0TqTyzZCBaIlognKUumLtwgmcAayM3Ijw6eQIsAM4NCp9qi/dRk2
UU0kkzqoEpNTIKy7tvrxzxUxLTkLqhYpQoS0PFJzGa0dGViYLBT9RV4KIhBaeJXi25b/l8suWsq8
kV2mRvcdUrdjnYlRqhv18q4MfuqtDAXgt8AEXdhBE2UY4ES2yV+vDM7kNfJAohN9WZ45bvL/WRQ4
kpWcmTBj3DrpxD1HPv2NB9W2ehml93zMTMKlYVu7yhNSu1gw59pFw7uh+UE6QPlMsva+wCbyGb4v
4QXtQEV8NMRKB3bq6ZHRQsY4QEhenbIHOIZ8V9PVjOaszQPQ6GuuebWVIDbVoTwyfE6zZu0X+Qxv
/EuTgEcz7/REQM9Eq/tArjUJcs/dcpruHi+RmxpC8YpOey6gHyh7SPT1pHfbnhevsjj+RnkKgzRV
7uZBU/OYX2bIM9JMjGqQ0C7RIWxj7VaZnzbWyLX3VgwMzoaH7rSDQj1J2kUYNnV2eii06EpLzUhT
R/ZRitEWnFfZi2AodD9wvneOPeTMySjz1Xcnnauvd1bYeLt3c+BWPHqDx+1o6ZrcvD9Sz6HSyuHx
4clAWCkkBqWLWpg0kQaNWZ77X/3qkx5CFxEBcDTS+G30D0OIlzvrR49RsGJs+MPxgckvwB8VVDuM
V9OwRI5Pyn9+Tl7OfbXAAV7bsDoaBWtAIWajRFcOlbYxCB5e6JifmrAQZTjyXTbfKMM244eQP2pE
iMvtXfab3IL50/gMeLCobtUVm8nWlcrphmEku/Mdn1yCw5aX8dxCb/ky50dM00BC6R/dM+yZ4MDa
sEK+Qn4+f4cH8FDpBtBoO26+Z0njMfcdmwbuT+Igew0yE/Pqxh9BKz+afjnvGrWMyJ9NJsUwJPZj
XxvtXWjOMGhAzHdWxJpCaoNqVrcsbP/sLM8ydTPCrsDzieZed4djU95OoZfs7KtJFfc6ZMDdtEE7
7CMYupVMSz8k8y4fmB+5KRj0OAvyPdljhqdbivZZi3xuZXvFR63usgkRrgdgjAfdgCm4P7fRqWDy
74BJrMJhqA+F/oamGulj/kxay++OsiOLIoxiSS52eQwuCF8yFugDHl5Q6vUf6DXdVHc6+ompLcSz
daQ350zK6uCPC1Zw/SK2/9mXBNskAfCP7RLMKZZhnGySyLsWJRZS7MvP9R+4xDrhbdtFuUuLeuIG
KPq9NaChWDsl22z23NiRUmvX/O7f1eXV/c7dCFbopIUCLJHIW6pl9w/pGrifzWrm3oL9Z++lPvqB
x0O0OZFU2Di6nWENZ0GWddBxkCOjbPa8hrH0XBE7wc9iLDRKI/twhCfApo4OBZBN+wXpoTUIS++o
A46kXAL0ARtsr++9ofCf6elMGqV3qhtJNuoVi6TEJdF9YAlL1r6veiXTtclAOHkNiqKmXSoy34ps
mD47IW6rMQcMvxpZHqxZ8r61lnOhPLoEo8IZ20EH+Fi1Aypi5K3YXQuhCA7s+xLGePEpBirEDi7K
+z+l7IXdco7xyh8lFi+9RJL/vWgzQEv6FX4Jja6cAEkcz0L3mazjjOAuIL4BRzv5gkT08cqthFxv
gFE8nN+3wvMicuk9dD6fpN28XnQ3vYhhwRJ5fJqQZrvrlCwtiqSI0faliT7GHrJl5FjAeIHi8jQz
+W2RUKzkAPcZ90N++fK/Id+KKK7zWNdVIdK6A9ihhawFwgZUtmmEYK4o+XDQu1qDPobAK6VRhQXy
hmoJJrtryL23/LGkg9jCZNXIxCC7bo/S7lIZy3uLMjB/PMx2Yte6rE0LTgehPqGkA1uULrZ8Kyzl
CaF9yk7rmJKg7iT3Y45pejo23PO3Ze8NDpw4ACKUTpqqeR0MxVbkh6CLBac477Tv0EOoCK0EHtAZ
XubwkbNVlQBQrQkVSqecLmirE1IlAfFm8DSJleMyYBxYPvfQBuLqSQ6KAtiP0iCQXYs/RAFsJ1b2
aRbsQAFBzbZP5Dz9o1MSqLv0FCbPf40L8SFmQUgW85ffJHOCYlPQWj/Q7LD/QRVmPow8NaqARDWF
ARI5pzUTTqvRmKKJhUmsyASRqTH7GNiGdocz+bWNXjdkY3vMxybwmFwaGZv3ozcufCPXZ8rE6HQX
RL1/omuccy5G3nmkz1wkJjIAD+Pcc7n0Mf7PcoGcNXQU4X7KdXkXkAv3xaZVIs6hW854dhBxR2es
pqqWaw5RLRANW18nn5j5VuYo8hDNn2pHj96XlsuB/iAwEr5kSLszPR+ZD6agGiJTE0N1a0Cj06l0
1/QcEJweRi5wT7iUcn17+MSNRSOaWpW0ECxoHGolbeeZgk2NRhAzfJVoirM+hhw8CgrzN5H0ke4R
phmy1n8V1boDnY1aHi7go0UZ3MowAaTll2cM1WGXI6Uf6Nzpp9D5um4eoVnmWS+wUPlDLztc3bYy
aiOo9HdbEGQDguvApTCyV//wMDNcIIvQXPfXuJLpkV3HtYMBWiFXcz0drmPxb1Mf/TAiRlojPbJf
PVssJFuebuhko+sIJWYQD2ISAXFlxVykDvWl4zE/iqf6p+NhbUqjTWSL930HBOUdl1OnoiWfWKBb
NsJHmCcfKg3PjYWzzESKHNKGlj2hL7+GX4XQ3a0Y5YI/wanC7Q5RI726NCJbGqBUOfZ3G+ZGCaob
Z04K7HcOs4gXDUfmwQn51++oHF6uT9XWMLkhSirfQUFJfGKFFHtQu/iubuN6krcBD7JI8DLI/+ki
YJWsipqyGgZCw00jEjXUD/vAbJI2dH4iDt7Ex5tmAQmpa3PYmxfRPSWZnAIQMPPfxJ9rrkE9FcV3
SYf/iz0mN+DRSrsOmc8sUKP1KP9nrsbM/vhZXbzSbg6ToP4TrK59HXfMss+/KlE6wdMWeS676L4H
FzWQVqnnQY0xS+KAV4N+sb2ppXy8YtzQngpEI9im/6QAiWAlrNpFIh2+sCy60g0W9EZuKZa92j77
bSgR16Dz+WGZsI8ZrrITPi6Ekf3oEnrapPiOsvRg8xObbTvobmtuDIaJncY/U131n4sRMStQCHhJ
LEEvuzchj+FxuwAoSc9QuQwSmOYQmKoWpELiBDUyTwmrqjsQrntEmE3jtdGJ+Pt75M02fk7oTrs0
ZZFcbfMgphbJwUd8x7qdehNYH2auDL9vdMZ85qxsknKRbpnuqpT86oDazw+5zHB0oEqkUPYuDaXv
kB+mHC5PC3DhJ90RkPec3MxC7/stL4XizRBazt/FD81fq+oltmF2f3UTY/W9Kh8HDYgaSiuU1GBj
gXIMs6xbzdmYx5M0GZ2iCzyuwoN71AyovlpCH34MeCNEYOwu83GVombmtnYpcviAZe4GLPCzRqLh
XUASE25ByUQEHFYha/FLUpc5vsmbVyi2r5QLSwZN1sJN8g2flcUdbpPYjqM55e4yW1pod3kwi1Gf
MfwwpKRgiPS8hWIxs4Tu1FdM/gxCMI8cTlonTAqMANHbt5ZG59UDpceUxAmE1zo1bpUe7CA0vIp9
W0myI4blG3CDfRYpyehWxyt1Tjaeg45b5hyrhMri5JO4EasKJI69NP6e4SWZmHdmct7qrVEKnoVr
h+87xU2pCfqWDFmw2Juqm+hXaLgrkp5nJ3lnD2pVdk3FYa7PMwJgzxTgCYnYhAAKpIhGUnP+Fi3h
M4SNNEannE3/AfvPLMgeJBjsIRdgg9cf+gxLl75zs4OtfaE/YWANUWdAoc+XJ++MLCPzsWYQQHPH
hlhj+XIkS3vu4RyyhVR90A3FEZzPeg6cI8HCkWzOChfPbbfVnjsOXcTa/Of+R6rSdomMV07fHTBV
T8YBI9dlWXSsoQelC6CBOdSWi4CJbKxttckRpzV1t5x71wUaoqSozjQKaNqgxA0gW6MsUgG7bljA
cK3+sJ5GI6CCvR2uIoWEsvn4UxI4QePhgWRwKeEXosFfOvTue0ysz8LtfhAuXyFskhrY+PoQ10HZ
WeEHLd6IVG5emFKRx2kJ9nn1scX1M50iHlqnTDjJsNGA6kjjW54/HriwKwiXHTftCixwBJrSrik1
GMdajn258FtVqO+nj7HdIyv0O5FCPeRplXIrmRcXnMEIHi5TG2AHyZh/t6FMZlxyqW5Cw5ZtbyZY
OjAHnP2wUWLVD4aMxQkY5rFezjk5aKFhxIDIfdwWCgojVN/Rbfg2x/uq7rtuxuTg1WwX8y8hdzip
b+80+ThuNsiN9d2R/eMAJCP1TA4gCVstZtYlSepiIc1/Re8BXCpHOYhxD6Bz2Na59hNWpJA9ZFy4
mlTkELvlT0oClC5HYhBDjoPMusS1g5Wrfqw7nw0zAsyheRC+CnFnOkIvq4cA6Mhh3gP93pdUHIHR
M0bePtJVidUdmbsdYVyFC4/bRv/dldCZ1AoKGHGgx4jkpIGRXdLoCmpBs47yujnhtzGmSXfQR2Yi
TPzWFzEyA2cIiJIFwG+/FqmZ918iFo219FVTEyEJ/WgpHu0EOKnRfk8UdlNQL491VwvCilSnsI8k
ZuRFETHO1up1/QRlVMzuZYJqtXn80vjvb8ngLVqKJEVFwD74x8/20+L8hmjLQ1GUHkcbI9Rm473l
e4lTW6h6Yhc8uAwTJ+PqGp3N5Gak1z20jbHChZmP+IzOW2TVyFGqj/2chPwM6Jmx/ckYCitAMK4I
Ld4ayfFJt5CT3jvsaQ1atyjHsaPqSxJL8x5qlzcuw/7OisgF+pq1CekT5cvjW4ZtWOX2Y6c82VOx
By9zq9+VpV+2RemiZ0bGCKXYgCugy3Mz8OC5fb7vE+A4B2yAXczapfZabx2qfe1gp4NPYQyxlRhL
w03/E3S+04wHzg90kK8ILFT82PaspPtlodq7RXv46n6tlNXiW9dvvT5FhbSIVosg8UqlNm5Cs7sV
Wxy3yv//fjseqR2+jUP6AzWznUcLutkDWjWN4wKCMAbq0rb9Kc/Myj7t0xk0xR7f5CfT+3D2Y+Pi
Htj8cu1q4wAoYPsi1C8ByBA1EEsQC3IU5+RbXSKPE++kQ46Q7/yOyiUWRdlfioc3GukRziRwb1tx
EejYYWXqZAYayTxzMGqe3D+JzmyDUnX2s1u3H13ltnjNTcwlqquXaAWJ3fOv7Bgnbw2qshhPfQeb
Up2OxPu/tDm0rRfj0PoGjc84ISjDk0CoGcoxBEZA0ZtO242vVME5mP2+8aBWTj08ZR/TypHoeRpv
P6cSDaqnF1U9W7rvGp16Tn0hIz6FAQ5B2bKk6PO1ZdgxMDfQnyRHBZFHkAFPnQqMuiYAnm26Prqq
cRFtdNswL3D1ufLKJTTVj5oo2WP6Ikt8z4MspBM8ngDvgTSV2vVmquy27vmbyEEXyndCoTt8dXQF
cESj1+YvKYEBduhuJDxoYB/xxGPmtMNY/QvLCNKd53LBAqJwjDFc1pP2SHzBp+e4wldAT4wsJWEc
d6Yjp90BpK7ViMISN7mSf31+TfB9vLypYgtrrkwqIl/mEDfEXH2Ewxizq14hbrNYUIXX65dLaHYw
XnvDLyB9LtugJKMSZGFybg3Qzo+5Yt/mAj14qlapjos9zh/A+b4ULvsipCzI+IWzzs8hiKct7lz1
TUQIXoPlsQxp27WuPMcYe7HacjogwP2MxwzfBX5n7a+ugb0lP1TgWS+MIE/VdC96cjAfHDAziImC
IUOlHTLfrjmToLObQjOoQb5FvRnT3C6YG9CZG1VRCqaC6fa5vWVqUdJEwxJ3+7B836dVEeGQ01lW
UHZ2eIwHUiJzAOzgz20Qu8Qw5aL516PMyNdq1eMpLnlHcmwiwZ+zR5T/CRufAOVIdxKBcXGaMEEF
AY7tUZyvkw73N0fDvrgYU3FVEK9efOU73mEhdLPo6PRPgmMOJj2XF4M/7kxbYCDyKfjhR9CBTNm+
YTr7V/f8LIX9ZeCuwc7QL6Roch6XtUX5lhQ2ufjhx8lD6ebWcnFOWTZ3j8C/lpBf/7Lr70rTbSJW
ZPyrZZf8868TDDdyS5/kYLkMIMyBVne7ErQQygy3Spsnln5CWeVUNVp/55zu/5k+mQ/ER5XeaYQf
+E3BgxPYmr0s8w5dwVW3hVT3oj3Ji+mM5psmUfjJGKe54i1Fwy8IvZod3cnqhiv+g2+/smUwihEL
qRQmA0HVNDLHB+j8lWvMUBY5NJbcUb059kg+VTNUTg/PYAXTmF5pLqUrXxGICqsiRNV5jUlxspcB
WL/5dfKqH4DSOxnwd5WTgUYCLf3d22XppmlMBgYALhk8wpylEPsK/vu5uWrUhklQIoyBcAg/Ys93
0bUNgN7Cao2DcLCzYAq6+cWVN3hXgX8T57pcG2OElzrIi62URFsPHzLXgnLwyjz5grmQrTy0+oxa
Sb48JhJliPvt9eZtm/tUJIQLpbTghlg38jyxfKhGLwzf/ZeCyS/IV65zpobDHnCzJw08/tR5kMAl
tSewXjrVPmkAMPOX8BoF/4Am99ObFID+ei3NNTeYQdMSdm5ncoMbwtpeS8K03C5yxVjb2/UkOWpm
HVU6JsBXWkqqK+t41hqBrVQxy4EMfkgQGpvWNdR+nMxqNwlsxe07ET/lhMBywMhhLSaDHRORIuRe
cuQPiosB68Rgx0ql/96vh7VbvtstjEHsM3/AQCTgVtf7fZFd5s3YRrlnvdjlvXJWBLGYomFojPyl
54XZ9ObmL50P3ROWj5B3xlNLuTAX4sM6pqDBewqrCAmFZ6+thBfcNvy81s5lJ3QNyVFcnOngmayZ
lL0ZQ/dCPK2T7/P/H23SAMXZvRUWWxYikKFfz1zNMWm5GjLn2254IGLb6RK+ELfa8+tDV9P81Qrf
zKrbwYUalz3HJHe3rXMYQzjgiXtnqWTBhZZ9UMSqC0XS2fdBuwVjHxxkDkF4/0peBg3Cvu4elZj0
3wTU1Tsn21VulVs/1SFrq1Hpv1zaB1WiENCdumYnDIiZ1BMyVXD6dzldb6OSquhlOc0OCZc08GCr
T0x8xsK3d/HJtI8PpgY/HbnCjgpEf7nDf5E9rMk4GGRdYRR3ruzJS/6qcMz0cyVZa0AUj1Bvx7F6
Gk1fUTDqRi4Ng+1rWswz2xXNIEdg8G5ZuNBJj0tFXBQADYELnukzWAbuPnEij0/xmYWJ2Z3aMakJ
NC3+KagxZ1SZECICeTIIBZvBpLTbfIdIt5rfsEuVOk5MKNoEY5JEsIjGjD6clI1XQJxIfrr51K3J
Cuf76nJhq/BMb2cUemrMz1xgj93/fchqghGggsWdBpXbJDXyG6JWC1zgaeQfMNpuOBkupWl6UZIN
3AlaAewEegVD1wgu6lXgLzwEK2wXMGSK1scwv4rayfX6DSp8KF3HoV4h6mbCwzu8gcBIRFNMe2jg
JXx8h7WzzOQSdpH8fDYkxsJavA4V8rF4NDRsm5tPID+QW/0cwyE2cyIdtTQJfofk1KtjC5JYPdgh
gU/+vJhoz7GIPUQC1YtmWDSkttv3xSTs9HQYJWNkVD+Sv91w7asDa9LgI1Rd4ADjwxlJ11gkCDcM
iWKovi8tg/Yt6/QmIRLaJrOiWbOSVNrrvGT3CqPym8Uc9mZqWjdvyX5nY+PwjobVo63dVskrfZru
Xzcc7BaLp8wFxgeDG6xj4YS2fl4d7KtVFlsT83G2YOfznAtuZOxEFfxSKqCBOOgkpcvKeVxgWO6I
9fPSj4eBcMU9eeNaxmR13DFoJ+Ku8Bu5+Iv2EMaJc1snJUL52mQf6lWYyRfps0jtleJgXu3sVMRv
9pVJxGChRwzO/XSnvRt7aH/Vdt+Yp/N6p5lkR60sPkiOn2RaorQjpodxmRFGX/sZaltnBxhnO7IK
rIaFK90TkHigy0ah9SnOG1n5MQobxDkBiI5GfGV5skvnl/THc6eCedfroaO5B1HCpkGr5UA1Cexf
vlUqd/r7+dAfYn2pLYDKJICsR4d+5qQFPTMPcBfNo6rr1BAl2SbKxx4dAo+Feo8RTGk7FR+KGpqO
LEyQ2dkWiGEnXRLJiHULPFPhJJwu7CfaregfFXuX/764EXlxxySOcdIaLv8MBC20g+na62OenfBR
hvc7/aG2WJrErvH+w88U6QVNEdOM/L3Hy0cx4wbk2R7ZBpoWSx+VMoQRZipB3Jm/ajOztQn25xpq
MoINUAL9YXCMZuYfJemPslAKxQzDZEDU666WevBz8QpWcj3mpGzA+sZ1If5AlXxgPRc4/SA7TDQB
Ik/eafltfaUOuoKisV0brBEm7EtUJgGOUR2fHsEX2GfNV7e15Zrdeue9g8UP9O7UNcC+NlmlCHxx
dmJlw8JHSPEhNVPWsLfzX3YpWXETfNNJkzeJoGy1C9VBcF8uH0F7jAlOGXJsgNnjC3EX3KwRZBIR
BR9APDpaB/yIy1SdD4tvnkS0m3/vc2H8h/djNy/tMhqtjP8wb7AFXsllh4BE8MzusN+JBIAIQuOg
6mcy7h4B4RbgXwvscb3va5MBpwRs4994m4iFpl5s9MUW4MrYU6MeLJOjuAECg8c35jbj10Pf2xJv
RS4k0Opvlh2HHbuhjEjrgc0YlU0FPpQAELxWfh4LIUmjfOwKlMNRYVle+o8Ry2G1PwahG2yAyptY
N3EDD8SBeAO8oYjoXrNZFmkz2p2L/W6i6QrWJi7zuNe63m1H6dPozxcZv5b30wQfMMZUH+w/6u/6
wU/q94R3qUAGxd7MJGGXL+igcE6tUJQHqlLRBZhAq4aBK3wFstdf2IziRky0C8WEzQ6DfWjFaGsQ
DwUfebGMj5g0He49woHtShRUIJwAVTO8xRKVrbbKoR9vzdVxOCWm1wFJ5B12qLMD8OC8uIcpOttS
ikycJ/29KnT0T4CIB5+K5SXxboT9/7yoop6I2nFabYV4GWUU7rVZWAkOg2PBR8E2QH6cjr6o3M5O
mCzjkFhYnOA+34AwpqVhsy0eKGXRYa4jw72g4tCNNQuSSnMR3B46TFSIDTg7La+AdPLWZM0sisl9
/cXGfVbPyshnt5tBhJBMymOUZznx59XtMug3m3O23q05LX4Ory8tRj2DdMipWv1dHngpiLwSXLgj
jicwMYq3mcHaskIRSGfc/o9cCbxMe1OVkAFCPTmUbteBAcYbwh+c46cmNKrnIlihqNJhNkm5zNMR
Dd1v5m++rmV/1dndcyeJLPZtv4J95m5h+d1DRbR1GNxauculNts6DYyOuPqqkhNfjA5/VK1i2LLG
msOgPRCFFE1rTNnj8dXSbIC+6+OOjg4LjJ1Rj10Qnutu1t8LfdNSV2MP8uJO6CUUx/WZWxYm2ZaD
me3EzsY494IfK5dhq6vk8hNSlWueFBth6A30agCgKbD/KnpynpNqTS9MzNL/KulXhDjpeDLca0fA
3NCwcOrVlET8Pz/uxrUn6UrwskNZD9Dtk2Bn7hXnDh2rVRvJ1MFryT+K7a68y8XcaWOOI8I+HWBb
xV5IIWh/eFE8lYHus2xY/CaDZVqephmjU1l8Sl3uHJLy7n36BG3Sp3MNSR41UgC/pgXMFR1/KSZe
72tCxpYNP6b2OHKKp3lseMH7VFfzrmZnbjji4loUP90WsfiZl9h/UljN1Eu2a4aY4+/DYYlcN4OK
XiR+o9NfRnet4iIDHdklrKPe7etaq9tyEld/Gcb1v2GrYCYmdCweyclFrlhZvPSiCPLvV42EFm8z
SGM9lCg1QeoQzSVXpJb1PxlNV645VlJhfMFGZVby0OKYOVLXl9OKqVkB2VlveqOS0/2FxafwMVaL
rdc8Sm/nQinIwxjsi7GYC7NOUY/COXDL1P9xKyAerfRI8Buv2qw7by+bTjd35uEYGtI0fC6RjswD
S9pPe4Zm2A9rw690qZ6t+6zwDiyXvU8gjuWwxObxPYI0UhWYe8y/0FrnVTGiXbST36XXT3VX0Pon
PhCAIBafsPRf/SjvtpLGF4HQ/d+a+fQzX/VaggP2Ja77hn6HMRg8X0Xn5KgVP1QGflfq3ILqxme5
cWoBGusGDs1g7SsoxzwbzyBLftkVM1XoSxyn3K9I5evbGJA5IUSWHd/1K9CLePIS+Bjm0GdobUzA
jQ90+MdI45JA2zKrcUtBC9gDHQFVJ9UuE0qZLTR/YQNkmXSiJMGLha+aeaZH8j1s1Fi3yWHAGX0f
8dE0u82Vv2q8+eQatZ9l+72D6OH6lWFTRK5h/3/qW4UxiFeJqSvTUQNb9afRo4csXRpEMU7Q96QJ
HbaxVWvdTMCoHUWmAW2iSYz9gNJz+mLfqTliwnqXfQE5Vaf48dRiw4rBOlJD6OsrB6bSeXyl+UGn
SuNrwMo3OG4FwuRyKlZ8hGKex5NJjoHsBLHm1Xe64g9e2JV0/Y584M8+8zfVu0JSlUMnKKn1ofGf
C2+94iwBtXnFL0KmbBz/BardUS5cqeI0OJrnzpjYjdPnGrKW4ERYLhT6aXRultOHJZyGDCgRkACV
W8yNuHXI3FpW5bpfBYrnZ7kkzXh2WY0PzH5sc/wrGzEL/X3y2LFfA3Xp9Vu/jf09cdqAvRFDMk5Y
oGUwH8P+4JGJoClnrnUyy1FFp7XgFAqT+C3Jn9iu1V2IruDxcoqJrWBqT31Lss6dE4dWyi0y5aWT
Yp9y2B0bfhJG5IRJLClrH1TIXb9ddyIjVE9COtBU4AU/8NKuR+JIDejfnZzByuUkxm8VQ3mHmpNc
WmSzhiDs3d9/vHv+T8shmnvH0D1MZbN/hNagZuc3SJ5UFbkJFsR8FA5Ud7doBUB41UpDhchyJi71
Jf07h+InSxFH5LOrzMN8Kox8UVMU4wbUQ1ZmkFCglT5BmQeNyOkJ3Q6k1LYQukDIc9rTPCLxYyre
yq105evOrcu6sqoaWehLQR2RkhuK41dz8ikqRcZCoajvhEAkRkmXenKVIu/hxX0ozNcWUCKtzB4c
s0vHtfJnDWgQ5EILbm1k45yAqyukQxB8z1uK0n6b41Pz6xJVINrs4lN1J4RLt044AsnTb6ZIAJ0+
dY2BE5v85bzepANh6KVB+hAOzjkquTPfXm39a08zOka4iPFMXXe6/cv7JsDNJ5wybiwEPOIDiwUi
kcFbLNj+rKeleeC4SidRoPKWHir+ZMTLT0hl0Vr9inu5FoxzUh/O8iPBfmqgQlv+7amx77EObz7Z
fJnUBX2zYgV+gGEk06+75vJObtBJlCe5n3yUn7w74OExvdxLlrIHWlayLMh77Fwf5QuTe4b/IrLt
IfvAYmL8BTsxIGVaOH7C4cUZ6GPb7+az/pmkQWau1jPpX3CvyYUuwM4TbRjV+COgtb7khzAkaoRv
2AuSownZBbvZK8g+HbJLfP+NIZUhw09ws6/lcghyVcTCgy0DhbcPe9LCLt9IrB5IG/XMvwglsoVk
UxM3uMRV568JojLRjteOr0oh8QeuLVtAjCt1FiJhFVGTDSa/2npwKnj1hjYghV5uEOxOrCvdU6fo
S2NQ+V8pgkLIUAMp5Ery/czN6xg6C8jsXWI6S4CEsqPuFSRUvlDDPIdA2FZ4m65vGwCLCyDe7mHE
7LXFEFlhpUOq6EopT2B6GpQca7zHJEApspgT0wU4EXtnTcBZYslwOlhkDD7TxgWbTWVEFADvTSnH
6ccm0izXKiLYyOBBU9UILQaQyuZ/PeU7kx+P5/ILueNBUbwW3CGkEvzSFMSXD/GgLJtmS9SFvUwE
23Je6mc1mA5z13ka3RvD645tJDqdduTxDo8hTG7VTq0WTxj4lGaTVv5WhcIARXdcoaHu5mwUcVJj
dJFSrhKpYxDXkGgmcztDw9/MfVwWZjxmFF8V3osdh0yhC6HTNteAtcyrbF2WXateQpO1cKg1xrbR
3kSDrOKA2alCEJg8FdznfJyO7qNw4idtJuluBLIW6kPe1SrZXkfPBDAlvhZvPEhgRm2e9ROwURvR
bhRGf1+4RwdWsqZblU57RKdK5VR1ETCSLEcJMJxPeZ+Xn5qwNAo5lDw59rMZPNFGqOD463/HwWuT
i4kSyLSryPzScLvgHmIMvrCvdXHd+XXDvE7Kvk4emwG4WNfXQO3U2QV0SWnYeJO5Kfo1mhfSEhyH
O/X4PxwDU2oBkeVJgpPmfuzhx74O5LkwotkDjQFnaQ+S6z3JcJFvIUd4rqmu7sXFC5HcBxCOZtYk
RcFcqT7gDu0NFe5Z7zzCq/XES7smWy/dZpbiwbNupft8+D49/xgLym9RIB+mnep/tR1r3LTA4MVn
/xAJF9sORYnwilGInoDJKfMlXoPDS8yShueT8e/bMb26BCaK3VjDwyPU54hEd14okU2GNqn95rXK
mgIzowdSPuBRNfOVeTHac4T8oW7DDGGzAwGfd6S/PLzHA0WCUZibchfvJyv2xAhGNYY1mxAt0EJN
YLb9x/Ifdld9Ziulz8VkxLrV0Q6Keb0JDoR9+/eyZm3Wq39aF0Ul2MB9dsNOvjUY59BE4yL9SJ0f
PSKJJpi7wo3MC6Xb2JQ7b1rOl9cagfyaIy3Joto3mQXAPGpUoXYjHaRE2/hCRXFUCIn4BohYVUkF
/V2QVe7jO0SRTtiHc3XyJvu5x0VpJfPHvT/rVQ87P5zpJvrW4YdY+8Eh3LzlsL6ZoKwn0ltQqLp+
mLzFdMeYSxqDZKXc5HX4+z6GnuqoUe599WJpQpgjFf2QTLWfowPytFpQKW3EKjHtt5T6/UsidRiZ
kLoK9Tl185dCbbK4ysSQ2DYLSQ1yfDGUl9iphV3ASo315fDfw2oWQbpXPMa4m+mt3hGfaeB2iCgz
BVEDt3F+GewRYYfgfc1zUe8LaSGVDZzENuatyDt8VrFk9eKNgkImC3PRJgEra/ERnDCqIyXraHXz
+ZztuyLWyl259XFljRoB7xo0RT8XVmtVxPG+PYemYDuVQqLbiTaTToP1Tdy83BqrdIPgOnja6hj4
xPV6wqXqueZEXEt+slilKS8cLYswFSxGL174SUA+srOVOyxhhf1FtDCp81226UJQHqNWOgaKHBZh
ECyuHLbDHPxWeMTLrDSiKN+hkkORw6IdJ072ASWx30U4dazGrD0YeOClpODdtVuOrVB5UdY2Tw+E
v2MmrkUbPxmLy0a2cRxqAaBHc0ZPCaGxleRO2bfna3Z/8IDgmmkswXwJIvXnPxmAYahAz7b0W6Ic
4mME2KCUasiDJlDOmad4fZBDD6mlDL6UC5jNKmn0+tpE1YdAqRNQCMcPYH2c8l6ziEE4R5ydzt2b
BF6uH81iY3KV843a/p31SoEhM4n0vlTEgufViOYWJFKn8GYPCWuOSvIRDCn5hEjyClqA+ImHQtU8
kAdUXyRx5T612W+Vilz2CRUH2JLYlaBdh+S+W3QRydEgedUWRwgUuoTAgAybw2L3S8Mdw2se1Izs
IZCq/kojqZUDgjsUZBJXn0oVeL+8IiiSqhJvZ4tua1m1kscri99lLtzXXG8U+jevAoZqCIz20Dbt
KfYyq8MP6yUXM+a6PkBVRx/ftkTFfJWpkGtcAkneGn3sFDSRJWMTG8QhL80ipjX35wFCfTAWGz4P
hsDHruVam5rVNZbzSKr8L6slClLh5/o4+fJ0+N0lN1sy4TJxmVtrj72ROyPz0Ax1KV12cWooqsb5
6gm++TIsWmON6ovzOkJT2XrnnpMu/vz3phVyPh4TwJZBWME/3IXyWKKVg5RdzNn9SMQXXYWSc9Ux
iyEvhz6luhuHtzymSCjZ2XwccPSKyTjJQW1dghgZQIy6n/Ecqvwvw/UWt04S47mE2pnbGIh8Jc3j
liunENtQdJ19Cdrma4GO1Ve3+J0Qkp2Ibfj49xrG474sc4FvKlHStqW7zkfIAJHX1TOiL4FDQkHm
9/c5WbgElyNZWoeIbUuEiGskM0O9EVnSUwmQAwTRLw2Xa2h3wz23xqwzQtAWchIeMcu6lK09vMfO
ZHFJT34ULI+LykncuxiKBTKmQzkfyLH4NN6RTuWFEDNAcSwy+2+ZQrpI9JDrG0jJTd5VkCKtJCfe
Z7PH/ZmpWIwgEnUJe8dITfXXQJy2/pmtu9uIqTsDq97kLEQGhpLBDjUKQ8l2GWwfP68HHrD2Wsl0
v1S3gNXYyJXt1WAYnMOKYqz4caKRQ4ynTY3NY9G9INJ59z+H1J5JUYWlwuCRVa0qHOUdFb7v7hHf
inLjwmYkWi+DTYX8dHFgBH7jIMJMWiGW1j47RA+VPayFTdCRlYD3fSCSxSqjV6jJtcZmTfjy8nGm
0+Nj1LwRUOEx/n/Cvp6M3yA4EUXag8Kc4UZUWTDseTDnoKqI/3Igwr5cAohBaH1/cjjotJ9CUW7h
+MmNFY2O49Vvq6NLC32up77Y+m2yc6kuMAoOo4XXPVyFsPMcLXVXBF2rnUDCZQnL3UfjNPrNi8e7
AiEUp08sB0CEBr1odcTX/1rXYktM32ItmRmQRJfDZBDQB1kh0lINW4niSo/3t30ZK44rQ2NXxrtW
w7XdiDMLrwIdKKMsHbUsB9VEYA0C7wKYmNI00sKi4fJvn5dGqlkG/AiF4OqT/o5Ti0EqoYFWMcej
bPVKYIky0TBrTYBYb6/xlt1HZqqqUP4q4Abr+GKwofzh09dnA0Ft5ImO4lUG3k+tOyGAjYREFWB2
vIwNxt52uLqZZyFsO63WdO6iYR9Y8hT1XrtC8ANHcA5PwDdjQBCfQrmI5eW7Fc08ODx3zB4Ev1cv
1+xpfI4uDgo8FmpD7ALCK+YOeN+StjIISI9azMr15Ax6AKVJ5lF476GzPR/F7wszsE1wrS8wopj1
U6yH5N+4aZG+H7ZQm9K47/WJIWf/8CRi7PeFRQLLh0+we04kjrV5VvjYBJZWE+OQTZzs0NxNgSl5
LzbMO1J1YdDVml0R43yeKZhdCkZ/SFW0jGLN1E6ebwjsaYU62X1Z0c/LMp029TUOa11MsnvCcmcx
fL563SltlKfzsjRySnFCDtrWIT2pbnynOUlWZ6jwJVPnvh/PlMQEh0hcsYxFXaSovgPlwLIvitnX
2Fpg+H0NUZTRFxSs/2TuXFf26dCn1pVA4JdhiEzzs3PZzXKdhYicvpaVqcpNVX0vAFaCQC/dpHH9
k9EYiOv4qUIUSQR9ekzbwK81DzhYVVvqv+FY6H6X3Nr4II2LtLH5A+1ZIyAt65GjQDUYcbl8NgXQ
lzwzc6YEWW1fIr0SuoSO45XqIrfOI9igRHuDA5zIqhsubZT5itahQsuP3WQFIn9I2LPIioLYQrk/
qlr6Fj6POuVrMGlGQd8EkIOeTkbAHVIfM0h9LxgE8wXiDAJSnNoXoIseVoHahnLxiG1vMdXFflys
asCOZC4SyJyDD+LiEEPqmRl2L0nC58L0BavTSqVv2h6LcgbyXIiM9qMNemBZvWLm4qpGqcZzDBxN
W2XBPntMxg5neKlK3aoqgLDEdoOqlizji5Gn9tAKt19az5x4+VpSgokSDZqX//D59S9xHNiMLnAO
5/CNj9F/AVFTLILG3Gly6rYuRm2AcZ1Yj+Cea73CE3gUOINYed6wcV0xsefPXmmA9ozggmvWdTwj
AMYNLcCpid3P2aqYCyb8r8rUKx6mXNemuMxHfif7Vrl6ztarZOApDbDpvMAujcF3Z2LkhS+h/m1D
rE7x6TReZv2iJuG8GURTJHrGwPzOdNf0PTsLst64NELfs4GDl6I02frKvd1pXm3DEF35hELrwXwa
OCJ40t7VxF+A6YSUbs2L1ikWnR0rG58rETj092fdi2GJEi0+7TusCvzKuZSfIR2YCayyWTkWrI48
Lixxhf4tHqUQL8G5CrgWqH6P3POJ/AZj/CedU3j6ofUF4y0Ls81mqja+tZixLTWGd0sIy+bA/ctK
AK/vbeq0mddwSfT+WXLRpjufDkv8MyIEuR5ZA2/tPI0Vmag/UWb2Ck7HWlr7xS5M3ls2uYCh53lc
ddEiqw3Ypo4Ehkwh/7fFsmsE7xxHFB56Yf06eCNwO+6ij+lg+kJhhNaq315HnX6Nl2rdbx/XZeQM
zychHSelKa27HmSKd1ptD6+un7oaD7e1F/H7UKCJEnZ4p0YjOHDlSunfsnmFi8wUmXa2tBuXGqtP
rE0PlVh+5SCL5Zq/kIX27bgPcqvaxIJEwlp+os0LJ+YtI3A4eRtmyeIAaAvzQzkC5CLIE8z08MHE
PUPCZkMuXU1QwMavcGv76LcwzsPWkC9TH9+0RAkpofKL46PLCLDIiRwjfYO6DiKIvSjKb+7FfoVU
iT7j4r2FpuoJeloPIWJ8u8XIlV5qVBI5vEyeihBp/yfSDHqX9B3ggxYxf6qLLQ1759cSUHdNgi0G
qzgw+4RnjYKjOEdHesIk7cbA4JPd5IWLLuripzpltX4qpX0DgLgULIqgKi9A4R5FG7+7XLcilpyE
/okNsX2Ftsh5oRgea5xV8Ut5HMkofK1wG24eT2FCSxRbWl6UBK2rQHQyAux82uCLhMdnNn45cv+v
7OoZH2vlD/1QFEM4JL9RqpAoHyRe6+c6nzBfSBiEj/PZyi1PLCU0scKzs27dbv+LavmGCEI5w+wE
0awkWNHxraONs+Qkl881S6kmqXZvGC6XdkacPepsPglzp74B60C+xENdWQjg+m5QBygAmBJ8O9Rj
9W3LgkI0QH8zRD3xE9dHXwAYO1j/jmkz1vpwsA8PxUVX6Ze2CKgHQAhPLB1ea85E13dccWlWXTOR
3qaX5J1d1qz1bHKLaTonto1kw7LQQgavGcWKbBrE9/icH0Igr8I3Py1Efbcx27hs2+NhD6qJv5d3
MACxO+B4rtQLjHr4wqfLCYwlB9dxqPYEo6iDmANwL4UNAxKLYHMdq/cneMwPAgrXAJhpTpB+K6IT
wS6QTh7vhc/kTMcxTJqH985b8N4pbUOHhdHrIEBOQ0t3dhG5d8ghBqmy6R+BmVRPidI2VWSg7N4V
SZw9VV8TSw27oYlyfcPL4GgZrI3pjpB2Gjcr+BFpxNUiu5E7RAKbAABEOfDo1Il+voflsjACrI8m
6cI0Yj9gSs7lI48IXP0v2OrjhMAPtHvdV2Jkrtn4XHEdWjwYNJrjoqMcbS8PDZ1+PVJ1BIFjck0H
YXRL6MWSmh1bhEB/je0+iGPVv1yyVe6veD6kP6/C4n2m+w9kzlbYpN+KmUKxun8A3fUgr9EAw7DP
yNxnrDJv+hGj6DH4rGW8pIbT8fgtWzD/xkSZyXCvULXidYqyLUAW3x82KC9MMKuAha1lcv/8pPyQ
Bqp3BpSRa2x2QwTYZfkuO+XOtcqUxjAztFE8a7kjU5Ev6CbdE4rKuR6OhkXJhFZ9+L/ngw/JaJKC
HtCjR1aL9vLlcpN4VfPWE+VjFS39+bOrCQi0Oqo+kYYVzgVVQr8PLsBHqdASB+aHGNdfAO+5LLIL
Nr8I5RkZkeW5mG77GimoPEVdwrZsxi9dJMnWr3acPcK+giFt1dTKINCCBAx1JUDjYJMnz5VuG+Ty
OvkPS6bOy+czb+j3Vwn9CLmHtc382n7IZHD5FalxibyO76QYoI0L5qyX8zH6omCxBfJNIR41qerF
O1+IuilOd6YKKmNi0MzzHZUD+rdAWuYxiIp0bdMOa73M6Vm3fmmKopafrRfLiU2sSan4+KvFNivZ
57O1v+T5CVB5O3Pn2kJDgvS7TUHltF4B1FiLHOeuGwfE7FuRC/n7V5scTG0Sl4TY+uIkYDogQgeP
gfLYn/tsQ0NMm6zVxavXofljcFpqZvndo3rgB2quNkJ3+sVKZKApK17Rnck+EO6KSrn7DVmBAmKv
gyjKa/ykWuQLd1vqdeg6IA1pUOiGfoA9FZGSJwh8dz9Yf6GRBUD/bn9Q94zWpRxFP0yzLWEP+ppV
u/3R4hiZZ26BwkJFHz3gZhgoYt/hyVGGvwKK6wefbKXTvnXKLBD7lB7MtlHh1sTKTGJqL500WPyu
/MgoEQBIudjuDCKqlb525jKC+rDhwFGrCjxxhZNbSJvQJ8sl0OnUud1pjgmSV3UpR5OSOyitznEr
6JHEijkOSJRe5am45Blm6OrHvmo6WWXA74ArgX+yQHmfrccqWlXcCRZxyOfVx9YHPWqVJbhPxf/x
nwzyZ3Pm1ymkHe5c15R4ee/1Sr3RKW45g8U8Fbac0Tngr5R2RA1qn1fOckISZ4lq8li18VLqF8RO
42ef3elpJ38k0gJ/F2/fDnkG2IH6nR/7y8dHn5hYkd4ZP62F4OQv3QYdthbEe0lSzVhssw7UqTcY
jON5Vnu9XxCgXfF1OHzjO60iVgx8JdtMRG46HiEQtHxJhLS1IWH+dqHTJ0LTv++e2G0+uxUNPNaE
dms4fjnJkb41GMjNzEpNlh7xAvVr3ISYkxKEuteS1I3ShQZY3eOK3YBZ+EeQd268PE/huUtzHwnk
POEOS6M0Vq46l1Np/+UpDzOkEGMcJHbyDTejllativUNtOHsO7uZ6ME1r9XWYjvx2uSI3ylxe4qS
P0k2utNmk/we2VGpHuOTphY6qHCV4EMy33YHavoC3YEYXnvjHarAGcUag0HeCpJnPGXdZQydVTdQ
gLqDl8o5lfKq/heD1JfP5mGlSt56z95JE+mMvUgmP1YnVKQ/BtaXAbf0kmxYRSdZJHUxfgZ86zqV
fpFQlrn31F2JIjms6W1z3oNREHQnxq7KYslT2iLEQjXTuzLjJsYQNpjWPonS4njh9WkKuwdcIvb3
v0bOjZf9otxzxW/Sjs4i4W9xgD0zlLzX+8cNEYxKUebjOO8JGRS92i2NblgjlBmdoqUx/yMDwuxo
i8MH1GR6AQohFJcyQtzOUdPEGcpUDdziObi2vwRbpZhMp63K0qO27Cm9MWpEeB6IJIQrJH3YDQq+
mt+1jJGPTJu/3814rSDM4xksA4Ezs8m1IdB91dRxBEvy3+5301tUmeMd+HExg6wq+azupeYUXx5z
RLD5Ma6W4fLPlXAr2lI7iLcB/f4yh3z8JwQmXIfqPQmcakGyx7wtHo+75PPOoid8gOjIGmMh275b
fQrCD+K8LtiB6S5d8yWll8w2AUr/ZakePBnTRj5mOWAbW5xWjPN6+GCR1j+CTilqY224ys7+32+f
yZbWs0D6QLAgm75qAZSW11SWXXJr0Cbm2uegWS6Vhl4ZGV+MCLEJ91WXTB0TCT77iFRNiCQHyn0N
MPTs6Q4r/Y/eJQdEaEi0LQXfIUhGmGQAooq5AtPVhZppfEkQ62OpEplnPIV8i+/zBhLuDhpuATVd
4FX6kf97Jn8tDn7fzwwixVDheIjig0qvqCIkFr3wgSzrwNXQEi+HUI/M+fPuaNJM3MgAuvosRIde
3200OkUaB1+uck+/UOlQQQ9pQCwguYbZ+dZA5SzMLjFV/rA2Jy1Ql6xTH7x55ATK5mYk+Qtauxc1
Alzv9Qjnjo2sJxU9R7NlegUV80Cgj+gZbgiKSlTOwGNjn08BzyzT/6DGjyTVQLWt1l23p4+iu/76
/T/VCEmL0/rJTxxZqtqaYBSs86zKsqvIv28ON4NJVbY9uRJUd1OY0ixZLhIUFOELa7rNSLEtaA3R
7U3lPKqYUd+rZiAateY3K58WvI23kR0qL4hphZLmB+Lr1sjjVTZDUaEpsvPsavFfyNFOOyV8x2LZ
8hjBftVzmLuRHqOfFrCVsaeiBWAruSfcsLrcIiWolgshBTXXPJ0rPr29cNBHNrXn2S7AMuk2ESNL
h4OxirHXceDf8nMeCQ+WLfl9Iz4KTJ4zBEH6r3G6CP4Kcph6Uah/ikikw+c/ExA8ghL6ld2ADMpn
dS/5fMcwiPYKpPs1tpgGcUkdF1rKG7wBaMTJb6ojE/neoDpoVmSAe5npSi2a59pWs9izr8IA066h
3alNwIPBYul8qje5TFxaWUMf+0UtkPRbRfVu0SsH/Lh4mL5pFYaaRKK6RCCMAAuvWo4iSI1CQ14a
TrQpk0ig+F0UH7oMzr3C7QjKF8KTEqHZq717Ce9CbHCtxAwziYEEvqgKeTlWWMepYJBn2T0qdkI6
71ZBZ6b2YxM13utmhEzIM14CSnpQhpKeXqdiFxhvzZeiacBlGTzmDLiyyMz19ntoJjV8UiCjABfn
CQe2RrmXifDNyzLRjixy9RG6mQhIZlPrzIJCXxcBqNaPl+vBtd4E0ceoesaJLRqQaEu5gOBnAHNZ
dxfqR/6eVNIxl3qbYOFr2WSa05LBCQMT8JerP4aE/B5DAWsQAJj1/nbx1HhpwlDljdVfpKfBxPGm
xttDBjQnJYHruVqy2KaJ984yn6SF3914OCiv4+aW25riQGD89xXwKusfTl6WFvomt0GclXJ82BY1
pmOtprngsdJuSIRTtwO3SKdVbsQNrDg+/hlxyJSX1kj846Wj2BI3vylzU0tk74TFEMbVhPOxZ4Kk
6lVhbbSVxVhNmH09JaP3GuRMZc/YK+LktOKQYnMM3Pc2I+BOHc9eVJ7+XhDz252PqTcaqQgbIT5v
0JtIUXILAhA03LeUzn1dmjQmJ7FIBmJdNUZztfrde8pJaFrlKbcmbWM77emqycb37qa4iEX2VE7/
GrVPGlUAwKIR/a95GoVQtjxJPgr0cBQgc1XMuNsP9Fy7q6rSUY3dmMNReEEwzViWbK75UJyY9Dep
4TdMMpzSHACKAcU/u+z/X27qSb8pqCYGROi2TDsmdjgfVN82Fc//HSCRHXGNIL6w6KkE1yWQEAgw
8jO7cbXGZZuOG3rUliEkxjwHWdiZV7Wep1j+ho5pFc9JftzkknGyYG7D/+jYw+LkgRUJ7AkSfRvs
RMPBwhsry0xLVwRHbPtoCuWyHtxZ1p2GDmEG7mLay4LhTrFx//SPRCHt4BshgLVaNZctxGDS6RWg
IWt4WgX0t+loQ6zcYBj+xneQ7LHUVHwNZLRexHkx/JKlfukq7g/gjVnU6YiseHZTtwWr5t06vm4v
jituyPcPp/NzgmJo82F2L0e2qkHDvpWKSTIod5lIsR6eOmRVQfE+7YEjH1H7DuEt8Ru93m8bj8zF
erZlz7eNwtl52+3ERytpq5MQEQdJ+ZXf3/KCTI8f8zDWXTpeWVnIQ02lojGEzuB2tC7s1RxIhi0V
HThpvhumuDBOWWC0DVBG2KKfUUR9UCx8L30UfGi5VinsESHIihgb5agQcY/HPcfBOFknhYrZ4GL7
eBjIXMMHfuHGToElaqpL04tuWTLbT1oMeLI7AxFYPhpmGSNpJbkw8RLGnHnEdTVqa8UjNQ57TEQS
0/XOi4uAzrttP0v9Q43bzBpPlDsno2zr7W6Vub8Vcx/IWpGrQyj+wNoWJANmc/G25CP5eX224AQr
2xNBuphwIQ3PTS1LhaY8JLjzq864Jla/KcMFiww/9ZrBnHYzX7WiT2l9msU+FsahgiFt6FQAIA3L
H0cuziQm1bM8yPaf2ZA3MWUQLGJQTWmvR8H6V3TttDfMHWwffmlWn6CcjazQP/jHyx8YHusi14Rt
fwQSNVB2JA1lA/HLmZuh2VJlMbxmKa0xWpNRllKAEZzb24pVRyTHeWp4VaRtGfM2RAeBTua5hs7G
OBfVdlbINKOegVwHCr6g5QaKi12GeyFxoubc59F70tl3J3sjlNt1yu18kd75Sgsr1qcIwPvFoNiz
tEGFw9QdPkAb+LNwyElPd6cYP0nQcJoGQfOuSgefzd0COpx45rwzIJe0l9MZSH9YSCms1ZSPoHqo
4qiJ9xVYtEemsJN9x3NVHNusr3OMeihiNdiaIYeVYYlKVq7LTfICu9Xf/9Sik9UxCswBOZ7i3Wlw
ISLbs0aiLXE3INKu00BwbZfpxd8XOaamUCTPPX8fhy4q2SWNowvOoacxgXVIQrxazHLqGXnTy/Mp
WMNw3+V3VAEks3el/1QUKIs3gnAWvyqf114nlcmzlLwn7nBjd6Kkbcr2DP2tsn02ZtW6NHQpHdD7
X/6N0R3NVollg6WEAq9nAOLXJjQTv+UrDb2m9gYsaTTzP1J7caoZ2ynVQI9iEzVzNAuGsZWbZhfv
WTe5Sum/8S8wYbAm0v2dWYP9l442irYc/4WZ7eqzLyYKbxSNikYP07B49ls27fH2VSLkjiWj1nJo
AEEYwUwCDh30uEiD8Hm/FRgrSF6kT80Rpl1ufahX7/2dHftpLG+VtxIXctVUxEOA+9JYcSVsLBuq
d1opV4KxRff8EO6pYGYeRLBrz6VO4DbllDz+DjZTXG2Efg5MgRojG1SfE71KG5sWQgKcxCHg2ab0
nQ+qDP55CLM996dSLNW7zpd1i+IlUTuu627/IKvmuDzwdvZ5/WN0JaZ5vIjKkY/9Xc6xn3swBgur
LftPn0dTTwW4HvKwbHesVRJYivoF7a38vO6CFuzp236+q1m+eWRXe5LTRMYSuR8qigWC3b4hltUR
8o8QvG5ZpKGsz++SOJ7gm+R1NbJs7ncmvFqpEy6P/kJM2eZuHCTeBePTgYaKH+Z2v7ELcUjItjZo
ZbHy002Z6Ak3tKKx1CyV4+6nC08TJxWnsLabH4pxUz1fnCo8UUEbgwcefxKP1JuMvPyxdvYCyxbK
cQlN/yCPgw4t1zZ+AuD0XVTtMrAiExAIvKlXZGY/J7tXOrGI2/hQiyGu3HClACavJufhoDnwJV0d
EgHAop4jlqF6ieQzgHqdSn0/yiE3bwskavLbWtSvdmcEX3ZPOvj79gDN0HuF+YjIXEPp5nAsJE8e
TDVDrqRxVWrEmuYgwLtWnEZ04ZK5d/5J1nAQeL2KOYnfHo4tLTW8+xP5AgYU3vHmxMq0LfhHNgCo
1ON6/8rs/318XLxFEJKHaBT2G7sIx11R/zH4oydHiIyQ1MTWvSiLlAFiLnUBZa137fMOcBf9+Yq/
auNm5cjwkZCK6f4hYqXyNeXHQcISKzIRUw+am8eoc8wBdznXzbs3kiCWWPzs1R/XBoz6e0+SOs97
P5RWSI664WWGyOybdJEmlVBl6fTcrFQH+bYxVQU8faAjJ8PuVOsWQu/lupOKxUVczgnq03zqk415
GaI9L8J6kK+c29u7lKk2DtI63FPdQZfp9NjVHrC16lZ+ssAHg11kW5vxgDgegZXO1VMrRISP+JZH
jDLGfteExQsoRW8cTEu4kCuN25c/+Fh+gnTC2v5qwJiqwirPyukg4odfBtB64cDIgRu+oGpP1N+z
aGzLR8CXZQ7rVW687B98d9/R/dIAOooqabbf194hcMD+dBP2VmgVAGfgykN/kIOM7VuzEhhR/FNv
6SYIrIApGtvk5L0ou756ssmNw1CJXdRYZ6FvPiDMWkBYxRB/uKJOB0C1kBBENjYpWxc7ddXNFEvn
55LGCh2gQ9XAJfmufm/+HXy2IYs38A18xD/WJnUE6H18vPvs6YQYJUc2/Cj72b6EDDGh537m4mLq
p7eGrfbQsynIpkEczQP6xfdtMJuhT1i8+i64/4Abr/KUuZj43gxq1eq1Cs+hRPfRTgKkXD4Z4cW4
tMjjn/kZOcRMMwycZgQ1dpBEoccM467AM+xv+j6lYVOEGA6StoaiqPkaqLQZfcehiV1aWtPtbjz0
geCGKncUfyZjwnFT6SVy5DegGcbNAKRfyzfcssvNls3yFHWUOczv45/kFCq+VQwcAmx0Bd12o8jV
PWCuX61zRZ1tQmRnhcTgFiV0bPs0eglVxRxl6zWLlcpWci+986ZAmEmWChEeD8RreUYHv6Y3Urjr
+G5SiReFnMvGYiEqbZcSP2Qr2IbFsTbuxg4pu0r5/ovtsAtF7M4DhCxHVdt+/qUkOSCZ3ewNPoKS
RdytQcA+4lvl3fPqyNauVI+gRThqTaO5ZRB/o4PorPJsIFc6ioISUV7mhhntxXlSyELsHZKbz1PH
WVa59QsUcpQveCcIIGRPY9KxHvX66DJkrqG+391/d0qk8ZjJejXXcFse7WI9o7S00kR01ouVF7PT
A2/FsokcwtYQcRBGljYAzZzCsahSNUQ8hLr6QKC8ZbWgtBhOonajci2/Z8S6qm786rhy4rABbymo
qwptT8ye9hGhJM3K4Ml76fFN/yMBM07Z7+4sN08KuF/o9Cr0wn0EsIEcrsldT6puJxy5LcmR9faQ
y9qkILM1lrOMCp0tQvh7F6QfgZ3kqBbz9x3r7OnZQ4iDo+wh3BGZA1IbvdmGplgiW5lsRrtzdwQk
vyBd+KQSZTXHHTkg5cITqIR7yzATzGlMqIgUHEPIR4AwRdnh6Lg/TwDNlfSafgPAIAbIBI4WW2b7
NbmIiWITRpaD39cSd2qfesfSQdEyIKPvT9fr8BKcpxnJekINRDj301aT7V5fRoCb3CpTsGwXLiZH
/CeFovRA8De7+Mh93mN9sxU6Umxtfvv7FCYhOYqy408rAvvoWNs9XeAK+rpm9W9A/bMqMcXyxhYe
943uLTxbtTK2Xm6pdEV4/O2v5lLaI276KFizR3ibJSWWYzvKQPpkkDBeJnWINEfe+irZWR+DKEy3
pzVnKKQnIAWRy3266XtCb54weidfrf6AtfflnxfAw+WwhPdJ9T1bnxQhw9A5856gmIns/gkkN2XN
C3Aa69MDZvVItGYFjExTPwsWeAkKTpyepFffruL6076FdczIBagX1GiAsRaLIW0s10DvjgP4YL9p
DD/QREATvQLNQfGmgRsuQOh4zTgWeEZhVy0K6Jr5aTK/TuZApMz3Abq5GANvL4wMgbR+Vb9pcF+f
Tl/hO+M5N3h4UXl3A8VP/uADP92i5HaGuWzGlbCBGzM+Pplsh+ZsXLuuWMP1ByrKdQJLWxUBBQDi
A4bT9YQm4SY+FgBhXhTl0dHUG3MdFBP9NYU55MscnKYZ5wozz+0C+z8ujnNqLDVAkUl1+ozUlSvB
gbfOQxD9+n7C10r0dXCyhUGSFFZdLFymV5LBUlLAH6X7Q92F6D4XwSP02HoG49VQkcGI4tECUHET
/JJdWwb12PtY89FUriM7RqPVF/nczCVmVj8yT6d32nyK/RkIcVSQ8EPjvM3LBlNZlGUPfUbRrr5/
7FjfCIY6HnEyKpx2bIsHgDb7kpyE6uzR0jTMm5882v5qd4D59huip6CS3pmuGfYhpGIgtRaXnQgC
qsqFCyhKOuzK1Faf3UUqmKjD0tkRSQnR+nYbXeTJAZzjGLlPl2ZkXjJT0LvKy3JDy/mwQmb5/aPl
qlpzMmh2r2NMY1IPhgxrcqSvAdMc3GdRNRf4Ll1CwvkWbvLJn3qnundNFzj8IotQwyAv8N8dV3Zo
9pdtUNOeUgt3anedbOvdVD7V29g+XxlF/DA9K4kM1uH5RoLqsJIxvBwyXESgucfnnK3yAWpKXRrR
81km12VAeLiB0RvUmeXTHPcArC7bYKwZH3sXmCMCI/17QG8cQehIczQd/q+mDjKr1onvN0fDgqvt
G5M4W1uMOzsi4wJWsCXBQ/TedRFoPnrnGvgml1WuX3pkRK+jtGLF1oYSj4VRKi39FpaKrVVW7S/z
VLljXHG2eD87VmxGQXsl0EuuCMUOwo8jh3VAti4hO4kO5j5rprNajMM5IVLvVR0sx8xI9DB6PVAH
6IAnmWcZalqeor8BK+2wtezBwa/KGCDh8TgcAHhxMGCiNaanfUuneeHqEzsJsk/hbEhBEV6CVNdR
CGqUYP+cetxb88+/z0qsjli+CoO8/5msuEOl2n6fLKs576F7yV12PHUs0FRoKDBwY6jLSvDzaipt
7zZfqyPO78bsu89FzU5vgRmVLW7FnGMOYSwGb5UU8sF+qaE0EZpFguL4RwqsgF9agObpnKSsc3cy
0rUpmyJ4Pfh8dcQZtxoRzbugNabK1iwB2G8M1HnHxunsTvA1wbISYlNtxwFfgd6sNojOwj8T9RVc
ozU80Uh+V8VxRN62qZKak9AywtryIN/1hYNX86tmfJH5m1zUaUJ6oen1qHnoe4NAlz6RP2136bnH
DT7nxNmNmPcw7gMN3QfPmBmSE7FcQQr9hH/Qx2R0O/MPQ2OcH2NmrYfNLWH5ZTMUChhQEHbmg9/c
4cbeurmqqicn/5CFwvTaP6tXaGucKtym+2O6mHk7JBQ/NyBqG/oyClrSHM9L0BvZGWlpo6Jn7u+p
2e8irMd3f2iQDOBatEki2AXxY+DD0s20BEy4wOMhN+3PkeILanQnJczKO41Nj+dBs61bVSJjF1s1
BMb9PBhCXHtKhMAPcx2LBbq+EDbZNlElyHJ0l5lZdEiZ38ix3SmGhZn6S/nFlfDTjQDtoZBt+FoT
4X9lwt+rvLHH1uQ747PLLrGYR5WWuy0R6YmSaUHTQS65FlL0DZXB1TbKAIpq8rEZ52rswtbWGxus
G5FAk3AK7eoe8OhVacZ06GbsTKaiTSmxgBPPWqaUawwXcm/e7gTzoMeK7bX/KeFOYfb83N83w9sC
/R35NLnF98oAmCI9+Xc/EvfTq2V522zA6y8sGZUoaUZn2XGq3WLghgnPGjXYcZnEuv8E1JiTg6mj
b5T2ZL5PxWbOQOHxrVn9qjoX56Qgl3VyO/Zetuih4BUU/A4FVjDF07z0CCEdy9hXaBDCW6G8kFUu
csKNVb7lyFnOKQ4rqzXbUjAjAl6NiKZ1GNUCXexEn617HYowOrkGBdaI5Z8fEwbfXKZRdcqiQ8K7
mQtuDpXlTQDRkBR5Rs87uaW1JZzPyMVvhH4/lHRgjJevPurEOzSGVEDHCn6ekG6d86gNoxON10wK
A1lGVClm2Xl+JBX8bHg8W3srDR4VA+ytfcpYSCjnpiem3yE2HeMmrMIvItRB43BeqIOYC++sPyK6
/dhsHB35Y3r+d9mYNCKR9tGc9vpqjWD2oe5zWKZjAVGtxoQKffzNB9FcAcpNpio33YWyl748I6qK
KcgrncqO28tZTIgJKelKDsQlcUZbnE+Egf43MvbOdzZfQ34QqW8lR+bTTOrmNYNAUk/p9nnLQFHF
smSmKJC/qSw2kPX8A9Sj4S1EW1EupdkKhR92TXuhB5BgEvsAhlGBqXsRzZrtLKFVSSZd0bHHliIh
6oQHc7sxmNsx23UKkv+mYcc4RJo7PLxl3gV5iQiFV3qDIHVpeVAkfQ3KisxaH8ta0+v4OiayL+7F
80cqu5dJWsm/LV3FF2bpphSetht5InxRmYQAFcy7mD0BiRQybPNTeSzmiIw4PTEd9+tPMoZwTgdg
9h0Z0Nkxf50514cdiw2x4NP3xvZe0XWfttJgFMdJ9Gb6BkTWrhd0FClQ45F7FVJDmP8OtfB7ptn3
OoWD7+ggWczH6ldVidLcYoBEjcaxEBkXDZ5P/d4Hh8JDG48Q0IrR0sw7aQff0G/lepsg9RYeK/0F
YAwBVneBd//qvw958rEXgTGjcAXTKWgcLj1IeNLsFQmTLfNKj+76SqRo1+u6EOxCHXA/1q1XTjS7
XohSL8Z/UeWYJVcjkEq2kZ+hkg0BjbQZIPJm7GW11uEkA32h1InyUcKtj6/b/i74ECOWbRFzUMQm
sO1on8BO3f4rFciIh2M10xev62cGvNt3UgUpMAHpWbD7spdJ5yN2NlK4EDG+QyGCveEJcCfZXfL3
cyxOH1PBrrrLI/QdQuTBKUOosgFb0cMo+XBxWWVgiEOiK8DUFM2qFyJ9zkl0NihASmK6TkbXA4VH
COpHnyJd+kEWG8Q8cGQ6FnoD26W571noUhVKZV3UvfGq2NGaN9d1VTiHoUcyR5OK2UmhBLd207nE
avpXy4m794YJH0Sij6wOHDH/B9thIXlOtNOpRVC30E3GDPE2n8vUwcPcNxCTeAP9paSgLNrlBV97
DyYC6c7QVkdc7lD0cVO7f2Uz65EHfvCz4kF3kzvVwmMMjLM1gaNC2ZaQY/Y94qs44+Fjkh5n8Kf+
jYaoAAeQd7dNqFBWjOFAR9RbQO3f3N0X9qQts7dd24bPIpN5RemExNMIJCW5PBU2R+1tNhvw3Vky
7gVqNLenS0J5x8ewhGI3vnsr27HnH96t8VbHs1lQ9CzZSnan1ZkvjZAz6xztxTHuknJemAFMIDY2
wZL1qRTXdS+lfMYl76iavqgXl4ru6n/8kVt48a0HdCUCjEJk3fgcR4tTLTdyivV4478wMLvN+Mzu
29POXJw6Wzdr8wzyudefh1BIcApPY8qPFfZgCSR4TfmaIbga29wONOUPTLZLfr4/y0oTiowgXwth
gFXrRDD4o+jK8nerDzniNreFuhLHXtSf3QbjonSLLBsbbJAA7ifPWPoQo7/LS06BIE0Gqbhcbg4w
dKZF7EaVCgalnDwVyQjeOo/BeKnHWfWFZUhEC0EnjRlsNNVwZ8OStX+z0IKHGtxNZRUTgh8dY7Jk
cAyR76i84i1BAyrzDULhNmYVuFjq6ITJHM7B53eNPNGTNcOUjQhnRbRhXk45jOLUTVoDD7iHFVjv
fZA6sPvV8ucrqiIJxol3LtKdS/2SWJEO+I+bzNBiqNBRbHR7Y9R3R0xqCt//yl1SC+xKv4bmB/Qe
m16dK+BNd+RA1UbVD8ynORYG7cRBKF/MhrQB6J7qkbQdp31LzbFrgR1VR+r1zKnNw1FRyu/LkToN
7LqyLNoJu16GdUhqkS5VESFhoMbHzYjGSOH8XmsgZLx2gPecXyQx5WPxG53/GrCas4Uu5CGoq6Ee
kOztG9cPdYaBBv3fK0F4rbTFBc+UfTW8UwFB0nPAhXIcIGSPwykJsyHMaqcXidgBK5I7Ta8YgdY+
Y/uUGmuyDy1RF1uJXq/3UI9bIntMFK0CbU5YZoU71x8uyKVYGFb6FuaRwBSoPaMwYQjKO1KZuSx5
GLRp4XP0NaaywdtAvpnhIsZAkX4XAuXEd1puJypjUrJd+iyDsJ7PPBz4g4NP3eoz2OkKZjdaNxsP
kzelbDfnLmReGs/6hsQoIUnGXZTG6UK7G7pAlgYxX9T79oUePv/IfP+zP9KN7WNVwD/X+p4+CYkE
kj0ypvoUr4Tzb05FaSG9FSfOCpY4XSkeLyZq2qOiF1GsFEke8OqobaZmFtdKBvgK6UMZ+NzbtAlu
CjJfED+UatuUUQge4HneyzzKynQXJITsYcZ7Xw38ehBmtZHXxhIIpBjcyqlaHUxufQVhtHVStp5C
0YTIQhR5nmnqWct7YLo5Ejl5dg30c4ZWfQ6/GwdcTn9ZLOrxnQH/V91i1soxNjXZS1PTBx7o9m5b
3eMYWXlw1MefeVOM50HrO9ZghVWrI6+O8sSfDDxZpmQGopf6vvqesQR6InpLLB956bIaugkyJbCg
i0unZmV6iC/w+ET+lAya6sk9YwFj433iKFRVP7bTOLVN8WLZeZ3qrjEUIvER49lK40qZoOZ9cWyB
LaVRcZKKjENb9L6f8pfo0C794XXHgAelKwzW2xrMZ2HTtiFB6VDzHiPYLiG7rO4kYggJmqAE/Yw9
v9Ke5vzsEf3lsNysR2shSeyzDroQ5cA7+GBfoOPfLbRoKPND4TvUd2jirKDu+/TUZcWzIa7zQm6b
eRP8XjDplsQRUkYFnrzuQUyEb12tBwDGqsyEyYQ5zOW2tb/5FpWHrowTSXbBeZCa4OvZiNVz0Ne7
9u2E0zV2myFDMSu4MmVjTtt4k/oYlNEhyba30uwiFvOITAiKevn+Zsimy3M3m0n+Tsclp8HYxo/m
r7IjDaOfrJFRocYkN6PIJ1YqV6+f0mcxe1oi3LAdNlMnYNWrg9qUnLUD8to5IghpVQy9MXsbuIjA
gTUnumuYLIGsU4FFnLvZseaF3Inkc/lnHKdbnWoU5KgXUzkmXIsI+U7dl3w+h3CpoyaL6A2EHaWH
U+RYJcJCIQFNv1aTMxPcCkzH8HRaVp2q7ngerGwgeN1SlIc9ECt3+SjPgH3IGHpEM/HhZ4usV7UR
Vd0/51amKJcj4pvL4zGjvm35zONUZtNFemqC93koA6qPYa8ORis9sF85yM5H9jph5H42lAF/dblu
D6e/jcbQNqsUiE1lrR4YjioHjUTbhaKN2XCrKh5kn1H9NaIcUZoFuhYkuhoa1kFL1qcnTrYS+i93
K4xRqDlsrsP6ssIlLeAgCmcAtwpvIkoCL7Y1GKAmHn9eY9X5VVsj3y9hINewcXCF1fb8T2Ly6G71
UfrgIoCMc+ZB/TCG9iXBK0x0sIS5pNolYqy7OIzsfyMv266qH3JsZnWjUmIfqWMeSsGRJajt78YB
xOiA1QF71KaOqo7gyZW8Mr9vqVD2A0Nio6VDgViwmGOgAHV2+8XpfHBJn8Od9pESmy8qWyS9kRIZ
Vh78sSL4Ae2SVAVZPxXj061QWjZ7MTh00JMtw+xehsqdujGWDp58Kh+38kixJv2ZmoQnzDZmIEra
ydAf50W2tdYptddgHkYeKv1uvT90hNY/NFHaIqf5yJww1lL09tzu33AvElWPDgJPv/WI6vd2pzJB
uDCTINXaVUVcgPTosd5G3Iq5n9t3QQQX1KquCAtfaijoAjfQOjPUlVYS6/j3wpSviy20fCdCtyid
ZIb/SorAwJybAmvi8DViEM3JW9PZpHVHA9fgcQH2Jpz5RkRaEW5NuEmbi2F0SJmpo7xqxvCE/28r
B0u0ujgdI3yaZ7dfePVGHDZFn+cgvo4lBSFAbwvn0dMkSKlWBJeYuR6Gk2H6oK5IyxdAxbyxDc4Y
Qy4i5aGIx67sogon63q97bSuJ6EbJnLstB4xv/6G2juyVzU15+kOSThbmtJaGVjc6HbpHhDYpxEE
h7KuInYSxDdO17hH5+Hcmv5KUMGWbA8GO7Fpfy8VFvFbzbqeJbElNv1TKm0gVtPaOgCDHDYd9C5v
FFKggo3+WX+48EqpIauC6ZCBuMXMELc3B+/B72P2ZwUxylaZTYfvaAWXq+qzC0G2xwfIQye7bNra
EqOcvWyJWLrXl0CmH5tPbsA0k5XVGcEgRtD2uQN2oQhuitpgUpr5GV6BlicRsxDR3JNEY9vHuacG
sZVybX0UUTPXWo88jx0/TlKHzoPFST3VhVRO6wQIAfUKAa6e/MNVF64I9S1XL5i3/K0ccdPSuzU1
LARS2Zbu08qAOiF55WCBspMAsSXMzKderd5SNXmNqC1jHJp5aKQJIA789ewDosXcrBHBlhs0A8pW
AQ16qTEsXwgRgFH8uSrPKrzpDI+VhJAGR1MjBHaKkoJ/dA+OT6JuENeyKWWziYu84+pLBUPNFsOZ
UAHHtyomLm1Ic1vvf0bwpIEMSCn1pUK3nr0woCrQiY0/10KTKjIh+SV6tazcE6ZCM99SXI6GYuR6
L4cDCIwDwYBF/omvXQOLstRh7pj+zsKGhIqKPorGMVhlh/5NNe08tcr954l0NVfTHzZFOw0b45QH
1bD88exHBnWFUHlikPpRjuU/1YXoXymheDwEiIwlYFVM5pWzsiaw9YAfXJrtIfrZCKEgxIB6xBFr
DszqK+SQpVmC19ukNqK3WOjYtxCjrflUR0tdkXfLfJjFOc/s0e4YnFscYBwNfobhr8we9Rj/xUg5
SsOmQdWMLlVhmtEfdFm9PIkEzxT3LmxqMubXN9ackCML4fZK/ZBfNkV4b+6iMWB8KqG9z22JDwd4
JqeldZSvR1jqDe9br1/dDmsiMYY2BO2uqKy1PS7x1IsiBkRcNPavQz74GE6P57mFK6jffx+M76Hq
a+Nt1CvkGO9T6daR3hZBOLrPNGW/9DriOfOHTJYfS52eTHPq51vIyr9L2AL6KDR0osNdlD1tCAT0
BES0zv8G521/PrTPcrc4NbnbAxZf2/stUojS4UdjMqsGLbWcJPAfzvgsqNCngPst4dzqBlc0JJnW
/ead6L+62yIBjvCyNTAFF3592Uqbw+M6TAiZYT+1W+z6OChPdWuOnPO+vS6q98VgMGkd83ppk/iu
+JUoteoMw7nCj4Fp/k7Jqjewavaclq/5vyVWEM29C+xVKerYQIPXk9n7oauHxrPVmfTcJaFX9EIE
4wyqtrDYc9NjX4t9p3pOJAdPCiKylcXZIMSZiX6N3Hi0KKbdImeQAqWEXPuVvM5Oa96lEgMVSwvO
2eLhjhWAUeK/SCymT78zsR8Pr5QWxXyvD7GfD9px/gE3HzSbWwzJwl5qssRiui76OW1aMpSzvJe8
L3jSvLqzQEkebR8J8w0bLVHGwZHilTv3cypKov1flUiABnyX2aSxJtqlq7kpcSubS6585Kwcrlnf
zEoB6Q/8x4dRAADaOZRXsUT0KDfMmyMEoY6YDGaAhZb2fsRFuNsE6XZT73pP/0/k3DVTSrqDp/4F
YVYy3daWtpBN/csWpx4E+BGfDAzWLUHI07cUNS+jTc6RY/QNoV5DgR8c91dXn56zd282FpL3n8q2
YPYi6N6Bt1/hFT4JWBo8/3uKSzn4nGhSVy1fHZVAtoUEWHGVGQOuW8LpcguZ/SgMq6HFbqNz/hCg
b5HLlwQyynNq2dK0AkhFWTFjOQjI3HuYV/ic0AxBU05DPRBEwv9s0hExmftGNgsSnzilBFU4zL1C
qpgC1pWGWra/dhfi5QjNKT/ikzcxlCbYQnLhoMZ6SM1iwEObWRz4MaTHM8ENbnHLoABBmtZWGGBF
Zu9VPow/JxBJLZfNqV8EO1aGoa+vGm9H8GoOEbgAB/oBAxhMKRbEiONxFO+VmWtREk5z4hk3kls1
ubmZoDbfR3b15yLhhW5gxz1MFoHSEpsUoyEhwnIQKKIbVm6trdxPYoBSAHBva7gU35ZDzeNSwdLe
q+QGflHT+HuELNnrR6WSS97uycYCXZnzujRVwjNpcuvG2qxlUKdHXpNEPKJc6KFaUz5eNQxT//Dg
XJj7NyTj72Abn+jMAXL9D1npeQqLdX7E8Rv2OQXTJaTyXSep7jleFRszN1bJiDNThBL7FrR3reUR
2lEKVRG24FEo7C3xAQQ8LjqalZuSakZD7MywYrjP3NdHsclAZCGQnPKyEwgX280bDg1DW/BLKXfx
qgW7W5JU8KTG69v2EWpXdIEQFoBLNnCilgralkl6wtoxdISJj6jMr4n31+zw9uWMOfR3KwREvfsk
/jY7tA2I1I1R656X7WlAErdsKIvp15TCOg93F9OLW+31pPpbebxVpW9SYvrBk/rxMJEL82ScAL8g
ttvvy6ojCGFEBrbTE3pq7BQ4jH4vIynW7UAEBMDMpS+CSBkrI5d2wNj6NhoQ29CumlFM+Q3B+KDO
8Tmh+6TvF6Q7dEiwr9pW/Q3tZFeU/anjYjJivbyJDIed8D1HH4c+Yy+o7I/HfBM/Gz6VnYEVYvW3
al6KvpzWO1JPqpSiBc3+lTO8cyx+JA25nkLWvbgq5sbfK4Qce9DJ4pj9QoWmvHet2nRce+fCi+bb
LfC7l1cG5Qfj9yKt4M/7bgpEhZasLBY2iu4jFouT4IOLoIWluFdf+wnbWGBfmVwDSKl6efT3lMq5
XGl/FKICutuStE/jGfl3vh0db+ATPxqGdgan0rOXyYj3qgAONUhTncAFcuC8wzgD8q0K6pXHvgSo
oq0ghEoWGobANpBMGQ4u4fqaD8YFyhlUfs3k5Utak/CkRY62aOSFlXSe9doyLwEbHnk8BCM0GIEe
j54zcedgyPepEKUNqOfTAYVmDchXp6NB0oGufbaKGiRgD3o2J51ETrYyFKbN2R/Ufq46ASLOf+k3
v3KNyBYXgj/9eZjmdZv5gnaTdSNl/OKroHV6JcWtVaemGb3DKfVvt7IIjpZwqgLVu57MCQo1G3BH
wFmKplXotbsr1pRRH2+L46T6o/HlobuViHHNlTGrP7jCmEjtzJpbeM7rua4DoGPjXJFNDPC1R63t
VK0VNQzpl4xI5IKtHQ5H8A3lNfmFrCsFA/8MUhOsbfN8rUKyoXS6CKOqygsDVEgCC05ld8wNPWH/
TeccHiMCLTQ1E35sZD14FTEtVzsH+5GlK+5Jz/0Gq4vUSwraRqKZFJL0LLgKncgL27rNPIYPQ6+J
tUUAoH06lKBcGnyr6bbPsowQbyPx9WJVAfhgsQoKBwZhBsOiq+PmuQJSTen80ZYEoojZEVSviK4l
qS0mD2ty1vAxauoDkjg6IjaZ8vIQlpVKsp/ON/tg6b1MO6bWt1hK3y1GfDKsiHoAjj6tVVckiO6M
tyZPos2UzwQMYDbj+8Jfv/HaVYx7sTWCwZUe7KXZsHWhhnFvGTMitaopqOaiYWJeSc+InlzJMwlZ
rY8WoR1PRhisRzRdd3GTlgmGLw+43MDfHpa0YA3hU0mFRbzFPvRx3NTJyTbWhrHYfabOC8A6QPek
hKT/yYWblV81ObzXh9C97Og8G+bLNXwDjfGm2ZslCi1+ntsfXNaCIyNut7jFrE/wCm6A12h/zLKd
OWKFQSE/d/iGKz9VJgJZIbdlGpCK7RyvkksylA1tgMmzIB9k7yQUrEAwLsuSR5KXK3gRr1vLvbxP
U8FtG8t5sYgEdRx915x4RhivZ9fNzsHuSSOgdPcNUSCVjD7XLJoXA2ZDpANt3GwpSAg5tZJYx3Vk
w3THoquUTp4DPTEjkQ1/VCsP77NzD3lKC/QRMWIAhyaFbmJwcSf1NGoAE816tuWXf1RB3IuUBXfD
qgIcwOYiYm8OItc7UhtEXVOkhOVXYFepfPZMmNw2a7aScOsc3EMiP1rDldaRWHC6mGhGCEJBjD+d
cVwmnptVggazYRlIN956Ct8xMmI5vlhORyEhK76fcKhcHmB0AKSK3kMO0zujl5jj5lZqFx8sVXQu
fon+lFyFh3V9ORj05ZHvfvmtCfTvzSs31KUACPGtsOjVwpA7ZVIacJxuhb6/vjGPz/Zy9X+VUcLj
RANNggtbjK7VMp7AdJhmfKoGM3wd9W6N87d1miSxTPrhb04GXlEseHMrTuhELYzrCiFmR8zZ60D+
M1WKd6ALeTO5amN6ZPnCOGqGyN25jOH+lXHoAo8kT14mDbkpZkHwaljvEQC9xq63g7AQJv6MxDtC
xqZ/s3EzlzUgaRo0jZWcksJK3sy5ackrXmiRebgRzOSqhu6at/EFNW6p2MGX5UCCQfnxMXsG4rz3
PfHpnn8TTJmthnbUP1HfL/FmjQ92Wa97Ln/UJmmr4KKGFtXe1ARjTDyfibZlbH5Bl9CKQ+iuxHha
kU4hCHmGwtj1O7KzAt33oFrCpwlquVuVYlPd55KyprQGDZh3zNYbMA2B/FYOb1pymz/cHxpqOf6H
htuJgQ6k0vSPMT1N2KWF6Q32f/bWDG/TXVZvuRVDaMp0+EtP7AoT3lJb7CePbCIHMFpoLz2ZLIov
jKOLXNc2uk+rcXcoN2/OlkZsCnm6dWNplR42z8gNzboevZbOFKTGGlF/y+DREt/0h6osSA/KP4mT
IZFCtqGdC3EGrZsBXTY+Zu9Msydrr9Rlz8NONN2yVNiwUuYRu4rj7CvQKJsdf8hwZAWBCiWLiJGH
a4ZZTlLVZ4VgxC9cHybwcYKzbbs4XfAuVfQXXwNGgLeScxFdC12WK/P8heQafSc+CZhNUS5PG/1W
uQOdAb/NsgTSXcbKPMA/B7lzJ07gYfuKYmnLETQM0fb3e2E4knml3xfcRBbpbGGoviUiWMqwCDaQ
woGPVSSuOe5dpI3ep1A1iRWy4xiCNtCKDXfUV60lvhvBPX2B8s/d8byMfHAmlV7SbWrpKLBobKNV
vVZvTlBztRW0e44LznI1LcuIFjekODpm/9ymIaU1NWnET4KQY1j/k8aJaJCZDY8vsvb4hdJiku8q
25hg4NAPz0EV1QC/Dxh9LLD4c8oNZmBnJv4VpZesALZvgirY4BnjQqMEbQ/GgevRaviZJFGHhzf5
ft0QNxFb+UD9t5q6nqOixiCl9kA4VtyB1wbAYVNI9caHufN9whZa3LVOcxBy1E+8WRHPrxmONOxK
djwPEfcXXG2/l3GFr+oigYBBlqwUzAquJ86cudl9NY7b+VVYC534azcs8JXQg8abnPUxzCrCaboH
nsZBpoPx835wUd3YafcExtwK5msIXc3bWbISJodbFACoxodvpUtIJ5SpLOR0+X1vXQda/xcdJXw8
UXnmNkNGm4/lk0F6cDOoPvGeKSnrKU1k8BQMfMNFoBD613Z7pwlTIPM42b015DHxDwLAFy2/0gh+
whfQBE5p9EOsHWfIxdMaLx/nsSpGLWtZk8Xk5CH0s32cHHtTakxii6hqkDyvRIc2tpT7bNHyHNp0
y0qzN3659KxFjjaEsAnQbPJ7csx2mpwLA06+7Bc0xpYzCBc52fhxSdLMsVAYGHxNyJZ8XgEI0SxS
IFmrqi6+mJFdNweQk001A1Ap7lWqSz2646Nh3dOEeLlvtyh5FEi3BuKMD4tVwuB726j9wTR3U25S
7MxNTRUihug9uYMuPMrKN6cr3jgyRmA+JQ8191B//B6kXkyqUG5pvADhjqqebgIwCWZ46ELft9B9
78dnXzUzBv9/R5znmQj12Rh0MoBeYCougNMWl6ymE4tFITghrY70jZ8/pEJx6Z+9NPA2aA2ldmz2
zv1W5pkQyajHzPV6HfRrGyW+Hs+re1MVmOGqdLxVJeuYs3Jlh/JJJdMFTb6ZCF+i+9mARAEBhw20
1RiMUMkrTJHvVUrr2gox6rBkBtuReocb11WiKIe0sXDLsi/Yxzy9G9SnNAl041rMJSX33ZV/QTnf
aQeT4+t6KyOl2n8yqV+mljQ+owVU6Fz33ZF+iz3rNyFRSFneejlAancB179cHLGtPgLegFvHvGkT
V1JsEi30agdSW2Ay347Yd+8R6pmNMiEvpPBTvMcJ6o82ZH7g0yXfq7nUGO2bsiEMalJWQj+pU0bl
Cm5w67TmdtHGwNtiVrKhTIQyq2tiZ+nmn2CmRNjnz0xH2OinrubuKFAKg+XTssWYk+B0Qqybosos
Dt+MGYvqgyjR6XifJwi7FZff/u2xahlpgxlCfJDIfLPamOPll/Pe04oVXgdnCfFCYLX2VU25pD7s
Ii525o6I74P88AVCQ3Kese6pPHAkNCUfp+9s9YWIeOSoTnY5hpC8T0kyYJbXdQDxt39Bn0zL3sDd
x9AcIbMNlbHz82jbL88VazDPMR+6F3jQWDQq51oTqM7O8O24wz0B1sSpeb4m1k/z8FHEzBvc0ltO
Rl+62MahIqlAj+b08xyFYckyas0Czf5BXotdTUgjUopGtkokC5TUuCeRosmWR5YYLJyKCqwlsA/g
NUlw7II9kNnjPPFCMqW24ljBiQd0PpTcpHf3r9d2SG1E/GZhZnnvg8baWGs45upDUF0EjC1DJ/LU
3asbSAETtuMwZfoba7GdKCt54YYp3vk5ZyyWhJARY8NYrpDmLaiMyJy13F1adDkKIao7AXH/Ny8m
JyXQDBdlwJFd5UpokaIaaa/7xz5M9K4ZDYlF0EcsRMx+4TFk8WEXqleIhXT1KBmeXKbY+2jotrIL
bApAwmfSjoYGaKF22WVD38/ST5cIUQpIvhW2rngO6PhItA8zSoQUF9BXkkRLnKqs4aOe8BFkvkQt
K2MMkpuv3T+4mrykr4S0Gmg3U+dcLHisfsm21vI6kJu9lJEkcupfM8OWbx3tVCbNElDclKghELAO
KjqiJtQYuSGht4MKK2sc+8uoMCKQAan4oGN4W0TRt3g92EGI0YZnrh4qXXWHruu1kbmsyAFRjm8i
arhh2h10/L0ts42F6xgGyjLudVfa5vOFBzutuzEzyxZ7kcB/vFQzdSZzW8mxr/YgokXclgb4d3ce
0BeOgq85AFHpCI1gzuIPHd379K6Wz/6zVJAsKLZFf3XHB6TQH/byH+IOMP4y1nr7O4DjwXQNze1A
InxHu6aukP4tFoMk5GwwkWcQj8y7k9MlHV0RkRhbWJTyeHBu/lkeApZYBYhRts4Ue1SlCaV2bB4J
ZEJpqnTR/v1Ce0oIV+0kkEuvJj/mvmGxEOvWw0aDDt/BKfSrYCdEqVo03DPmrJvi+Q0gMbgiAOwF
iiEcY9cvA3Hyp2vO0JDBBy5FGM2A4dwUBPSKty93OXBUWg4wwiRs4a2gVmAjR1eOKv3DOiz6urmp
8hHHVwJ7Da9yK7ea9onb5jWbzkHX2f2lrAcUCL8UFY7vMvObRvAp1VM1sDCtoA7QtCeZvPUxn/m3
+LOXGT1bbNTbPP8LlUPu4FIMkuhr0lWHecmfdki8nZUaKgoGcNne6X/zWlQnrj2cc6WWzjNqMRSL
SqQe0V5kXM3rJNQTlQsy/4KQGe7fusTjzTCMk5IdAY43l0fr6a9msrPP44VPTblrNwf7GEH0aBZn
EpbFuIQv6+zJ+qKoa5B2dKJBzwyHkVYBnvWFPQJEWZIg31OEc3JKq9Q+0738gBKjtzU8GMHmytx3
0WhoF2i+ohhLbD76PJNDXWT3ck6R8etBSvM1cmoRUytcQnQFwGW+umQB/L51zEr+7srPi8GY82gg
BuWxqcNFXQwZOTNK4AW1hM11pWGGA64yAsdx/hRWg35oy66wmmzx6Ufblelgzw9ZAvfKN/z2u9ZV
TteijtrEJ4DMzD2yrnQjqS6pp2FaN2l3TXarUSNEom9hPUvRIsJaMS6PzltAn35hjuLZ8wXiVryw
n+rW+3azQVRs7ovdiFlejgpHvQxmY2k9vd+tU6bKZXSkdD5mqm5hFXXtmHW/qgGkkLAc0IixQxJ2
1+4kld3W2d7Vr7bevznmQ0z/4muw27178hwF8PJr+x1xD0rcdx/X2Jgy/5Z5dOno2VCR8oksImhh
oZG4ZkWfUZ+iT87IWtXWV9zxBP7DqGIp3Sv/sDjLAHZYs0e3hd0o+76HqOfF4+Shoe53tGXdujWz
weLVKqjiU1BLkSj7vA/vjZSoGqDAgQBbVzCdpLRHvcncQEbBhix7pw8Y1w+GfNozed6FfnXWqiXX
9Y70LXLYypyyCL/cl2KkpDq0Q+Z2NhERSSnrorXFT+kRSUHZoFzDvWV/pYV2vjXWrB56/upyXoKj
tV9un8CBFsFoUrA3oITTNLMvVjeJ+FQF4smnAdtGfSE4THu4ubt3FPJQOOT+l6WigRAuR5eUVCuc
AYWB9OxlG+LpjVOYhI548i8B1rdgry0Ncr4oorzq0Kl8OcmIbr/bqt1KAvNv0ung7Q4n3FOyTIhV
vPKSHNszdeD1ZRPUMnFqgiUvprzNdyVMz3+eyhSmDlklp/WSf2bI/jGOERENqe3P2ngYRzCt55Bn
/dkrwW2wE1Iw6u1dUrZFpmaNH6YQlZrJ9Gg5UWHR/q0s3ne1gXy48BSK5PJ/bYLpjvZSiQtUVeZH
6m3jtaWR69Syba0lB3/zroxIjGQ6/oVXuN/dtDHkeHELA4QH2av1n1DE0vVFTENRJm1LIGAYaZgA
ZpLGvbgNEJtivagVDrmCVYf2rpK0wFWs5/7XVzJGK6AhL0wSek6wmbY8upY3tHlEmTCl2QE7y2ca
yRc+vVcjDfIwTFBO47//GlXLVKntANB0+OhTgZFd46KiOAgIUqTQcXH1aSXU/PdwmQX6NRPl3eqE
cdHV6/mLV7pN09Y0F5tNYgqxkp1EPgo9sWk00h8cRoDMqJwlFv0Y9LSc6gnjmXNTaDAARpx7TqGL
u7DvJwlyhkRJ2bnbyzGrSmZS1qHt9KqT4H2bEAGoXT/jY6UHCTzxh32x5AMj1VwXGwbEA/xOSIWx
gXJkqHfAA3X0eQaFhK3QbHLIDKnKG5mnYsK01HvZKb0UIc+3moICVFBG4NVvRDQ+S0ABZ+nY+lR4
jTsSaTe9ynuezjkZJi7deliFHMIH/ApVhZH3cUXuYDC0kn9tm0IA2PUmUJZwWjX6fYeyLYUrmW45
73G1bOhpsMLPI4osiG0JkPve+k0lJLFN9Vwz33OBvgu42DLwBQgDOt+2gTiaRcYwE/Dr6OPhEKve
2dQrGwVO21aXb5AYgpIJGHXeUktEKnmwvqAwoQ7+Rl3oF5fumS68p0okEMTk3MpNCm1Z45abOTlb
oeQ0z4DN3Werw1GdNvj327KvIhb4+1R1Zw84iqKEeve0cP1Hw2lM360qAA7kWz9rh5IKYp+V+ajQ
jUbNo2IKRH1QTKvTIXttAPd3rjsDbYvkTkLl5LzeFDsBufLPZLvQJuOICO2R7XrMGsFariXZIDrD
k8CEFm5Yd4+sryTwE9ldM+aT2dsVJpIIY1PjTsTmImsh4JdFk+ZHayvB8Kl9GN93M/UPGaGtFotn
UbutYB4pTFgNnv5rTmrNBTkdvYcX08wB0PQIfII7TjlWlQlOSVgqfq1LOMe0oISY0X954pQe/Sor
H3GKuX1HQIoVjwGlxmBbispIUmSfaIoNqbpWtw6nKb0qzG09fNp092l0llEGhDurHp5aobWUYZ3J
wUZbf0Cl7zh5I/vTQZi77HP6PlbINvBwhPyNSfxskr+5/ddpzfl0JgBRuXS5LI8Y7nDsI0NRWnmj
b+/ZMJbwJ/R/MWdgV+c2H6WDUe7K+2WXob6JLUbgzDgunJ/6L51lib4KlL/csKrgNWNqiKDXVjFt
Z08IqKbCyd3LS1PEnRgmQQSkDiaBTbZCAcV/ZZCf6yILGnB3neJwLApNKKBHusfXClYNQOR9JxIb
cUPHSnIy+X1XwG30eQ4rfTUknKDH0VkpyVcAb0MprHeTewlkLciUux79082HB7RCmMLmk4mFmzn8
gja+TSJPoM/UvYB/78SxAvo92fjLTRIM9bf0dQa/CF7LPRSXNc6lceJCEfMq0oQkddg1oNWKBCnh
Gt+NpRhfA5ctD/tF4GxL66KvMmPBMl0OfcnPzxqoDfSFrsAD2BjYbTutyeqLhVJQaXBLPxx50a/S
UZ07HsFBB4NntN5y3GBxaVe6yvLeJHvZDB/PCA7nn7Ofwa43NFZuz851awDR0RRUDN6+QePaGNkj
klQUzm57YUspzdtA8xWkIlEmZZIvt3+5f21Z8F7yN5LS0rspEHC0xal6CTI6aa0Q1riLNlPqvxRS
bEAgpX1+SXyD2zVCoG48ysxdV0CM08pPmj1gf5YGgHxt/dJZvwDWGjQ6JSrycivzpjeXU43dsdB3
3qAOFqpZiycSxpIbgQ6UDJ/PIIVKvktuWLza5gsAGWOzaRmrf9CrEazM7NnfMh+uhuAHagOEtHSb
iBnwgffsAy8T9d0m6GU5dxygoXI+VQPtHftW/Jerujz/WNl7KNasjDNFnDY3N3PrY0WLr90mkd0K
Us2zrd0FW+FKjDLlVUxDApvuuWyUawY+f7EJ9yAJ3T27DkJiJ7qB3Ehvnsw7rW9kgufye91gC68C
OTBLiuzqMLzHwwnhnPTgXyfI9Nh4DZcl03B7KR+ykrQ6+WBMJ3xCEg9xABDJGM4fwzP7B37FSi+l
mF1VtrXz6tkpxsA8N/tg9yv6B99pi585cyubdxHGvpoGWTcCWewNzx6n+5DTg9t9/8IAWaWcQAUA
tI4ZV1GiFBfcZZT5IM3W8171GzIFQsekAZGIbZ7+DvRJ7QKTU0T2UIVFGkhl9gmKzGetB4mLdLLT
VDfpgK8a8QbLcMJvas8Mu0PlUryVwUjXIdmZI8JZmtBekkDMGT9GuP6sScbW6iznpLP4U232PC5B
+415IBmifIooQVQoDQHIJQqf+sZ1lhj7UC7dhbJHkvqpboMuaeP65vymsZG7q/ZdNYczgoiWoJ78
uud/gYcwyeVf2NPIjxxLRnXivl8aZY6Nh29H33H1npI6BE5zdQzUVs8xUMX5boYj3nvQw9KUJ1L3
YHpz74x1OVv8U+LPEkOv3C772gvj3AJBlCN7ZN5qVmiL2cafcjGuu4VqRlG8aGoPMH7g2lUlHFHZ
KraKdi4ppQqnYuSPdUNAYrV15mg16G2U/PdcsUCyW0PqkAn/4owWhTxfo8WAgHO8kpotkA/mzSyu
jJfMeRqv5xVGOt+07J9xAldOb4GqVoB32dbqyNJG/4Re5EXtLVxdH8v4/9KOwiG5Toanvf3N6VSK
t4twfCWi3C+Oa6pqSrA6O9dqlBtmfEE+FtBRpmpzzRAxRV7lFGySZuAY0X8SoROx/60lnLrQ2UvN
UBxkNOBCdCeoobfjJhJmV/RPJ9oaxZNNlUXY8Z/PTfZ8UnKcnbRP49lCtYvekh7To0hpo9o0oHMY
e3lPdmgaaBvG8jegz3Pe2sZwwFl/8VJGaDfsO/Y8UMmaVJUfJj+B0UTph5s4C4++x2oDv75FBS3I
9iZt/eQYEJvg6Pc2RgHhKypPxyNxKKbqyTIjkrcC3y+zB8Tqo2I5/M4PPSxk4E0nELg0i1dfGv8N
Py31HwEPX572Gt4oZ6aV2gY4i0FsT1i0j+ypPkR8W8KY634STfbe16q3sDt0zvmbv965c7sb68t1
0LiRuXFnkUe8CiKnyedblgQg++m3JcipuFySOqDGLanD/qOQHPscWG/tuR+vZLyB4hSXSF0kFyzK
tMynq2OIjC00I/bYCW3YyCLpmXcCy+448t8F5BisVrsa1phnwhugRm9ltixvT+mAKLuK1n80gWv4
qH99ewO1AveDOSYzmmhT2FhyWykBQtq5a5LTCS28KHGBzxmfZp8v7cmqIyN2Hd1nY5dESu7xQ1cU
37l/LEjSCsLdutvxnZ7YFYWl1TiR43zU72iNTTeYUXfb8uSFLuaeSeIlLttQX4/HHD0FowNuCvoZ
C59L5AdXX7OG3aRTktmtv76yd+h1Dj2P8zQ0xviCv5VGPO69PEZfckPCKgbEwTqqLFI1+AVLmhrT
CAjbJq4m+StURstPagbxrmELr7GOe/5KSx6JtBVh2JvlprocQILdq4QSSRFP64mhmb9WoEnVYVOq
eUxRcmNKdH7soJspKDx+JMZ5r/1mNT0/sBgtbR/EyGzFeciq5qBeLAIJOcyebNZmRpcLD5D2wgps
IGNexdTolOtR5CgRdCfaZ0hpiKqzSuDNIxjn6WRdB+hioHnM3WEQSNSFy3RnaMktOipjAW36wVzi
a0D1suOB+qSIZirPTNNy5XyDv9Wbd3oxRqN8aVRLUP3hl0aUahVDrTkH3E7EbqHUZ0JRUEQhlDTe
YY6WdxgytVsH2xMtQBS7Dt6EolN0Ti9DWkWovsJVtra9hxgPFBOdAnqVSF4g/w3Ko/SPoLrjEX3u
hBoo6dLWdMkXWUm1ssQEeOm81Ob3YSsfueQz6xkomEHAEyjV6nLKCVTv23rpTyEFS6mpqhuL2GHv
lTR2bKRcGXW+2rD9n+pz7vvlFcXFep3xKcksrsQpIjNlUNuiy9GxPDs1CyZGImZeaWbhbV70Z5xr
vUFAbuFXbeRnjap7lE0qxby9mygWthrPNKlBzm3IRnBoCrSQNZ9lTC2LAjUbPcdgRu4XbHOwARb7
sPZPwdiQ4VNHzzWv9Ao9IppsG2OXDVSzAzCOhhl2aIiIlVC6VkhhqBmJMi2J7RTS44ZdM6fPQkVz
alnLKeXkLRMylBx5bxwyUqhh/JBzqUc4mFCtDsfuSmanvDjZ+wsQtq2vX89Mr2tOCfbHGkoA9c33
pB0EEiCr+L3ttvQBmxzeJtrnQFa/cSZGbpyyK75ppsPGuL0tkE900dAC3cGQ9D4auAMdanW5OsdU
FFAosRCkH3EeBTIbpt13vpX9lD+fy7apwp74xOgPatYoVsjvWaKdVxlks2/SZwM3lDr3ttbqTBKY
VMt3CBW6+Nx4CgrM4vj/m6OpDGarDiERxIcfkqkqwwszwthaifQsImDmpLKdVuMyNuoYXDpeHfiM
Wf0JAZ6//SGBADzUodo6HNu9bmhLVmsRHQEaW1l/MhDbtYBX4Qgukwkz3zSDy8gsNmSvNw15g8Fw
SJ7py+4+kh9xrzPAFZ4pf0dO8wnXTk6wOkW90alfDaaQhEsNnzjo2IOVOtYQxJ8ClErusKk5ghqv
qbeuXZBnjsXb3A2QzyB8Wc+04oir9QcUNdj4asem4dGL/fzjKzO/VYtJ2ynuRVQigHVaZyQs3Ds1
MW7vur3LY6NCIpTdXSEplkw4OuYvHCpeyRMnm3lPC2/ik3ikSOmcsCkeV5M+v4t+fwTA3kxqeLta
HzTAAQvrk7A4gFWluJx8Gr79sGTopIjXBkswOknh7mYVLUtZX3xhMRh4LP2CIdNHrCUVMFjoy084
TaZ5X99t0tWH1dYNH+lSMS4VgGz0RykCRpI53Wr1TrNOKH7BQdPtBy4ce3lnfqm2DqQV6xu/s1d1
ONO5XjoFX3ijpm1LinKONkU4FCkhVeC1i87y0lmlPbsCaszi6TwJnTda8ZPis/Q7XWCKEiN/5TPl
o0g3fsKEkS+fizoQLwEoEHiqYqC/YDRyZU6WEdnaZCroXbP87XlGJd9V3rlKawEoFupDlo+Yu9It
1Ve+ro6UcJSSWU2AhnxE+FjwZEQ3wMyWGP6vI57KVRiagWZc1h4fj9NxLbMmodwtmESOn+6ROZ+/
/t+vzmD5fXXGG22ywvIAvMyh49wZTaPnYKxNmt+8AVPAHxQQlmUpekSJupwCpQaqCaXBADvZlq6a
GlJrNy65JNTjsQY66t5R7jv+vQjdv5GbAYMo0H2RXDeO+eXlfvcuV/iUBfgrDRw4ozcosSykq1eQ
vqzkfBr4Q78Y71jB007m8Pohf1VZcOpjQN+86PlXXro5hh7RweX5cAyRhG4+EDADxCgie6hSyro8
EE8LvM1yMZuLD4DLI9ojij2KlwzafYks/Q27ian7Qo2mQNOkD32kGeXfOLJqTOaL9Hma5FSlWsTt
LGFL/J11BugIxdX57n/pWV7GzHLbyoNWruNk//vWDG16Wc/ydG6xYYGUM+2jfkq1bSnG8kKlZXSg
+DXPpxGqAol6FzkqsCekiHvBhRw9kRujALQxgEddEpZQrb8aKer5m60HI+5S7CLIXtbuaYlrp3h3
pxq7LGEsORWIsJ4FvDQBn1GpmtdmBjRXbhXvAcHC4wcSnxYWgxYnUmWgtkC/4+QxsIVlDPBe6Ikq
GWAKzMdoOQOV9xX/UrDHu8G5cdfcizgS7Ll/WIURpYaSlto8hSenBXe1PDvkJwLivFcrdhRxymkb
PNtwep7QMiFHwdJXlt4eMW/pB7quVevYQy/CCpzHFw6arA8yqPOHnHIa+UDZUwLaTeQ51z4S13rw
I4Umj8oEnJJVoab814NE6vgfh6nBCNAnLzHQSNkeL5+YV75l6J5Y0ntre0I+0DcS/luUmmBDJgDS
tSJ/yYmIrGqS1ogHop66CvCubAfrlazeONr0XPcbXJyKLz40yhTvsB5DyeKYB4f3mUoEsh7644O+
DbINASc33e4j+0ERdlT8u45fjDZc8pcRLYFcMzdo9MdImYEmcnoLe43X68TAiolXoNbWBf83Uyo7
Ec4m7nDxd4tNaecp7nrmuy5sIr4BoWxGUw7I6xPAOuxk6LFuF58t7YHXASVmu+HK3B7myEjV29LB
V6erfsNGlEEuUjARogrXG9SGf4rDkhwHQiTM0VBMyBgCWQFo32awInbT6LQWnz+A9S2khWLvSCeF
yn292ZQooZiz9toXzST8GN+37fxlKdcfsjFKyYo6/PSoiI+0J0vamEOQyjBWnJdrKWMuDsb7ppvO
uSQiyDN2fBCsDOWR0ky3ZVx+7pCaBJmyq005Y4eNts1UGq1q1hqW01O4u41zL4hloBU2ch/OOxbB
6IPQHHqvotVvpj4BVf03V9U6lOyW1yHUTEwa64re21n407m+vZBpXRdEAbUmysefoLJfd/NO6KbA
CooCLyuqxFzyKa/bJ5eJ8QAhUp/VIcbPDQ0+xPbcXw801Y+m/KS5yVw7lkIBmq6P6fhMOtVmr+Q0
RvVVkfjdfya8hUwJ3l4qABIOO1+F/RmfGVZVxELC24BWY+sg14H6qSBnzh7zx6Ud0tb97pHHXI4c
qtD6dFquEcGbc5/Rjr0PZBmOy5/VmruNXYcaxlirjNKt76IIYLrtJ0mkNCuDoc5x3yhq7elP5Opp
DTOcG90SwcAi2w5RFHNi8187Ly2TOB1JQiw5BgrYnqNno5Ccvgmud6sygweyVPJRoUIaaVWuaLha
0szmAvjIYJE18z1NuFvhzs3EUgEj8oGOIlW3ra6lgtWv7FlFOdSm47P6Mvi4Ejc76yC27kdnEL1U
4OLVTqetRIuoj1HuDvSGn71EJQPktvCsIdPTO0ZwRcMJ2BEvgj9qDVs74xhFmH3E2aeyCesiLHwU
hoaGv2cn/m1AULXrTNkyYvEdWPdOrbZXkdnuMEVHSfT8qAN8EQtckLFYc/fNw4LNks+YF+Y3M4Jw
fzb8/v0VOgQ6g0uw4l6GhSYnBa+XJD3Y89B6lxpBftMYmGsmBeEDo3AXBWfAc0J2w5GtH9duGHAu
rs1oqWK1lbHXkg9PBzpevHo65xLjMHr4vyu58QT/Kop4PiGIDlkMZpzms0Cz2hhSfPfF8ZOS39nm
hjiGzd/pAffmOUq6gxD9DBEy7cmDfhp49SuF0JRC5xziN4wttAvjn0O3Qg3RaAdrnRh0hmlGsp5f
2IfW7vQnHEoHPdp9qxCQNeo4cZ1fHE2YS4SZTSrCqL8CrycR0T25FxP5DavlmaYGlp6qZtiDFsrA
UiXPGrjJNkMJlyTtE1ztg11KIo5CE/opsEO8M7P4TnTc3rJ3JngzCZCQM1N9FdvmLeKC88rj9X7W
zCjuXh+3ME9ha0A9V4XwGc36BbS0uzfPcoJqt+I/NarXVCSSVVzVtoFVqNiNKgt2SQCvWGD4mRzW
CTYzMOLCYoPgggEBFnYDOdaQ6tq4UAr1mXLdQzwOKuEbutFk02CyNXyZ2U9uDKbk+3camAUgsbco
CGOVSnM5u0rwkBjup6SEhphW+tlTXKpTaf0Vp9kMK4uwqmDex91txlHBEV2yJWUAnvKWHVurv5VX
CQi3gWbIuKFo6AwBKWr/m64o1+GCV0Ew5jOAVV9Ak5nfrxGs4hvr6ZGfPcWk+kQUSkM4CmIB0IpI
ofoU1orLTuJy4bOh2P95gfFoHrg8LK+fGywTYUjEXTWQwAiTOlIo91m2igwl4DvSb1BRs0wbRGxi
UWU+voUYyuN1cDxJfxWzqStjg9jPBQ1f0wodit1Q0VoEm74Sx2SotDrQN4lKepga9uzlIpiPIImD
AS4/x/Wk82PwAgLMdH7pFUoNV1bkJyI9KgO5IP5EsBfoYmlvIAEON1QvBNOvqsEdKGgUyMH3A40r
bKobarx/Xoj2wb8cBK6EWmxawRmna/JefVreE8+mA6K6Vzqx9eBGPZXW+geDatEmc27WocHB1Gfm
/9A3hZyQakvBkQT4nkohycZ7d8dZx/fEo99tdvJy5KnJMv2p+YIkeotcPondz7GZ0vw+Y4qBMZE6
VI4HDh13C0c9lCaC1exECkQ+d8FSVpW1EtFVBbym3K3/KM/ec8ZAyQxMMroTQmsDBaaOvsKsO6cb
c/vL272TrjhmUNf6D6mDPgwRRlVu+SP4Qyhj2XZ6ug8GEd1jZzXt8hFPWsa0JeFB0lU02dqptH2k
vLoyQkzHfzojRN9jRxiaKVsKtXutI/f+z4hsfOlnaXYfk+/bqI7iSNB/4QnNfP/um7gdtbt708nD
5kXdKvBdJuoWP8O8Vm9PwV2822UsPD1Jbvp2Uq22ba1dnVDFMFomEbBCLKOy5B7XeR95ssASL+td
lJFjl/2VeZcyRgVuMPAK371YzsY/FgAUtUcEoROZJg7m2tKWnXHSV1sKINQhMhqS2eG1Cs3BTZXA
eJ4XvQC4Ah5RW5MlRS1nSNzaLrvZCkx/xhvbQA7u2aoUzJtjySAGa/b9stQ0UqjJekhv04oXOYPd
wa/wAyNrC8qqddMTPV4c7gS8SYKlCTCnmoD+cZJz61oi5mo4ASjt3xhhE7jOOMJt357yL3hv/yZO
iaeZ0qrRp8qITBM+qEYOPjZNkdzZvzvMArVwP8AKD2NVcpJf+MRKeTunx1TDslXPRXStvMH1fsEn
SB1/YEVBqhxetidaL4ZAFiIcr1wvdVlvfSVNzxuK0vQ+DkUQvZ85o3ZM93tPXl40zgd1T5vb+5/Q
p7Uuun49V59iowWnv+XoRqQ4mLlL4a+SDky62mpYii0YRh7ErE29GrZ/lBmGe1WtCm5XIB57/rG1
0b0zm7TV/dS5m/mFAbvYqqG+feMllZekbyQmLdoBuaxBouc78xMrONeJ5nUdnXKd8PglQGq0gcs/
+e2i39Hunu7jHQ2hq2c89V/fjxopRsu2V3Zt4ADTAl0Bg3tnCOp/3alVGMFx6KlPpgm3rUklN0NQ
8AuMIgkye4+Df7sCVEcnkS4WUDc4uXNBj8jD+xDFsPuS91mzga2wxHWcWZ30+lSu46lt4Tj+kuZd
HFCz9pfrd58RyWW4KrUaiM0tY42Mds2Mc9ZHJdVHt11FUoK8Ez1BMrDL/ck78JrLKGE2Ft/a0W1C
YzXxtd2I3Ors5g6sB7UAsFKXrACu9CkpiVFuK+o5xqk0R5ZWfrcess0l6z/3VtSNJhSHbEOaUq6i
lVJmqohlavvdxNS752+/jhOPobhuo/WyqwkK9znjNIFAFPnQubx3Xi3EHIOoxo90Sl/mgWhyvdsn
9oLi5eqvvvz0T8mc4llYkYP0ux/LECatnwYw4MP6IZlT901+VCdhzls1zUJp7zGY67t/AoS71/g/
ng3iJfm/RZ7YmUz85KSSYWE3GLc8MARN+FGgSAOW5reY7hZyIdFwQOTu3hQ9o/Na5upI6KG3nWze
27nzh18RHKkSeie8g6J4fHwpFPdKYgbNR1zMUCmmky7uni3OatdfAB4QkF4+mYKCOoloHVjAet9c
nBatU0QoffUitm2OJCNKzS564nbn7m3WfX5+iJK4dHXCUEPL8LLy7cURd54ae0aafYSh8Eb9yK9B
c6OxZEEX6O/04iWvVAeFinNk6ob/dmQMQ6Oshhij6XW+Orqael7b/iQYMSyEEaawasMIiRXJI2J/
fkJ1Kqin+ylWlKSKZoOYLXyliY3s6Gctcw2II5lVidKQg079lZdMArfwItYaa1NcpVYc/9U65rGq
9+gJAxIAU2HtdA8x/Gm84gqb8AvYvfKmUHXsaJ/EkrPAweNmfREqimgZKeO4Sy81aFWPKQYd5c4g
Yf5i72w1caUR+DCc1aEba7CJ5jmCepGW8H2wzd2pvIO2F/TRzmYYFF9uhtGLAmmrocq+MMzlJnub
LlRs1g0JwXzUbZGIFu511/G8OSvAjufhzJx4KqJpafD3UQ3GR6uWFw19bDa58cYG5LyYhU6zs4e9
kc3wa7nWGtETeD6Jl8Ly38RYPeSYYJa2kSU9S/j2ucUOPqBfxGyEOmNqWQWP2xI/WukcYEp1vmdX
06e96rhRSUFL7XsFA4TLbppWzB3sbiNi8HdMufOxIGbXUFMPpBKYWysriCIf6VaDSPLojd5tvcow
bwwnXiz3ncBuX23xI02ghtoIhGUq4TvMI+W1yr7RvuFrdtemC93mt+u71PhksGf1NFmIlXBz3z+t
kFHiX+cXhaQfa5IAZsArZN/6P+svr1OLTESsnmQDdwf1NTy1VijbRosLtQNvS2Sm7eF3YmsUqHjQ
teoQNcICiFiScpIVkslh5FtOMWmGkEUjgDelQ/+jOhNaRoP+euRhNxCwmzMuHxmdlfHpss0vTyIp
NhJ42DotasbGzSTjQNUBHqjBSVW/1EQppHaEpha3/6N8EF9WwgsyPSSD2HBJoYxbHZlw3TaVTvn+
duowJaHn51elVVCCseRiXCf+emSd8MNcRvC5oqz5PSr5ZtTofitE1kUo5ANS6YSmg9k3zpU/AuwO
eulGY0XjRC7JWKZR8ctP9+cveeMqS/92nNZjilSiPfwJ6XL1pWQflLq92ErimyGGWXOOX88RsMhU
XVvJsWxm4TnDPz8JXU7BOwZRULtcyZ1HG7KrdbVnsbX+JdUZpyYSJZELDoK2LWq+3bpboaHUVXie
eCLNBiME/gjqupVSpQPXiOxadeDycj2ySjIeswW4S4JNwrYXPRgX4KUbQTBa3w2UcCyPvKZnLNrc
ReLLvmDJ5g2ZbIBPUQ2ZzbTA6D0UvwxG3opZtmILFfCVFXkKMGBjTJxHwfxUbD/jrtd49GfxIGRc
iBU7/T4JuRbfLstn+2l67xTJ+CBRTGZWvF4IzqLQNbJtat9N1vUC8X6xnviUz3tz4nDEY1KZ/MDU
lmtVf8Bihnz81FnBi+hoKGvP8Qn9NG9kBv7i5xfuI1jqFyifb89VHNXDBq6MahBsJsPltDREH9bS
duJL+G3Thk1zffiH0nB8cWw6D85CIav9Lc0htnC2YyNVPym47Emn5LAfkNXOA1gGhrCU1dj9v2aZ
nizuz4qUaxwoKyGxzesYy/OiCdcKIyun2z6KRrlYLOfyVWQ7yn61T9l4fP+Xck6S2ELvoLuz4gEv
i4pEmdEn7rtuTATi2Eu5qqHLyOCOiLA2ikDjW0GgFtREksAkkzodKrgP4TQCiyPiKW5NEZ23Ajdb
jmhSLKleA76Hf172rf7VYOWUn7LgQJw0E0U7r8dyqATECDK7UY5wBg48Ffz5WRa4YTX/BJVjgn4y
oYctSDbVlJsJlHmuNxHqec7pCDYzHDdJSycJVxsnWvzzMm8jokjMdpsJiwwuiyGOxpnVGJpEe1G0
pJyci5t5Ukywbf88wYGyvO33mKHGnrsEhZ0da/M68tTH+7JWK5+bo5Oq1Cmi4UyFMhAmfJhO5sg4
IfOJ3Oru8yX5ycc719skKs3o3lW6p12rIOA6+Vh22aBiEBkOIzoe26fQqi8mxs2STVGWaWQCjtnj
t0+EHDdfCeEjWgwudEAs/EeECGwIDlpYZNYEn5teJLiIkp5EQd5r1qJKiEfUZctTXEHqxhasUQeq
+zYxIqdQLPbjO3PvsJxK8E/TYDIj3QqlltSEzV+Fy0T3ZmhwOE4kcZbJTgTitRDFm7I9+aDJyvd5
PVkPKkkjq3IqnAdZS7LOrZQ3c1Us4DEXXlMUtp2LQjQUwrCGpaOpRx7GOYBxxaYQd2WO0JacRymk
XpkKnzyOwKX+GZg4kBaihk5mih5EGDvYWXjL88HGMYeyD872Ux/+i4qAiHin2fPig59gwiZaLU1e
pcGI9xpHHy+Y3qie/NAhbmbhIVfVH9YVP1YjFCMAesjmQ/3S7qB+lkJ8tpeqCN/CmlsRL9mHcTh4
q+j5L1R670fUuGjzqKIMz0TDtYZDVagYHXCDSkqViKFDQmixCls4ukzeCGjcw/0TncLAfSRfJGfV
epYGa43jF3VDX+jDdmvaaMdQuAtPXcivUNDPvEC12pRHHwVx+mp6thKssXamL0vIvomfmHNx0i96
/Fq//E1ol7uVSRi83BXf2WuEdQZz838DAw/XCHVlKi1cehVT/rPuzpXhxdXTttgb3u03ZfRRXHTD
nIb+GJp/wkFk70B/3eyfG6YhIexcN3T4iTwXzHdzt94VUEHU2l9KLqWPSimmE78rBVyB+FKMCauB
jlgmU8FHeAXM53YQgsx2Hn1fxVYlmgqyVGt4L51yZsMvFjThK4O2X0IfdusV7QaKfkbZ3rm0sra8
smAQUgz0Dzr4iWJ+T/+SOMw3gcDPkFNjK/N1I0ZKEQXQ8WVr/dwHOwZ9l1XjygCQL1y+MGs7DFvN
9ecFps8CQMiqFXMpySRC32nGTOrQeIB5/n1wk9tbatM8aKdQ0CnoiHJPEKdFqGEPpsMpIt2pTjXX
7dbRbqqeA17DBh4g0oXZqbFd0M7E98RXS12RmCJe3MJwpRnpO7wQx6jpx4eS+F7MyBfO3/6Ivcfc
xTb81rg1tx2KkyMFGmo36wR6m0AuAfsWRQj4yVyaO0upDGtP6nLhrHhmECLUilwuUOvQMNsgdTWu
0kujvoFmwoQ/U1b3UJYyI3KujESh6EVu05LSQbI3V9Y8LrJVQMaTMfJjuMKZOA11nBShMafHTyFU
fm4vz6jCEMmO6zu/aPPkAqynmue1WZzz0amh6q4hHI3GbhyMA+VHftc9BFV+lM3sTV10mf7cS2eA
CGsDuyFG+EvuHTi7BmfxqHvtfhaer8+bwqR699tqQnM3QcM7pOOcuDMtJuG3lT5SA9Fd3lb7Pvlp
7tFXH0fkb5nA6kPOP0EaacJqOFYAT4eCg8mxPlRcjmd84x4jYiqVrTq/HcTp95KzDA1l0igLoE/w
tRYyGcEdh5675W1I6Kmhr2ALVbyZByLT61yqcvzvYaHNOGkLr4w5JMT7Zp9/7Rp7ZKmG198nu9YC
j3u83yz4zEZIY7Zs5GNwRzTZL2OlGPVZPZV0UE9WGVlKcxHcCCCecr7SotLg4EZuiLQWVPvfNuVB
bmL6Saoio78LARuGJyVXLLVQs9YddWIUmwYS2sGv8e9o29iCXwd9cbyZSRIE/LIZLErvjoZP39Xj
Sh0Tn23ggLSph+mKnbnACIV8bI93ko8aUnHmrNzIgAXUuykV0jiNrN1eiLZdGLvx/Jf9RJfebj27
ZraYOx6HwysRyvvjY5S84dsNeThP3CUo9jdh8HzJUV/sQNoyX628NVgx/ky1pgRi3AODtZgg/Fsz
bZVtPuYyvwI2Rjsuqn7jeS9Lqjd3O313OJz6I6RGTJWbeC1G6ZvW/7kBxjcXIPDyLe3WldjY/Tfs
4sXUn0vvAUlgUO0Fa9aCVRK7FJ3BRI6dPgtJdSKXGfa7lg8O/oHmR0PCfVNo9lmPFZjN2VQWq7uY
Cg55kh6Z7pl3SDKeLmqJPDWoexFsGZApvHOZy8Evh+kax8iqEFY7n2KapQQFxVrkRewkr15BXSLN
xFaaq1ygWUKQMDa/Hm0zc4Lq85/mXl8my0G5gfiBdgP8UtH83C5dEXdHLGm4u6p7KprE10LAgsor
1ekCXo+plGprk+uM6u8VhiFkDIBVsyNBJw2LgMZkuqbvfVXrL/qgRV30u9XdSeXCwL3OvH5gyqib
dHMgVp/9E4osm4IbvR6sYvLlPvFxV0vpbcswhdMdvW6UQA1JVOSjbjIVR3GDvh6fY2yB2OjPxjQk
E5vyp6tgHN/0Uu7EeLrvKr2JB7ONW12EWkv7pGweXxl/sKQaFGdWT4QnvL3f983dDA8LupbLUJAY
pfoiPidHO+qwtu2Bj0N13HLesnhtSSUOcIIk11yBUZiMKBQiCFqFoodA7GotxmVjQycVyLeR7YBP
MajExL3NH8Ki96jda3EyEGy8y+3xCgfp+aNgl4UnTOW8qbM1VMLfvpBfCLjlMWUD/qwA6pPR5re1
c32CfPnaO5cKHF1DOXacHgFJ8bbscMK0OrHf0vp+oWEPo1CtEOOuYn6u/t59PE6CwPjYwa8q/tz+
sD2plc2D5zeWNX2ndXw5TDfT8kHUd80sLeE3LpXSnRT+cNJg+bntlFaghCouZ+m5KpDkFFMOZBbE
RtPMehcJFgVgg6oX7orP3R1mp0B5fa39H4f8/ZO1GJ80JPzj29o3YRduEOGbSnBOgIEQqSxG9Q3l
fQD4prhlrDiXEl081fmy28Duuke+R+6eW11DzQWLj2QF02jftvGPUwqfvLHIsBEiFbLTRguzdRxu
rnAU/nPvNdQqwzX5aNTmbgLgxRnfNctoOgtf3PDAnb1m8UH48f0XzEVDovIDyUok/vHQQAFSKVFN
p1u+bWONvoIgpG1AcdsHLKqov4HrS+p4FziVZHvggVxmHyq88Rl/BRJBDJWckKCBXsfIfHUUPkiL
dpwM2Ig44tP5/m5Vu6l4dp9REXKN2zaO1LkBAXNu885WJQLL49QFIqR6+FxF6UOJPCFdjYftn3OE
mrsyN5wfGGL6d1J7orBu7ziobnWtxv8o1aJeFZkmGpUYPNnIcQG9Qm0+oMMxqY377ZuBB/rHPRq0
VQaqchTg8+rCJqy+sRIUFu4Hv7wr/hojaqMA233qzvjU3df9Pp6KmyaMZsf77gHnH+I74iCu60j4
y9vEnJujhDKs/vIbtT6vIybApB1xCDAMe5C4p1vul/pg6eT4GmqlQTF4NDy0eNMjPG3h/OHksTwH
EUkv0eXsSpZqw0VS98UE+6Zmn8vrocht13KfpxW+7G39iFnafKaeNoM1USMrms74/eka8MjkoHTr
6o6QT2tMiIPzUIawQc/ZKJusc2I7DAGWQvKM73TF1ZmV3gVT+wgl98zR9pZIe2erQS+oIZahO/PT
KuZojyRagiyv0z7uzUp+46FqBU+S0eEO9LCPhNIhMRZNHNo5Giag3b751g26/t2WolVXrE17ScxS
Q1WgVq0I734uyA+4/lBkayWIrgbWWcWjjmwRv8ORsCi1FKNHZkZCcbnHJdOictL2NOoBjEfn6vdM
bDTkFuqUA45bYKyTuuuQmxaNuIWHyd1u0zJL3yp+rDNpIWNnMdnCAnX1IGh5ckax6mZpOgR1m7q1
EFGP+rnYSy6BAsG3HIj2Ku8r8VbXE1vMignlJNfvCXXxCpJsOLVbJ61LY0OG19ZdkJ2+E9k+s9Lw
5wkzf+u1Is+MdcMrIQ8AjdDZg6uG8mXq+DG5U2HLfsmT+pY3pv8nOXuSp0kONUmVhysLHv1+lzKS
/Tkgf8/uRdkyHNEWUbsXhod9do7esjoVzazdrfDPiAAsVmmYOUlrCgXvm/DIxTKPFBeruzpidiIF
2pZ/NWsVcM34FaHRflqOAFm17nr/NdVSLjNExGYmaqMQaS2TmC+3v6rw9x4jzfMjGFzhq/pJp+2G
unZLf1RuKSZ6bRlO9mIFizC1mPJXlIbjkiOPKD8mxAOBJdqsVZLUe3EPV4aRy6aFmsUBOKvTIzck
fVpRMx7m6O+3TDVikCG7uoniByNveOGuL3UltRVdHwZ6HEtJXg0q9lR7EULKA/tbSJJnFHRaDYa7
jaJuv62rGxDyplTSij/zMlMmCSVhYB66Q6qY+S0lalbUbLt4R8TRw9vw7xiyVNt3y4eiIXurQdOA
1cLcwQjLWb/Dn0TNSPw5P/Yt4F1xbsVuvtiwKpVw3nL3tO1FVYKcwCpzQ+W+k/iuYpFJbMWlU+p3
Bdm5u1sIuGrbnWZ8inCw16B+gImaTnaUEAc5dMHS9gAi0TZaoMu9T/ooMDFgmHp1DAwyYybMX/ya
A4aqOrg6c9QEKNxdi1QxITBbY7vBHfj3r43FshNm81MXdJ2FcFwGdpaPdl9yLfHuaM+SMcitIeSG
ajLJhZab+nZpqDGdMy2Ovtfe8cm3vJTYHGZ0rxD4womr3Cch7CWB5b7FUglVDDuOMQicqztBiZ5t
LyXuRGQcNw5I/6EuVA+DBchU6igySZpKUzJ54Rk82/dM5mD2TgEVN1nIwxOChCNjnVB3EQO/fAZP
fdyIvf2xj/9vvXxWhDKBxVtIDsoYw4nkU/ZpFLXhM2rKk4fO9BhtLhVPId2LHpwT8HZpji6oRF/O
gq1mPTez4xGAV/PQEEBnajy6AZulFFGteRK87ASV0I6iEArhJX4UUu+4aiMcWA+A+zimMrxdt05S
+ARiWLQKwrbS0SqiTR93jFisaOWmIJeto8IKfr/jTrkm3NB+zV8Owdp5xeWZCfJeHDzum4ZhYQNR
J5x90HPsOpxS2GzV5T/5GAMWFrkCD2wAfKqGYqYA4YYulkIKExt2R22paDo8R9gje+Fi8MiKXp4m
qONjm1nKQ1VRL2h2R9kCzu/C8nsLI9LDtK5Xh1xo3w25WiWT+r+t14XObe/WxVL7FkV/xrbf3SMp
f7PwVREYY6fT0cMIqno0vpLkFvsc1pIS9KKbyGsA9+zZ/nqrZzw+8R0pXWoop2VbrmYjWSZJHlrS
TVX9aP89TKeg0GiVpGOF0yl8LPFfCRGH7+lBc2vGTQjl7NfrX5ssIxpfyoFcc4udIAK3+qdKsuhU
gw1y3u/bB4RziGWtFFoM//nk7rBuppJ/UnxwQ0l0VcVS2JVNqeTJP7QpAlrfP9I27cdxgnrCyRj/
6bwDFC1VXu3pLuEH65ywIe4cje72/eXW6D5SrM0AY49dNIEkTvqN3+b2CLZL0hzkriuVLfzkQtIF
ewxjkEsIhvJyTWHgDU+1PS0d46/GnP6YY0AS6u9s8c6itrY12hLJyequLhL6xHgFd6i1FSORbKMB
V1WIekNGjptk/F2+vfL9LFpgoz3G7YHThuQ9r5WEBMStWuC6BExjuz0c7NREj1qH8r0cU8ldmz8q
rRwnmp0SYTHQLyCJkjcNKQLRIppvZVX9JOAqzPeIrjO699E000rT65NMRg0q1OXa63x3MU1VHI0M
69CWT7aXykqZfQS6/JPC/kFwHhrH57Mh605BVqQlz/bGx7LVWQYBswNb1R8ouNxgU2kTJHOefad1
cX4X5iO85pqDeamoOPUv1ujaG1FDIutcJLBeBCRv7JT+9vEsnRVaQQBiq7J2l+imq8hTaFjeWweW
Qzq65tKzSvRMmTH7e5Uyr5UNPU0KAS717l5eh/pFBR2v8W1yUtOxBHSBNbHU+Z4mW6G/tdRc6N3F
NZhkjpxONzGJJVRFTWny6QCQJdu7KDIiIQMFJJGZB2O2Zi2T5sZxymJOPHuJKWJyO90m6s77fvqv
MotxzL0K1lsu/SYdkO73jt1zdl3ufZZUYGMosG2a/zmNJEjLWpw6h8MO0facSZv06LYuFGUBIWu1
0teANbhvCHQgTDJpAGsoAFHntXT6p3Gv66P8zQWQQD9CTOuEiYp8G9okrYqcVmTAH8Kyy1UAMS+D
LUhXRTG7TksCoGzk1o8hDn2UixdAF+wbt2iHpgoM8Ii0+RBKawAU1HC2e4lUSz/ZNr0sXVvwgosv
k2RdQnwtRPkLaTTiwoAHT0Xg12plzZS+1GZjH0lChtiJFS0DhwGMse1whGYB5smDcTxtnj9YAg3H
rrLNIGPy0yZW1XbZgHuivUy9CN2IT5AgW2bVkGbo62BNmQ+z3kIQK51qx0PAcWPUCTjNZI9HDHq+
l1qVY0qjPTKvgtFzFVe/zpTC2ugGqTqnSsu0kevkN1C+D1TuVmp+Kq1LWcd2KCAJ+94xniopSUwh
fDsYAQlZPo39lPTcn3SBQJ2c7xqvejy99k24WIaBCFkydaff6+LWyxBJvjuBQamz3l9iwajuluZs
YR6MQla07Iuw9BRXFbblrJ9tafRPiC524nkb8TP0F1Kyv1PCnSlwjS0PRVFjWI88DcO2keXDTJgb
CrzD1yc6e0AbBAzGTq0JdvXskNWMBAQUZrMvXIdRxfAqdsdHYxIlBGz9Zzu5o4DiXzeFHt/m2tat
0mVDeNhmnlU2IwgSeuch90K/HM/SXx6VaPHZBx1EpHwwMr/+Nl9WMEoWwx6NPK1nP5caxy4p2MGs
QJ1fdH+l/rtGlryEHrg5MNkKRSJjszlegmzerKiYV4SsFStIqWJPb1pPRV1m2SdROvtAqdNAQR/D
q4AmUcYDzywVzKtvqXkp22ciuEiw9UOxogN1Y/msLEGJfO+WphKSYk7pbJD5yudGtWwB3lkcguNI
gdMXrgYUgPf5RRtgu/KIvpuu6Gw9FxQGMtwIFEeyvtuh3OMhSpE+s4bbPqYQjWa8ALS0iEdx6nvO
8oX2xraWVtGuM/GF4e9YnuCN050JtfKeit4e404HW9ksqLUACwRxJZKlxWVgT3GGUneESk+RYBWj
K0QD42alTocgojK6c28nB+jll/28jIPa7unXTuTJUpaSmatGIlOw5djCid//sNoKCbgvBWxy1lvN
/hXH72LS27KM4s7SHCYZnmnjfFe/WTGTDjfyDCkVGpj2jsqXh0uyUpt9VhPxY0koL+iuH8KoY/CC
c7cUB7I/LsmhHE+Cf+tvnW1EGmche8KwHZi6JWjzj2v4J2nfhjEfEe8HtCp34x5WpV+zSodK111E
bZsg233+bEoinlvou4PDZZj8pxK4sL+Mas1Rq8IwPdbf7ZKBtGXLY4V5GfuHyJIk9AZjcV6JsX1+
6t19CvGmiDON+aGzFZ9h1TuPdhPvwLHlh5yUsL8zna2uZ1R/XGjrni2KX46DDQqkmmmg57w9XNLe
ToLmLNho92Hu9MColfWLoPNFIGJkd3jOeOiinIApvBZri/8BUaa8A6TF+Ejm7Ethwd7O6bEdzNiq
kAwxWzVjeKklfuY88jPCVR5DqCyCbO3VO2T08eNcNkpvlY8+b8gjPEo2qHPYCbsNoI+q2RiLA2Ks
xY0LL1RUjmCJpdKG3XaKHzDiZ9g27Ko3KkVw9Tmz2U0ZwwLUkj71StV2E0jl+oiXMLQmSdoMYL/f
nIkdwFEppch3S1Ln9w2xsQ/mNwI9arJssswZbYEGkCp3fgRKHPhKPOymf0oXF0hRwUWUZ+cA8q3m
W5zOO2s3+bP1Wkvbp/7ghVqAiAqqr7d8///Cvgq0h5QIFzQcjQEr+B/76c1efczXqbZBmKInCk0b
Sab9noLWGjvHddarAWu1rdgQzgt0Wx+SRzGRBZze6lcSLxNzjLg1tVcm82g1jceYT0vENe3ocH0k
xWeGoF62VxTw/3uSSIM/YBoQIDOmWXXoT7IHXUWrFFmJNl98H5LJDnJzU2G3fORTWeTnJIc6CkS+
DLs1EkHv1mmQaXFMZpz5/fZOSsE2bqCYjGQVlKEEF/c6AFzVyNcMgpFOaLdfqBOJAyXJyw8sZ+Bf
tCp2xFpGHCPeI2A+VXMSU29/iDvwZ2I8ZW77I9sJUjo85dw7XgQSpkzm/v8voeCgjqxrJTnX6f+x
o7t6YUxXok3gHDAsMxbAIcva/BRrrJpfIRg2rkClaVLomCDYXOUoHMr/IQ+lbzT8PlSoJ8pmm3pB
XdEJQfcdjgkyu0iY2jaCJVjndVVLvWWZ0zkOljBMTZ+7FUosYEeoW8J8HtPHvV3qID9wjDj8zsD2
PGLRDV1Fa+NFvBPpgJktgA5HWtVmfUtlVmjNOrkVJ36ePHdkZTYqkb8kWgdwqHM2A8LKyb1JqOj+
VMEsTviVL3odOVtfZ1h4eoc/umPkAiTXvn7tkfC0n7aW0/RwuCev3Dy5AzGhV4uKJ8jTGFcaOZE3
7AAbCUg48iEi6HxdwcZDwwAzRzBqzJIhjiU7pVyqVFkPVyKXpZhgq7bZNDhNz3wdaAki3Jjkaxb6
7oC1C5LWNXQtqaaWvV7YHGQgTca2DiZgQWApwLbDBHrjP9zFikhOcrTZjqLT/2GL1P5K8cqlUbpH
PIZcjy97M0jciwpfR/1Tz0kQOnEY/+L3cPPzlEoKDZqu9sjG4pVb58k0zYsxvpYUYwoyNprVNZpb
q31Q1RrfwzikkzGoemDoy1fzP9ybF7c8Ck4j3+iq1xoaDVZrsTsyZ2kE3kfQ+eK/BaLuSRFQ9the
gsJn/HOp5SWrGz/dR45nId1ntqh1Hdyrhq8iqaeS9iboUO/SCnMdIl+OsHN8u9EUZhJ18VZ0sw5p
XnM4K7TBSSGxZ8tn2ikozvO7XeiQLh0mqr6fUVuuhXLeMeDP8Vxtd8dahwFDGYBDvZmPhwgMPmpD
sV0LAny5z8hucGOVZ4HJeAFRI79NixnPEZp3hTWY3DQRn/5NPFwIANiwXhlYevXHix9uLKUa4SLH
XXkHK5zIE06zp8AYjCCY4RZhpw/F41xzugpmudDqItBgwNCzQxgwQbXPl7IaMuAOZUA8tmUU4qjK
ng2hZWoxd3RjyNE9CLg1fxmmyS4e8XxfgpVO3o5GiSam2Fzow0nv4hMeGv+9lLp1LvzjWEHxVGt9
GioA9lY0rAgiMRHSA6WuaNB7pPVqrbo8LXefViGhGX30AQAWZksDpwUeNkaH/sGfU7vrwDz9hKHR
JBrETqI8zm91WitW+4KtagUWoCdlGyhj8Vr5XZJPc9qnTFWNOl+H6DPnRbwezQz7aIpTEKWJ+0Ns
7ON49enYu8dErS31SQyub0GrXAZZTWygSlHDXxP80jOmL0dlv1C0L2mEMZe8dy13onLAmfdRekD1
21odWiVOeGS9VM94NXBfyMebMg8eUqsOOtsbpFzEuWgjjEtY2Na5JCoK2wmd4RwjrnMLDHR9yf9u
jZQAGqGqetYByBPNqVEDZmm/SEs/aIE0QlYHoFpr72BdhqZzaVy3n0gldYV+/wEkQL4yZuRczpVT
QppiM4g6rwsCyCLAGSDgPMwdZLLFuENGW0uecUyiARA0jqR7DewLZ3zjzidbwEeWvtNL1xNgnwKl
QrHMP1sUT6VGk19YUJH0m8auYN6EgXnBSZpWcvI7N4fb8B0OyIOIRObgDoekMRM1WqyqZ6WY7iJ2
FdlQWCRuPynNG5XDJHWNZTv3JcKCDRqksiTEr5qdz8UNqa0vXb50Jq17mJ1amWuH5u7VVUFWj2l/
Om8PmPngLHHlsr6It4OIWu8QUYxo+sVpp7W+pnp70GatQB50bixxysTfGxsej+OomCrGMS89szv3
yIIGkTM3KdrrJR6MYeKFcA5J5Gf9yQttircGbLRywSjWYO0BrROSg+dQbAUCuS8aya6hBI31G6w8
WH+9EthrFVmuxXuAWOMfuOssmUPIQQpt8lhmYiD6uBo+pZI1mPDT//qsyJzr9AQ70CtSh/9GJTBi
89igW0xMqUTWZDWB3C51T5s+LUxaADdjiFEse59zfngA7emXJV44nWAMc9mCPYBRqE978tO/fFZW
qaDyMEqNnAXoy/mvhPsJtYhv5BCVNphzsnBNIVGt/ry/9rxnRkny6P+g6kmyGaktVj43ZJFCPhHt
qfqhqc5iknybS16u/jbNtRciqmhc5h/jywB63wXr8EoXurRUz+8D/m9ky8ztlgKt/Hb1BkxfLdp1
N9B4WofGxSaS3Syb2aavvu74eugvHsgPnMtEHVSOiTJA86cPjJywmwSBT9xo7siK4v93cxTLxoSp
hfEUU9Be12zjBIrk7jSNN52lFUXdBHK9y/cg9go2Ns8RK0w9ojBePaMpPWItku6vWwwcUdNd6241
v5tPEvWtdhjx9VDEw/6NCo1jeA/UcXNO9yvJ1JXN1EU3HApCpmTsOEaHqQqW3TZtPyG/DrfBpC83
PfJBlyLnKZCU6H0ngCL3jf8i5PPkpwTuose+D69O9biRiAjNklMGGm3yBmOtozZv52rJhgdiwrwr
QNBavVVjsxG9fXKiIVXNbo/DegxdQZjmCCL4RXpLT/N4k4tIL1Fdlz7AX1Aq7ozhp5LO43/6TrBw
o/EUs31webDLj/tPmGhxn+EPT3Fn2icGKNVdKAvbrpPkBywgLnkMOD/WZ+2XUvrqGNY19fMIsAqb
IcnnDt8TChjcAoPbRCUCnPcfQGLBfs0fxTXzWS0RjG4YvZ5oRy7SPvSunqzEpHqIu8bkW4IqVvy/
wUeTTAlmYY5WQd6gBZWM9c2VIio3kApcGzUzieW43Ds9aglPzEo3ODznLrA638YtBZFW4P9ap8U2
9Yuwf6kBLKTaRLqw9cHl//r1nxRTYBrVBv4+JTnrr+Mv8YZDPxCyBeAkGA/U8FCuU5dgb/rK9TXD
8mm8H9bAfC742KqDrBBNskwkF9p4vE8Dpj2kGnSTrZGEeTspVA4b9VYlerwLgYZ9mT0crGSY/QJD
g7vjMuSUdchsj/9m93GS5vgtXw+s+YhuCyRTrB89qOKPsRyupbk59xWV1V0oCaEprmgrhHtuTnT0
wenWLTOlX0xTXuLdhEsGRB8aCxGI84eU6s1sy2xdSBPD8RL7oR+U966FN3cgyCWdXvQ3GbZ3WTW2
8LH4/B/NN440Gaed6YGDITNaTRny+Of91WIIjxvS4hQ0V/u58XqbXZxRJunQX2MjrLJbn4ksFx+o
prSZWBOws9ebP/AtvSR6ftJ+DRFfbsjC7rG947HTMBn5kNivsA3k2XADrJl15rBIqAuZFopOJqKP
0jZRPVNQqkn2KEJJYjFd/btA5zyUw2fhDCpXKYwXTJ/2JLsfnY4CZ3IWGhzUwG6dkS4Psiw9eswW
txF9ZpMg2Aur+tc/4sRUCe9DfZA80fNYu0HLyesnfaShaboAQDrOgk+p7v15PIm9NGTq1lWXJM6f
aMMeN60dlG5tT0LMqu4ueDCxzBLDde6Og+XULKM/TZf4+l4fAEgL+D79K61BoxYuZHpcpRmjlVMW
Vn5nG6jf8T9B+AT1/plk8mcOhxcfNWbXSY8i09juJi0VdtxM4HDYHq+2F2x5HW9pjeC8GQm8TtK+
EhcE14ZHWZ8Dke6kxn8IERJW5J0oTUaX6RIePUJJFQITNrfruaBlJbUMrsKWTe4B3R/+l7q9E6rz
NPanTEjjhwfWJddLctokMpxZIyQ4yjvGXUrI2AOSfNHUqVbK4F6kR9x9ofimvlD0/2TdV6ItSyFn
novNmevYkFs8uNewOIezIQYcSc8yhUs/jmmkDIWOB2nDLf5R6PP6slN4GH1oFBTyIZg3Ji6f8oR8
Tm3Tu3/IzXqHAD9Nck3z15z9DRJBGuCHKmvafBotAhpVRzFnABsnk0/mCp1Z6yHFTkj1OfZ78Rri
TBpzkwtfGsHAxKXFl/JsNZg82gY2HdV1mPRARK3VB1FpF9eri6sOP6biKmYa5d0aTXGwg4wLX7Ls
X8fkk0vkxA3Ab46oKzC+qxNfPHSCgIo7cKfQ/Z3DOfPhnK98WEmUVlsO/OyiHrrFcQUwYBDPKqSY
Hp7BNRaDPNnPUZEmLMy3jstXfQeEjLwJ6vzImRjdy/r2HLeqvDzw7Z7pLmKsH+HODVQ+3GNkFot+
4KdBfa9O6ZSwrGexj1VyFcC9LQQ4abrqEdimTKVV/Vby8v9B1xAjJbVZ5Ijas3ASCcLZaCcbkNjE
UPYeisT74VS1jm8Xb20cA0VgvHhOwWvnagi1Kn9YvLTEQSvj3yMSqA9NogoagUSyR46a3tlTxywq
8miSbI2Nc6gB80FGqJbwu8h6DijG4A9pyFtRFrnW+cbXXL3XuQbN5+TTeDoVlzIW4jgnpW45+kdQ
Vh7PyZvfbDQeBuZhsX+Y2Izz3p5BNIMHwLMpDsdWu/+tb44SZRb4ji5nH0Jx78vLsiYXXcKhB364
hbokVoN6deWyWrtxtBxIvcr82XOXizdqvckddwyN9tzOpckTwZ16XGMmlVo4Fh0x21NnuiK2lmlJ
tG/dIiAA0lXgj8JZJv+A3HhoDUe0ZWYQK0plBjoP2FrxtH1RB+sBOu/Uf1cwW28DwABNaNlPJUzB
11vfr0vJ+b0wuhZTkQdz1b266Qt8qi8BM7JVmTFkBOWyKf/oxkvoqvDtBAE7x2xwTrOkDSs15ZUV
nOqX2yrVmESQrAuVp5C6xVSzCH5iUB0pg6dIH9F4eoQu8tlKm3ulaTFJLnywB2ZE20Jcl264X4QY
pfHD3yeig9aEBK3640Bxbl/jzVwsK4I77tNpJoyzTPIKsVWFQGfYYpmaVhV8jClZAzuwxuKTwJPN
biS0yv98E81mvHWOWKdekxMkVMSe5thEeCJKudZYJL1LIXcd5dBgiAN/yeOe7rZ39aVm24wmVDub
iTh1Y/I68a+evuJnXoS8VvXU/TCZMPP7pPuGwea2cjApevMOuQTuHJa9GwoJ6HMjsqDgsyHTBaDz
3pRw/2ov2fmWOVQfZYr5w7CAgK12fvbvl3UrWiIJkPA6UhaqPOVS6DiPwkqszEqySEeOqbi427vz
ZYwG/eAjKituoUydeUawpBgi+ch5HJ0vorJPfrFDTkx/vPw477NyjJlAlS4YvXUYL6u/hCkRg/wb
P92/6CxQNAA5E812auOrzOT4bSzVFv/EQvAAV9TmkMW5HS5MMLX9E72mCt7f2itNHvK2PpA6oM7g
TwuacnGbO7SzcpZbUaH2+3cvw9sIA7rTNfbnrvPpAs0pudp5XRKFtdTA57LTUr3ztQ9Or0xnhIkf
M7a8IBtT17CBeUglGJNr3HP5rk+Z3JbHFigQGZ9v84jhCy7ERRZtn1avKg2khiwUdKFB1sMVo3MI
bJq5W6edRvg31pwgsRRnO9PTfROskKJMwfeLnlg/0jkflAKYtmTv9NCIWNh0pZoUya9r/MFrBYI0
8rBLbpAmzJsVjeloTLSRAIfzBX7USrhwJg7V0YLkvomPxhVCWgHMG0xiBAs8KExPgkNIxQnpdtyd
wWfXeu+pg39CchJpTYivmtdxpJQh9m1DnotDgA31PIEvtvQr9IU0Z1KtV6/UHboEzb8INE5vkBmL
PPyJdh0Ve5muqq9O/9rWS8uA4CGwnxBBTJtbO/Fmo0djLoxQ0ELcb+D2wovBWpy24MH3IbJYjvcs
xSsHiy6qFyiyQMGTTwrSyQXAa51DRXVbTW67cjpGnXFh0JMc45MWfPuk8lQWN96oi952e3J/pT6O
dIJ9Rlv2vs9ihjNedOobUeTll+pVUr3BEPAEhJJsHSEnSpCaU6oIhqAK1/XQ6r2z+sNGfG0UCmec
Y73APxKfyodOnVcW/oAjcLv/ADMIIcmyxZca9mpsxG1Uiq5Xt6PM1mrmI3Ws8WZuktEIh4xpHvdC
2ESZcyej1giuJpPAIMwVxtsP5yjCZp+R7ybJJG0PN7NnrbcrT086OTEau1ErMS4zC4uc6T+aNMPv
Q7BTlEqSb4w8cmi9lZut9VwGK2zf3YS+MQarredSskBz1TTtY1r+jiXHv6ftCDDLwvIN2nl1iqwG
b1tti0YMBNOOTpi9QPnPBs6GABv0wqKtr/sE49BlTdgaLdmkp+DSq31zd442JaSdYCgPjd3qVwAF
eJJee+4fMXvKft0YJyD6EDxKMcvLX7DyF/mHA5uIoz7k/qTz/iTdS4MfZz7tp6LtIUjwniXKcqPu
u0RiH+9vSeYV6e4K811IAAV7gqNUgHJJWVZBpJEh70I0Y3/msxzGopvXxnLTpwjeo/I7RSnDU1s6
Mxg1ITSjHpSQz42eHIme/Ss2b3t5LCoVMdpNbee97roi5bVSHyfTYjbCBTj3KE+XuF8Gn8oDqnoG
/pItfv3uaX9tjbSswIc/Cx7jF/ap7VXHUHrcd5p+updEpXe5Qhr1r4p6HOhw0UN0dJm/VGXp+HOs
uxwSC0Nv+ndI4SUvGSIWPUkBw7GndkLyH2agBhJk56k6b4E3hl9Y+Eole8WDBLd3oMgPHXV6d5d1
ZwhbRdeY5G4BpKEmeRmv8T5U4xTGO2ejlL8hVxi4bBd5yZStcFmYcyNSRUGcBnAShszRcyVynMc1
WxVclGMZ+YUDijlXc0dWBlRKg68dFFksX3acj9yKC4glZWtiPxoJee9mfHf5CKwYhUiPpxboDQ+P
LDeDe/nHl7BremRm4VrZhKJv7Ra3aAt3qa80YtONT7oR4cHu9qqdkT44XRyT572dxg/uFCKhLZ/5
YIQ6/XudTxh8zX+V7cKxfJKjMUfyjA1f48DFNbvP7AoYsYuh5Sx3Y7XGdx39Q21w4NBUB2MMERKo
wANGz3Jx4yDjqJi0R1aSqzK6WUUnrzvSwAGgmBbqVU9B5HOhDAKv9Z98QLGWqaYr2ljBT0EYuICg
6WDpknF4XsMk57gAWalk3O4+16BFnq2oW5BSO5tlrItLe+EZONRYUeWBYwl3SyEF254TdD0Ib7sx
8qGnZ1fka96E33CNUPJABoedndgJwp4ejlJ/7tWuOXC61fcEJi64ASs6TOVUQEp5mNmXUDlzsvgy
txO84LuqrvFpECwoi9IwHmXL08Z6ScCz3oKKXlF2tdz6wS6WmSMJ8nOav5Xv4sUibsRGS89Smh8u
BHC9f/Sms1cZGUGuMgzFRbclQCRd6y7b2JZcPGEodSyFJ13QjasIxYGZ7LMGWtQvUkEmsa1PCdJa
bmqkWYvZ17w2N1a+0IEcAeua3+sTl8+QeMdZ0agJ8+KzumLqH1AY6JilD7EottnbgyAiU6+lBqDP
NJvQMJH9EgzGXBrtA0zMgHjZHZ/7SiwEj6+7bn2MGE6ftUE/brFh8UIZJBMdZfKkx6bkKtb4wfiW
33Z3FFobbN2CZxyAlAS4amKY53+3KIEp0FOQM3ZoP2IbWUjlo2xnZDpMgZ7/FXfStlgAtrBV7ghF
CMjK8WB7LYAppvaES3Bt3CHnUEqcQw2tpfIo5pnlzRzpxOP4keVnHB0GbzUb3dC6M5Zmzbt4zHB/
/ximkdyFByiRJirvHT8SRk/GkjeFtxoA0d1AXLWltJL6+b4xdWfzgTeVdMO6OAjaCNQtNaohCrnj
25fznFVMo6A8MrJkH2M2Q/JoQK/MSwkVBpzfWrUsrfuB1HyP4eNcDp4NPOBUOhaRkUFGz9tQAqMu
0hSCAB/ec3xINW+3ShEZcuaoCEKOFNc2GWxAvARy6sYPxPoXDxGMCycAky/E932iii7ITRXN+XYv
oi45tVd3Chr9VU8X42XVQqwbI45DDFl5yjTIwh1vFpGYPosqNCexLD6zxeFXG3LPTo0UG9tAE18H
GcQXv2Aijkjj/6oFWdIybZEjXQQ/0oWhRHixiJ+R5oLybpeaS0pKgs+113kC2rJRQsVBTk7yg9Tg
MT+xWq3tEf4Uf+sDCDFGMgBYTVV0BIRjPWfcmOy9poudb5NwjZS1M1g/3QAUwCChWQMLP8h3gbgN
1XqcO2wigR+9wcm3DUNP7OLCmQRJfqqNWwrOT690KYOxeHMZm1FJk1gKq1LnFFh19YGng/1hB9r/
qIduzhB7rH1AcXBPZ0RuR8+SpGUcX97n8d41gIZ6dOUCpaEgHyQbSaJwf9/jFFBSq9nt3zIgcJnJ
tCbAspP+Y1mboMC/D9yPWz3p6HKMhswvvkN58B5FKKXvOk8r3lI2EftUYljhabyTQpdY/o7zYX5M
V9x/GBnJyVky5omBomQ4ETBMsxUIZdc45r0crEvIEDBNs9bZJs+O145R/rLgSigCHm7Bb5ImQTHj
ClnOW3vTYASq9rZu6GAOGdJrGO2ELg8GDmQC+homLMhpDtzcLUzhwL0OGkGq5AjcV8IzEjkeYF7y
TuwBMa96pr9Em49NDtowBYXLb1NIKxXqjadhcHjyzCfgVALnIV6MNFMrBwLRARSqMznr8DZ1rJJ+
skhx7CEHFFbQT+2jgqMwmuedEasdxptbQEIdRPTsLGiHdp68SdF7vGKuIe8KhuikcCaHvDSviUaV
b7Du92ZGkizWSHA76qUx/Zsu93KmfYLvooumlSdudxM2gh2ezM0Eh4sZ3aKkR5yZ6NryqYkpZH1m
qH34ORfB4m5Jc9MpeomI+GX1620mdbx+DiWjNmT2araVDrxExlar0aGvAAdnR5XzQPxWKvLIE46l
cJlW1GVV8A1DWOXvFOY+b/Xfqe2Zc7FueKbPI4ctL3GgiRzGKMQ1DYVDoCcXgQAOF9vmoblchLJh
5cWtbHrGhEg8dJHC7Bv0qZ0IxsihmQVn/TH58LgdEjv9Hjr74GyapnNLmx0kcT4hkO3RfyuZSSvQ
85N5ggVw5vbZez9q8BZ9aetQvIvTG6sv7LgrYpLVkdnH3KZCC3BL8skl5U/qElehpN79rerF9o2o
yapQRsBZekNx1JHDtaCBnKTSXiyK4LRU/82khhS9Ek+1ny1vAA24VAPkA+WwTjeLJYPZR+sB8Plv
BBo8s0mwZKck3LdBNdzH1A5mIZ80G93TPjY3hQcQXjWxkzvu88bIINH9NODcIFb0k+XjVdX/TE8l
5Wjs9pxdpWLsR+z8zIMbIdEptB+4s2r6qXVa4vbqzFcK5A6fNIQ0Hfuz/nIhg7y7WB9QyORmokxr
8DtMzyGDJcW2EZXZulj0fojsW1EEoECLfBZLmIgBryzoAIlbbGyncgL/hDPjuyPMugeoJJuwXg6Z
8YbWZ5IFh/RRW+NI2r6OBlyJdKgjjGrW99yLUE3xfYpTDz7uti93sHwyM7f4eBcD1O3ssFWqg2qT
KOADZXz3m3RdYXbtAQnbslJWq7IgfQkVq+R868TXY0jOAnWiJVMt1n/WgopakaI9v5VlOfQW8cPG
me/4Cyvj1ZtuFQ9su/KBJhiL9zNYpVsYTYq1HaKgf2h890ZLvsWwlQ0VyxIxwYEoWqYCa83P+ysD
+dkwy9qnUOxHra7MJnWh4G+cRx9f+ou+bmkrjE94KU2/uprcy/JvGJzCSwP80z3LIJ+ASBCNn8YH
wY1fc5v34hkcJisMl65sO4hb95BB+hrUV9YRTroAToJfi9YPm/ITxGGzMTJ89G2rfohk5oFPiQaK
8gJsWhBI5iaM2uzYPFH+kCW/GEIvb69XH0HkRCVmlPeRPjMHkx0Z/1EgcPAW9k2Q4PB4bhcrCYxH
GJvU0Hk5RkWx2HiElfZvbfdGSD3c1dnHwkbt0KC2fGb35VJlokIgufgDmNqEu793j8LEI+p7cSGe
NNt8/j2e2H2/CQ3Utc0OUkNWC5rusbRk5IVcLRzyHZH5IrBmZJlZfWaym3HSKCWPYaEFgFLRmyKr
4wWtRhyxaCV54ej14RbMWG+YTYx/51Q91o9YBPoIh5qtHwTu1+Ka5QS+s5WtURgi9XKorJxZhr4d
GG/xNgIrflKZJGtNbfnT+4ntS84JMM7cH4I1JQ6GwnEvzv5pz991wU/9EMBvJFJ5Q5Iyq5PdrQtj
sUg6L+GMDvCmKOXr/3+tBMpde4VzuvnvIYExDpqX2ym7onjdPvPcpaJe+3n5AS9zL6mMUU4jx8xs
n01/q299Sp2oC5vS12WtAZzt74vX6xM8ePdDRcUaTMolO4z7XvCFEOgQriL474SXpaIlfJtJuysN
gAyTT012aeSnZRAvmbPHN6mvVXZ5rSdx0w7UAuXk4P6MB4cMlzU7SsBAuJ7s+ng/SWW1A56Z/W/F
svqycMhHrKkL3Mre28WH44JJgZeTusOrUeaMfpV82kdbtA9e0w6KG0uwSfcY6v9pF9jcQmUqgoOV
x5tX9Qjk14+gz9wYJH8PHFWO5t7yzSi3rIRjhCrHhs1TqobJAu5PHUvlEtTl5uOHI8FBgi5Uraja
s1QkDDZKKZg8O9nnKZ/16xWdsJIXLeqCkJJm5ZUEt24/BGuoMk2zX1gKECtPGedD7hEAtwoSQRMc
+KDSTmY5Xx5trxbEzX75AapA8hfOQbrNPgJ4XNlL0QqjIYbjHY9+V3bN5LjojvFAshs0O2Y80JQg
mPVwR6oc387TUR84nbj+IYlwbGEdIyx95WehSOTL7pq2/K8YBoEPeLAYRHhJESTsIDAphoXF+2Ru
NB7wjw/71CzWucNpulqgJjQcX8YinNJXJ9AZhd4+ZcH7elqKPOujh6eyzkF8Xj2809aIYdT3PKvz
jh30KeK71NtEj3r0am4uOLqLdsjuQnFFeIdrWW79lUylt0BGZdLMXWWCDUhqS6k9xl4BFGXVeLfO
tYOC5AofN7ZYDBjSYj1DGVrgNj/J6N4ehEgsCFOn7W2fRg4U98YaZrXXKdCYBMq0NBzF0sC/hIpB
HCgsg62MWw2cnlvp6Hu0+zJ/FHsltAS5qqo2rRsdswU1kZVR0io38BWas+yuLdn7hIK9PpGiDTPS
ry8tZNcir5MEphzeyN9vQyf0sEfI5seK0RMTd/yEgw+lvbIE+aXi1sOGjztzksmGITTK6/B5WYBL
fsrahj2NTDwp/nm7dvXnpnzH+m2Df+VqMHOel9UNYLU1LApSOBEnwFIeNqUP95+TnsAPK6TQKgnO
jTV8k/2I/fw3+izM8cuX2ba4m0Iysz700FZLx8tk1NRrQplTYzgV4IKprXeRC5C5Pt+IVs+kC77L
oXrJoGEseEjSpYhjsiiIRtXWrAI2ijmaWHhsy+pEaV5fHRPIotdaBDq11JR97jrd+JCF3kW+KxN2
HylATA3/ODOqfmxIbHRqgdZqVYM/Likvn0YWSZMEwpvFaL2MFfsV5WBT1xqEfDMg32TPWOL07PpX
d3dJGNrTCnWGAj9vUYws8Z8OqNm7wSJ/Pkqw6j93OWm0g8e4OikRxRp7xve4Z81kG6edGlVktsj/
UZ2qtDLb5jEOALlV4xlCichD66WWJUOAs6DDpAHj/BPkktnoiunDU7Zvs7NlY6IdP+4xOU0wUwOo
rYAoePti/n3tXsWW80bkq4S3hGFFBufAb4n7SLWX7kF95yy+ELzHmUL5W22S3erXmBYYU33/4GCr
UXw37UZUoQn0KUgArI1Sb6m6aLX77yv4GGD6ao7zigCqqtw0QkgRj+abxNIIVaBGnIhMxP5T7xrZ
peCVwaKhSXgX5+nGBtlt3ieHnFad9ACfrDZQf+DvsqpaTXrtr2Hwc9ydmb4DII0ldLnJFcgsmnoe
ye2NJ/dYhXDCYWWtRszwnMZ+tvuQzhaPtppCyoA+2ynpreR+RgppoFtmLdpcnHHVkzcmIwmYkNud
CPhkIdbDnCwFwL6SIJiHW06K4WVTaPuEX0Fjru5KtnocJFVQnJwov5dTd0EEdn8clpiqqucD2QS+
7CObv0Hki6PuAMYph3lfl9FUjxko9gV+SjoU0d+P1iK/P6x7Gqqc/D9DKJShimLVn4wIdPsb03mX
yjfJogJLt4v7PFR4paC/Te4sGjg82ZbKjuEHKwRm03+2SVBbZGpowwvVf/NzRNf6+EmtJcfCQ1VF
/SSEDkeGy9WSqs9uMLlWgcI8X+OMzHcmWENsBtQq2LIMuZTqR+vDgOloOQHRkUBeHnQybbVm8+ci
WYGE2BStzcPH1gz7WfTaKVdu7tEFjoPUKYG5wVsfCE9wf0MRL8b3K/mp7+UT6ThrDeUa1jvfN9ZA
/gdxLkTsxCQpvSLc3dDyWhArAKciv+LVHW/ySOOFaXo01hvAZ/AsshNFOAMXux/aoslPUqVws0rE
Wq/CKfLowplPRapFBOBzja6hkwo62M5XolX92kBPDPwQlUxl6v+4zN73dPh7z2oGYCPtANxKgyZK
gV+BdKBnMZ5RJdV1ZValB43DgP6XD/LpGg0lGJPMp2j2N1zLVd5Zf108CQJR4oDEYtTfN8pm2DRZ
wFeovOYsBC9i4JehvPtOHPPosa2nNuwgS0i5uQScLQMcyq61qv2nOxfGBPnml1Ar/X2IThp87e+8
l9adCXBzDPYYpCHSNMT7YO7fM6qWcNjZwV29Ir3Xi0G5pmqlqejOj8roqs0RMhk+H8Ns4uGtW7z5
wFZxny8pDB54iBA0BrhSoSYEcbO3k5BLsG1bhTXsCU11ZfjEkPAcYVKB4EQk/k70LWQjPbRFSdFv
8GyjnJkJDsieEmXn1dS+hgu0GelbmTttcbG6NYZXaY7WiV2Ws6MHI4HBeQIH0KV7L05Pn0tAdZQa
0CoVl/D5z6Nj1LoKPMPP+ytU204pUemUbCJvoLZKZnkKjkWK9wEzq/sMMnClEjDiZZ0fo/Us09//
WeFmyljRH8NVOX2guVuRo771NK4XJiYrE/upmcFBKRqYkhCsoZyJf4z/Gmjs5j4Rzkr9Vc2vUR+0
nc/R2o082xP17BiN8aIdynHUu2P6D5D8KwWBQ4FFqrd7Exyne8Zyb1XpRaXMqVp0sFuBK9yqsBv1
7wb3w/bosBO/9KtdECxMclnasotYJ2g/71LtZc0qMSmoZN0Wv7CjeZDAzgjhab4TU4csz2FEMaq3
zRw51IZpuy0sGtTn9L1NtvhamtiQS0ZWvZW8lsRFutvmfWD2Ez06WZwPGcS1srGHeULar/rRn7qv
aNqvkUXg6Oz7zZuPO5Xus7PAeTDeWApHBawy0txxLGXnClZgJ+MAX0COSRVQR5/h6yLFi9GVgIFK
qo6lzgWEQhgUVLtshMwje4sD+Bg8wnxRiL7rlYjkiBV03tEY6wjR8AVLS6/i6jfTMpp9O1e7VmI8
e3btl9GJLejT21UWVB0PepYnTzJJDuuhOzrf7vp042A6Ii9BTFkgd/8gxGl/4t83XTjrh5JIraxz
Gh+A5a0X8rf8Kyu5tkMkFWnt8q48cTTK+2ay8NCy05LAG0h7sNU2Ir5Dj5li+BVMA1uJc2t4Cpjp
4mQFoWwA6vt/YA/W75QoKun7zWGTsaAfmaPMdlEChDY9orOgjbNEHh8ULZkusSOyJbC3mKNvmy8X
CqpzEblyBLRp3Jsimd1KykqBNJOPXAE+bjaRh/KT3TAH4R73ez7SjMJxnhfhEvHnwMjFdnSzml5r
tmNzvazYu+Jh27prNLb/1ua2hLF4DuCAuvy1ysnNGifIYCKrs8R073mtno9hiAci/s1MMZWSyDBB
HD3Sg6uzn1hvGNrkb32pQ8Fa4vopDihG0DM/Rlpg/Nd1CMvJk1SM5+17vX7WOdJFfG3Ecd0+GyT2
i3tE6nleCMKVeanhJj/nrp6X0OUgyfBUPvRpaWaCSS9ZPwJ/wxo+nKjbIv7nCPhQb9j6rmCGJXdN
NNRWX/e2wuQRRD574PoVz/UhcIXRLHe8b8TUe6fE5J/3rXsV/KlCFMeYcpi4FvOUPsXmhir6FE/Q
N5digM2wQP+xJ0crh30EdeNUmp+Oxu/H1rV0KSd6AiW8kzG+kW3LvOHGAl4mj18wJgNhcTE1WkN8
FbskiKngD4PwKvNSU02J+EsaOpBeUCQiTW2W5pBfyynK9g7U2Z/HCXdfged6/yvB3UlS/asDVTzd
2GV+C/OavGK1VMS5WhwqGQGn0oHs2CSHLX6kUsn0v1f8m8LxPv3sCWvB+fUKoqeac5u4ngPtDDeo
2m0mHLQ+TkyQS0fa6c3vX831P5cqy4TlV4o7efSt83rARGGPn9gefjOMB5A9qz88T4GLapS//xOQ
4EEPe4A3baQxKbnllYdh5urXA0U82UbSmI882g5NVV3YcU1MuGW5De83uVRH2Hzs9gvTHjLC7dm9
Q/g9VGedB0LK5NgpN26sZoz0c9mAPYIvekfSPX8BFik+2K7bjDTCQtB5S7neuYe8gqmww6GaF4Hy
FM5Hv0FKb1pV2M8KexkFJ2jJ36aoCz+dEs546aWxGYZsnjZeNuquoed4oYQwp6HycNLC2aQmomd6
QOJHdtYAJ0DbZfm+bn68M14qYh7AFUUX5S2LS9MwbRCX6GiiFr8bL5e3d0MQXyNQHwQvA9ft9dMG
og3ncMqzrOWrpqm2VFd04XM9r1x07EKXClmUeGN+fPbSkUS/LVVIqbcO4x9+XV3X3ggaa0HIjZ1C
5kBXNK0AqjWShHixomo3LBpSQNNwKdVvwOSzb405h2USCbjbjI+ufe7HzNLOtEXQ3O8Z4lQjCRZJ
oPjFPSfgXJqRXfD89dqLtIR7bY+zCtdnjVF3UgIez0LyKSGgp6VR6+8ELjR3FCfGVrOejSbTG/6L
aOuC4lAMSarxr0VQRuinf+I5gyJ3S+swarfAxAYLT8frGJg22V7MKvu/B/bzkaEsIdrqM4Xm7o48
BeKFHUbHK43gp2wruT4+0KOOfotDJyKIK3Y5Ltk/B7LqrynKnw7iRQz3XOzlDhhD/1S/M3GIzxPC
+JSIQ7bP/O519tWLZXFh5B5lPRBRmLj7beSt5nZO8BWtwuLZ5WIJijEmPuAvgbrD01avSXfng3ut
l58zXjoGlwAEiCu8rwco8dci4mUFBuNK9VPoxQvF9aGjvrWqnTnbAFh0/zipQ64b/YSIZSB97rsI
oFagCdCTdCkUCrftHjUHe850TCjtodP/kG5J3v+npXaWUIW6DDmenbcNj69coRDtzKqnyPOp8AcI
etaTOl8+aXxTxY5Anw239hD5AwDVKZ9n2rX4Z4KLoThozVC6TfGS8sRFXyWSQhG0jdilLjMazJQj
U0MEP2pQh+FgrJSu54VzVdQ0bDzTqjBg+R2LHbp6HUl7i+w5Ihf7v3XwX3Xh/G4vOJYqalXLUyPE
KgCmExbRVIufvNiB7gohfscVdExuxTlrr+SIB9p5/U32R1pRb1JRvLj3svplJDXYoKt4j7UhzsU+
yOO0EKx+QPU8iI6edwwVcvJgUxj1ixqrVGx8+/a7Fed/GxxiYTfE1aytCnBO6k+ZuZbxA3/llffA
KdONrIkuURXCx23cRyX94T6ZsK2v8uksF7vban7kyBF4FkYH7s5vVkZRlWi80jh0MTqnmIMX38j3
S8eSUDhvrPzznGaW8GMHHOrsf6t7joyNNxDpOjfKTnPVPEpzqZNHLpTVq+nDEIJMsibfOWaOyJz6
anXYdQl4p4219Oo6VfnkqZF763twj75wtlTwWa2SlbSMNTYd9XEFCmo+P+Z6cdoFy/cytbVVSIPO
IGgSp1SljQ8w/+2Vjp3lIjY9zB+LuKFTMBXUDmo6fAbRyIu+UFEz4I0AMrA5iVW2QumCZ1DD0baL
ydY0pPWqasTG/XcpTP/JUlMUaw9r7XuxOrgWE1T7K87+mJ1KKB8U0US+XJAILD+pXNfFCD3Q8Xfg
Qx+2cstBxDMF56lcVruQSTvxjUSkN6QqwyUuwOuoNY37YFORqzj6mpFt2GuYg8sPo0tOukGOf7NT
Ujp0BnjVsXHVZcQk281c9nGQLVb2GHCtv1xt9hZ9S3i3TS05d0hHJhDYyrsHRfua3U9z5s9RG1Ws
qScC7acQF8Zjqcwb+OVY1uN95RI1smhc9xsbbvkCIJGjzL5OM+fN2v6ZU0WTFNCqVbgzO1nA9P75
eiJPZRTGgqcOiZvTm/bVDQ5KfHRo2Nui0LqC6/Bsc4K5x9cOdJIjcDjPETsXPuqt8LP5f17aji/r
aBZv0ZiieSv+yxdNUkJksGP7WGSeM2QzAKGo/VTqqRP0Kt4+Ma+u/v8l0aRElmi9YaZzRhwYdgoc
S6yYpYXfMSiDEtuX1m0douLJz7+6nFJVQLIMpGWnfsmDetNPkiGTyHaLPdKmtQKAqrLKe/ocNsU5
q7GZEVmSziXrTsRFNTEHWs9v1BTGGWKHIZ8Y0IoIIHprZoahVvVJZ42cjI/YabrMW2DS3xZiAknX
Qe2nWtXyweEEFzTvmtVEazNFznadNJMD7+v1pfvOxAQESrXO/sh8ghdCNeg2HtOiKhj35ozlFniD
DKS20Rf0XegrvE57kfk3yvYdNhsql2yq7KqK5OcHWILumyDYodxtT04WzIMtEAwKkPa89SsnIsv6
nlbevt2wpoFSSTcEgDMUJuRJw01J7G+k5VTPAMDsd8UrBzm+SRS9NcTQY2DFUzwqeR60XwXkRvAq
MOmMw8AsN/55UYzB9e3bHoaya5ok+xBn8RZKyeUGP8ZleFQDf5FCF/zaQ69HW11ThpEh9jqP6/gi
5ib7G9lTPq6JGPVOtP4H++Iez5ezCW3h8JVSl93cTNrkh9PodZWftYXIkhUoDbwFchrsE0D7+9c8
OJoYsTKXX8qA704aafDrQ1QkGxdvL4jb5psQmlLxPHQbU+tp8Q0AezIonPYNlYsF87043/ikGdD7
NwuB8WN9xaDhTkQ5DxJNiEigD9yj3QA5bOL0/yIHt57neQ13MBq9KKLLB1yre+GbTkPGgMwZwnoH
4Jj6d9ZnOwgjZ3rwMIUxqfu34WZP6zN367UUBuT9bkFYvtQL4Di0cxZvPk0vntAnKH54etu1I70q
YxHPI4F67QVyA+eM4BuDdF21nMvKX6InC42d1EqihFGFjH3I6kshopf9jaB62kupf5QMQPpJTJ+w
v/pONH+4DZo7ZYOyu8JCeA0XqHzqLoXCjH0mGeJReFQav9XdaFQpJM3muTEYp/M9xH2pgZ3L/fQI
IrJcZ92U6HMgIeUaYM4O/Gh7mo7hoic7p0+mQCHmxjsikDtgr57SvJTZZnRPpG4nkuoK1l5DYlqt
NreYBD5/dcBGyOBpESdUnJzwD+CLB/FuouTaeH/iHn4WbgUmuaxlQltNkOVGQiMft7hrNXruHFme
/xpojlhGgMNucEhb0inB1NJ9tmG04C/ZyvSCPDZKlAAFi530z9sDRQNSROyL2O6tRK+o7g6YHb5T
vRPO8QXAyRtd9+W8JNxxHXgPt2rnolylWmJ4Zt03Hsczb0A0WwBf3v+2m9sVHvXzrMycUliG9/kP
QtO0RgZw2+GDP2ljyHVDC2nSa/xueV45b7WunWww/RyPUrZOQ9vTMmklGRFzm408BPUAI2M13PsR
HP8yFvlMhalqQ0Cjpm/LDeGQdo8UplSlhCKb0+RdIEtcA/Gt2Ek9/OCoSPbP0506H6kw2mSayGvm
CpUAAFjks+Og+IJxFz9C3VD9bFagJwE1lK7A9Y2Ozn22qxBHHlKGhs882ljzIPIwh5xEVMNamK5l
+9f6UvlCqNY0d8i7VdGrYfJ4SXLeU4fNSw0nyowLi6Ip5Bp7k1rlxCFePORy458eFdeDP4GE2LrZ
h1MG88PIbyn7rs/jqvKphis4vGrLy+YqrcONbprDLHnaSYw9NeKy8arvOlHpUGKJ7npmKfRaWJNm
a8h1VMgO2dvXSO3RRXnNftP90IE+toJIb3NTCYtJ8PycO1A5yB/EHTtdEIkYz15syfUqaWOp/xBa
Qndpt8rXjrN+GFQA74cJiMWyiE/INXG/38HA8mhT6awAzx3m3egR/yhpdIPaZ8HIYYe7kqvxVntt
6wbb6nIgJyR1MFfnXkaQRs8f5F7GVHELxlo0BL8hqNr1c5g0S/4IatWV5ZUolcbTx7Ed27ctiM36
Bkq4p2TEJlmnkcvQsnhvi1DCCjPSqlcy7YXqzTcQ/YKjdCeUPDh9vQGXdQ+/RqKpixq2LQqm8xol
qx9Bt8RuoZPtgJR5r9ugKWs+hSHIRCizOis5LAA1MJsvgNcVbssSRYZ17oP2uJUx9W7+FHOzScl0
k/5Yn/rjY3oKK23uUQ6+xugG4V4pYt+E6fZ0X1V4ckqqE9rQ5Abc4gSEeJOCUrC6YgdoGK8ORo/B
+MX/u4hOHIc86ZZXa8HOglodLwbjdxsfB68wLkWko5Fsv2+U2kZpy72lprN1SBM5u1APbzrlD4TE
4ttBwYEywDij8YLLpY4lWzMq927CFzMgI8h3PxC85bq4LP0EbwVmOLCce4enk5WXcbqFj3Z6Aifj
FHL5DHlVm+GKv/6FJUHcM3jD7n3TfndMXtXcKv9moiVJwa5kV0VN0X1uxEcHQMalO4XNe2kz5Vr6
8y1IcsJHofrOW2SMZfzi8axbQucIVnHtsFDAC4XtUbtg9MWxtFIdlJDvPAbHpCHqb9Tb47wCSik0
gJhEhz0hpWgeiB97OjiJ4qzEvszk5ZiEtzvZavCpX1NQFhoPyiSF1vagWxZUXPgzAvkTb2C64mJs
XNrOyVPL88nXcvkCiQ7p3uhzkvzUqc/czvbqOLHbj/ttZ7KsxgkyY8a+mRZVrfpNrKdyX4tnu+Z9
m/k5nUYPqFt9pZ7Ig64QDMEwe/wa4bf6EwHfmqYejvR8mu/46hdzlCAOSi4f/Q6rfIWehnLVDWLt
SOOdlp/Mc7US2XmABrIwmpJb50fV8RuzkAhYQLtKI5Z6qh0v+MM+lmOUxSAM/sOjBvstTFl7B7SE
hkiYwuz0V71VZ+gTQc0N1pA4JwfD9lsWuDAHnfoQoycSJ6scT+PEWset9u3rx9jDz8daIAiuggwY
u35VglUh774YUq1pY/1+GMDwv199+2XS3PHiNuXm/LB+yZtgoxPTe1TlVUjkv9O3A9C29RQBK4vo
r7flWI2MW9B5PWWre9/VUeTm3RNFjHMNJcqmxgVHYgS2Q/B/2NvYpD4ekDHIg2rZ5XsFFjsNvPvv
wp7oYXSCNMU8mwf1QPj3BonYymg6adBQ3/ncUnSlxTJBZTTJIWg03eIgntMdmUDJpFlZT5oOmsbV
KUd1seC569xFgmAY86WO3cT9sWkqHpzNQxfc4jyIT57woeQswGkW5pPaxECIfyzRfIOfLhByMifB
H8Z+weQ4lX/ryk+86f9uloUZk86r61fQ1TezYJiEjho+iV+cqBZqrWpJxtXHkopad2iSLC79od4C
ZsBex0tsBHnnsYBJmeiUrmlw2EjaYxd1jX1dbi3353+2H3aZ/y23QqPcIFPukesij813qJmhahx6
iv/fyzONqEyWTc0bkWEvqXNNPERGMpDweNGrKFH8LXNr8T99hBoy57h20GoQ2Hf3QbFUH0kh7rkZ
xYYziyh6YLzVPFv0ZgjzY15ig0vkNNYi8cZKhg1D3P4SOWbKPTbsOBnLaiF1FocuZcG8v2YTcEFf
xsF9SAxA+m6+xv/NlWmajK/32Izqvm7rpYx64vbSpPoUCs3Syiglzf/bBP3uZdB0SZAnyxgo/EGb
791JsKD4GW0mYrs+yO5pTM02XrDccaChWMJ5Ty8PDQdJamExFDzYXtMYeJliXjK8fSnMB5NHnJeq
JIxiZCB9u98ldaJoX+d/Ic/qPGEi0VfpBp1YG6L7BU2s3dhBNRiPUB7EuhJXJ6v9UqdZ+LvCw8nc
oWZx5D4LTVUOBGR7G7qBCcoYi5cW8iT3pbpDAE29nToJh85RzH8+Usum8AJc2dYaMxGBMPMOS4JF
m2kXmGPkbUYOhziG+msMGMKBGpgP/gL1tUQ7axAzrhPMYEenX7Mm63xLgC8cbiVfdN8Qz3F4bcnF
O7sC6Uj6nyztng51C+al50hXT+g7xBszpmOoaVXkNxDhWguYZrEE3lYXaL5ZvM1o5FQGUiVyqtrx
mAfvQ0AA9fJKgDsiclM2OG1Y4tJ0t0prNtKMJB913t97jefW7Xh7aOPkAaDoO0FGfjm2ux16BPBB
ezMuerAH5+pm4Aqijv72nFscye2wVm6WxuYtqFcwBLxeWRWr5llrT3wMtNptzEttO7/dOXiGfknr
+8ec5izsOZF65r6D6nz5WtLOS4QF7Guw7fsu9Mci9fCEIDqesjCNoivAj4K1D6hAgUYAa3cRijTL
Q8/+KEx5OYWgnCvg7d4CoqR+aMGB9cOzNMAf4dzASfntZYwLq683hkJH061Vq3oTXX6Zc7FEY7qZ
/wf+14EzRNqqQCwDvxChGVtp35jxAz9SSHpCWnaeJnHqkO5zUDhawHi82VgP8LcJaF0C0qUe30rK
6jPdzDGHEorWqf38NDxUuWorrA1xz+bBqQLdaFzKLG3qOmeZaEUZZ9TEU+FltarzfKNSbpNIQ+Eh
6krTmVMj46LB2qdMFCRvjFAz7sWs/wRqZKrZTnh+csbt1uDoTrokZxegFxzoK2MmUS5SkfIzGAH9
Rb3m2LVlDShM9Iunn7schxfoYpCNRh1zom31qTBUXmf2hpUYd3N+jwxbvnuM/eH0gHm1Qom0urIV
MdcTyVhSe+V5XAI4n9TU7pMaod2E9/7etx8vFvqcJ+9pJExFiUwOBdZ1p2e+vWt/1WwqnB8L6XfN
MamEJfYrJ6VjkMQ2smAkfK1LQvHdP11kPCe2jKmlxIMj5nJVRu0Ayt0ktx2Z0tH98SWc19o6kQPU
MIgGHA6peXcjMoBZQSgy/8+Jf+Z0bytwmaB5deMZYVfgwYsBo0D03LR7zAK0CwDC1ZSDHPfPamjo
YfGJEiU8WnnweyKNfaV7YSE0QSWkKViXOQ5y3GBY1X8dYUibZHXUykEzFck838AF/S7J/tBWpmS3
bA63JcuxJ6uD2CAdMQO6o598pdguCshgzzWskT03JrBcOtHd7aKt6dLOne7bD0KTa9b0kbkGO5aq
l0ibec13vgjwZ+12Z3thMmsnWMdkk1L4SRy0KPIDUDJKv4vwg5La3CAjE7Kn0ALo1FTQoeYNV8LS
toNsVUNZVTZlaSfEbDCRYRmbEEenp1R/w1QmfzgSqS+8g3cIFkrArdEP9OyBUamdA4qoNPbfVTKm
u42Tdwyta1M+ZinmgptKsXSjcSk5zU8gl1MS2eIA4W+M4JQ+ffTpNForoyCNjIiOHE3A/v5fyXJF
WGLk9V8pxRJ3UcjCJOeOGhf7maeXMkliFKFQY6/nux7JpLW7R6vqB3dTh0vW7GimlDfOmTptQYdp
d6Czf14EQXVYYeW7mmsbhVfC7MUchkN7GOtnYNWzuyTbJvI3JMX4eVw7ZZWOpcfpPcTTjllqt9Lg
LWw5FDRYLIzvfAbXzUyK7KbA60JNTzDpguGRlsUDt2LzGQx9aNVfpBH8xsPXUzZv1/MAoQxtc6Z4
2RI1I5Ifga7eLZIBtdlrM+gZylXHzphPrG3P605otYB4Es+7kIli0c67JW61vDrE/tUIi1duH+/H
cfFQldj8FlYbzsz0zTeGJx6UwkzgoJ00IAHB777vg178Pu0lX7UnLTBx6BXCs39yNnJ1HMtpCYZ7
Hw0H27+uGXOm8LKSReDBZScwlcKzWYgHw/JZNM+LG+xJgvPq5rCerNGDwfnBvYal+KpODVl67iOg
xnyPoDEwvhJP4KkvXLX26l9SGBl5jTVsqzTMEwYLjWjD354sRsE8E0ycgZ6rlNZba+5NU5SgukWd
8dy4I6PH/1ge4C5EKvYQsJxOlgZlRnm7YNgMavugMx0A6R3RhFy+GFdYi8Kl2MLK2+hzYITtaEBK
XXX+QoIIvYcb77uFYAW/WBLhYS71U/2KWChnTJrZLFbMEN+UOr3bv//BD2e0Hf8hOMXemxRZEtTj
bOgCW3joveCvQcDC4mLU6h7fyIGiuU4KHmdxqtGtddglgETQp2ohgkJxfHWLDRcfYBghrNcdIRyy
Yh+vsJE8bbaRozbVqYpDbuiaEZ2tNTAjuckVCX0ncAW/yeprrgmheifuvj7xeq7okOJqMh2WgtzN
SfvpN7N+bgxP5NE9gHqf6yaPSlV7MvOIBKjp/CVMj3u3i8KDWgOMuBoRC5Z+HHPhLC4ufe4Wde0s
v21LS4sYZvMxRNK8jH6zAhNPkB/HmYb1/MPZdXfF51cFjQyIE+dCydsCEP4qjB08sPDlpyKU/FCl
uE96J3B9fHtzpO/zVVQZks508DUxHP5k7k81gEfkwekpnkJUSyv8YRmhH/cZqzddDAkvnxXL0wZ2
DZ045se/+mpNyhHYQRlDG2Pr5mx3T2PjCI5kb5VcjIRfCwk5DART4rPb0tylDAfUwQdcJZb+Bte2
KE+B3Au0c7xciT3grU5ro1F+Kl0KkjM6TBIqmPI+GKgCp5xZSY5rAUyAZotG8CnDInijYKbAC7+M
JBQNXb260XklWHHnngVn4BxYBIYOcBA2QG1XYfLN5K7U75mBcEqxsL/oeZbRXzRExvNFvEkDvQA1
G76LLbLnPUPA1Hem3H8EVZwCxI1uMJHvs6nQkaK61pqXp80ttgNCnihUSXuZdN4fnQRMoQumbi4A
YK6n7eL9DZIscAl4R+FTpWF9gvreZ1/GC9qCf7EY4IMCWOb6StqHydyxaN4nZSvuDIQeAiUA3TIU
0J+OaJeS8Mi3wdNjSXe4RQ7QUtdARnQ5wA0grxl/zHsy5j/W8HA1gi7f/w+iIbl7Q1XeqeAVv+GD
PVlFBesFW7xTkv1NYUAaEsGfvCs1I7E9jGhuz0yU3pzqfMC1V62HYiqbG4v1eK84Lj3dZIArDWmo
p1PyDAa1xTFRWVulluuas30seBS/nw0qB0VsCtP7I3tXyo9ogNkYf0xBlGDWaWF/VSVXQX2+Z/01
vCS/nGziZF+CAFlCSHg2logBxjvLICyuojUduL6wo+/miMhU4RvQmv9foO88qe1niIGcmdb+rqii
EeU/Ustgc7mfjhd0i6+GOWQ8ImGSwdiyA8L2Z4fWrVRcCvifLZQAc35pXSgfSQyBi5rBsOwPBfiV
SOiK1CauY1HP06/b/xaDJ8LRG7Cf3spl1dts/KWaFr3a3wAZl+Bn0CFlzqggxUQrGuKsmGZEvMIf
chyo+QPPrffiS4R25ekTv7AllT832+PfV0cKT7kma755tkRrLSNVDPVABqKs0abg6980hzFNGaZm
7/4o1xR8pc1p53aNIhYrdcpCW+qerxaminpOIhQlajUkkB9BR9WscP8mmL3mhiwJXyeupqgFysRm
NsoGkNRZsLkxoQzn5cpzm+zsDUEhrTX7m1Rc5o4ozzc3+dhXLM5J29oRRn6y0mzfBO5K3csmLm4a
YjD6iP5HOR9eJVEt6bN/0PwD1Hs2FLRcfJ2+VDhBKC/+oAut+Y8XDR9RuKjggJg/Zx8p690cowAt
PY+zgGOpRe2iMaVQ91TnabBChIFsgzhYMHiidJbD9wGDJnXllx+e1xv2i2/HnXSFaLnwSOcYLR7I
dkLUpoSUH5zjNkM9E1PwqkL6aEUFEI0/yrxlOEAh+Krpy9YJ1yOuebGW0SlYM3GtmPJmtqXMGwDA
QThGA35cRLx81XiMw3wzHthhVQ+NmKtX2t/IVSFJCOQzgqsCbEcbuLsEgLjnkGyn7SF/W9o/oduS
yOuZqlBP8jX4LwWKIi/QRuR0w2jSXRdO0xuXdqBmzGawAR958MOVpMeH1oZjicQfHelR5V2torOS
69hBmYpv3ab0DZXfRJ3ZRaBRIzVKGw5jiufeMoSZLz+fCDL/Ba7NTbkw8UUh4zcAfp4fb+SYNMlQ
wgTQtp9m80+ANhWju81wyLxN5Nfs5rTj1kNj7MddTp9CLJBGq87wSJzneacL42rBHDuBeWWE64Ma
/15Qv/grK9iuli3A0DPw8uK9LLAJQPupOv9vXhn2tsY0MKj2JloSGxTqJ/v5xw2lJpk3LhxvT2X5
nLNO/sNzbhwQK2qwyAtA0K0tljJ1VtM1o/vaZTFswwWHzET/jN7LRFVJA4gwxt1kkiEfO8+IhbIB
UTXukETpM0CVG9OnCr1ipppE7NwmZiauQ2/BR8RyimdKcfTZmd1sdfAnGXUCBjFL7DpjHQagFrfL
41qvP2OYK0671OZYuPO5oJ009v3yh5XGZH5GR0rchRG8ZkAyg2FjpcuCqHgec2NboOUj0j88Ga1t
90DZOgzB00m7GiBB/uAGiksDeNk3Of8zcgIw8gysmtDqINDNCqyTnbia704T2iBi8iv1Y/1wfhmV
q+Qwfu88BO70dlWKfajQKlMJCR/c8lRl03TmDVMuhJNtmbkXruH1W/13gTkGF4JHHWFQ5JQgcy16
iIWMqTn3whcjjJ+41+HnWiv6qiq3Ltb+9ri29y0/ISM2afxXr6xDU6+7qgOe5sEacPV7q+cW9vep
QOSK/SWH+BP8G0+dr7wbV0LBgTBiBEIaXxulQSCSdYUQo9VDKdV4gKqRxKjnr9DcaStV/AieB9dp
uMVc+7QzsU5YZ7XkItyiA1I0SHSMxkJ/AJgoeXYpZwnrX98C8f+Y7zxL0cUTtv31y+rjCdc6lagZ
PvVSlfZoFCxg6ilDFQRX6fSEllyGb/tMWICIyQpuMBtXrpHr++aQ4/yjlU3ZWk0HhhvCUpgj+VFY
vX/AeBt9veXSeXJaHEMHgwrKDUnMRCRdwuQkEYOfNTrtopBtxCGoDcl21HsNqE1JN7QbknOVhfhg
lgdFteInJFwf5Mv+Ff8UL5LkeebbK1ago4XyE6Zy4SUyB58+hgmomeERm8/7U1okZcEvisVPUMHr
RRj0kd0Q8aCdDXIo8BD8qWTfFKwQiOXK0m1k4wTlrvspYT4Zwag2qbbzr2VxomNxVnSVvJZ+dvMD
g8ZAD5gUh2cM27GjR9ZEz/0NX4ylPbKV8j/j4zvG2N3CgeMqdvsa9RjgYK9yRReMdq8gW8IThQGx
kas6bQf2V2RrBDe4L5I++TBB2yX2DoBBJqmiy6O2aD51rw/0RAxfWY3SNOCIIf0nA+8rJp1Bpgoy
EbGgJZw/oIOrgpNBmQBIROoM2jq4c5NgkrJtzjAxVLqHEO8+IFx6LcpD81gETirH4MBU/1RXcMdN
662nqUeaRI4iX9xfrdf/KR5ZCm1uOXEEDcgLK+dBh5uwcvv15Q3Z1h05S4AHhJqKJ6IC7j2voy/f
E67qNxRcF1zmla8Zn+xF/a70NRI5PQWvjDK2CMH/hGSEp8RF72vnPt0MolVD93gYQ/XEzEOwc34/
SbpJ4X3N+6cqunSQ/VhWl3gYdHt5r/+DaxG6enjm/zirxWCqPtvRsMJPnI5/FxckHbvdK8qaASx4
NhtSU4XVMncX4MDPD0pwDShkc1313koLj1UJF8RzQUeGnTDCExZdiJZ5w2o4KDdwNG8jw2BkjdvU
OBq+hSy5GB9/y2d3f+7R6hsFgt8mOzNohKGjDqOqSQFeKDUbVUdu1pN0IsyCGe1CpN63aTyHWldO
ICvcHSmOCGmwq1Q5dzxsK1XsrZiakCq3fv3SAIW/XvbkPpu16N8kFcbGCIRJZNPASxNADKE7DpWT
mEJ/XagApkAAUuUZLN1FlanoruN14lkFiaRVZm7r/U/qtNtnwnNqCDqJkgalLq5xB0qgeb7CbVH0
ZT8K/GBuLWb5KemNQQerSzqhQGW2nX82cidse0p00Ht01yvlDlzk5CO4K8oxcLyklVTb+ifVtnd6
XAA4KMt3AcHNsPnopdfk6QsjiaXn6pDCbockyaKIlayOS+1c8lp+I/7KoPbUDU85ChvqE0+XuWjP
jNCz4ksZLxINHNCrztXPzeLyqYvBWSnKTG9YuwlP5a3Q4Vd43UtdXvD4O2DRB9/yVp38T/17+m1w
3uowdrLXBllokH+s+Cy3dQDcp3R/uKPCMKq9OC4axuBZMGuBc6/zJAgIlbDEk0lu5Wka+fF6pLuA
FMPDrviUFfOsfbzyMNc9BeMZIOrxKAJ28uF9rJqoPhJOm3BB8wkqEQGPJrEhVUB/C6t9NHrsZ3wg
GJlywm4E6nZnMlErxey0P7ZfVbZdwVc9oLWun0vUjRVvNIZ7U2JGEBArlJBIiYOpgxMs3iA/YfsV
dT+YqYqw6jwaAPbFIrkNDSUOJW8V9W7vTEA1L2ksFWY3gxuPBrP6P0YNm/v28Zgje/y+tBAhb4Fl
PX6cf8b2W+hD0l83qbUIH7I3WqYZ0M9O+N6f7W8MEfthT28wvokFyP/w6qu3eL2bUmnmoKqXmnYx
Wq86eg9XbnrMFDxmnvTCxwlTdtJo0VlIQGwe3n2GPopgY1XU0Cyhz788/ompb97/VpwbP4+uz+Vr
9MVlP6CcoCA9ChHjHenzAemuVLgjifbuVjQVaRtuOZWOhtqfqYKrzGs6MldnhAXNmK1vFvd9k90z
3fvsiQibJOmtsyxkGq9o2zwpH7MuEjVDGACRn7VP4oroieK6DaN59NmdmyNrBKGNGTYNhwKZPWYk
SuYsoyzZj7pydeM6HmwW6cylr1JIjc6WOa/fsHYs6ebWlONKmAL7Z/OjUqSD6xBHhc4b91owHCn0
OvK1n6DDRA3PWpyFiF/tWouVw86IxCipCPxA4skI8bL2FmJKlhwr0bIHo5JoKFeRPJ+LuFnHF65Y
m2sZz1eNg/byMmIDVjwUDbNf4YoPoCy8W+EDjiV8LQvAyYztNb2g/kwJjKuZEP3UrrWRtpkcAr2C
9oPsZ3kbaGt9W0V6ODRTyOA1IrVVEu1xecr7NGS9oVM7EDGsh12Jxb4UnPVEvqaCQJXPAFg5qcrz
JPNmUbnZi7WH1p0IM4Bc0qFrxxXM45LCMKjdPUlLUE1pwmT/dHXWw/AN2JhFIBEzJjTOkoSEqSv3
wZnhVRyIj3o6Z7hvenskHL4hiE1SG0ZkSImV9qjJ3Ke5XGP3KKaa4fRL9iIC3Yv/YI2AXtT298OT
2apRseoMdzA6RqN7gDpT0xsVM95E4vNQa0AkswTzRLa8JaYXRFUWWEP1tA7tu+NFC7BKLh1ygwgi
GYNg48aiXAvkUTHsOUCrASuR6aE8EZfV941ZTaJnUdhkDWPAZNu97Trq/tyQ2kkHlBoAdcjRH+lD
QYNjmATe4GGRCNwcJ9spRgpbksn+iXw4TOLGdAIdNWFiFpWuU+uXqB/Dr1rrotsUbC2F4i8PPkXz
BzJ+bAoezF77JvLcaSaKwX5ZRboNXfGQ3OXekel7daC7MdTiypz59ef78f6hL8HmOBwpPDZRa2zz
3bjMHTKUpZUxj8s5VLl+9qJVe/XMtfIOG9rqMo6jvw2//ZZ/Ao3PUG03W7vRnOD6BFJndMhT4whK
qO7if6gmHv+7GqUQN9+gpRpWr54HjWmFPc8MTogy22ZoEqg2lkAnyVIngeiUHZ1Tto0jhmT8fQwA
f+rzpEpLGPeSud1DSksDGlztt8mgZ9fgcY0D6tI7iTq+hgPJ0ATv8o+9VUq7f2jNZyvIZ3Rj05fS
5Q350ny3FBz/mIqgnbmcMccm7v2BHIYASmoNwH8FvnlVL8m7bjUo0SWDxFkj9pd5yAFdKk8AFl97
9LXo3C8WwVhydnA0y3vOHJ/d6NnK847PBM7A8te1xYeFFodj66qXXu44N775hLa8wsHrJo6GCK3B
AtvamroyM5sY2zWcbzSWnUvS31lRk/HvQNbWxVi+DF9qrXPKDPIn66SB+Yr6BOP8Bg5MbU9TYxG4
FaU6BS8Ozyr2Avri+oHCtgWi1zr6Miw/P5CxD3ph6VWm/84LraOOtvCpr8KBJ2Zm+H7b8T6nzCcn
6U8QPVoDsIs9RvCiVj4lRv8uHi8/UQjZyRtsWGou5nzk2mHBCEKpofdqNW2gT+jOfyb6YbqWFVyi
9D77NJV82Jr232Mv5G/MGB5aMeHFDYkQRRiUtRUlQb/BZa9HK3jH5k0WBtNTkZB9n/1Sm2UWgW8v
oBeRbWAAglaYCx1VY1s0wRYsRfCJR2sUPBVVpl+aiXX1DW83ZoNV7GDNCqD3MWdMAMWOaaGZA7Gb
MvhyVYVj1DBGM9TjD9ad3eYqGFRAiWSddw5Y9Imu2XT8Hsv9vQRzDhkaPmxJoZ2VRsrKRW2REEd1
PFT4VRbFPSeT928ML/wJp6saHysB7NUWg7wjIPkDd2c2Bwe+ExCqpswKD/wiKn0PZXR/AAHoVm/M
wJQ5YvXCMceHvHQhq5Ng8/iZ9dnsgVLiFoPpGb0Kwt0oOVtBPx3SOjq4ooSJE9A2caNvr2dhEJFj
qZbnYyTbR3iVqlZdZEJOVghQgBVtY3omR0CMhHTmkdGGNUVJx6UyznAS1KW0kmkirQJRnhlhCCKq
GIgi4YrvKXy17qxjpg7kP7Y4YAHXe/8x2Du2KsKtFpUSQxRaxzgn9N99yrUU+35180RHncPG5GGx
L3ObX+4RcUfVT2/Mldy/8EvI+rM5/giZjg6pavpcNVkqy8W+mxdTpONzHY3ia0O9DpXUo9c7611K
LK523ybPRGuOCbCl6d8iCdIr2kMabA32PhY6kaKxFABZMb0lHZw1myklNT2jyyXfThv1vNPCLc/O
BH8LnkRUd39sNgIjYkTI1BOeCTpsh3OWIwvyk9cUw3pGjUZS3/wrLQrH9xQ8VM1N0q+ZSPM7gs98
FcLBE2Aelj6TufCZz8iSdMviMjbkcOiIpN+eecFVtIo1LKSbeuk+SsAXvTO6KBAuWkz0dbDtYMU3
oa02cU7iKjBcVG2r89wh7/ljzqAjCGoEH2FjXKNZTJefTcL6aGA1nolriGJoM7tqqntbVO8qaR5O
25o2U4duBBDpnMkIdCN7JgO3ENDPIvSOvhf1zjmnDwjZjsGzO1XWC2UHSpbaIl+t7cPPpNcdSb9e
3WWPXuexR8OpfCihpIKCXOdczY4lUjuQDPcSu+VW+ZTLmXpbwoNcLzaR6PYCkSy6q4hotY4nydTs
LE9C49rhazYMrx1D1crnS4zSGqrWQpi5eFWGiXslYC6jqFrt8dYpVxMSh5UD+0+3X/gT8dzaN8Ul
UQr3nt8XN4AkrHYP2sQ+8VKbdsqEhShWMlVafQQIJ+UXY5AVyFphOu3Z9bNn74BBnQ7sk+uxGEO4
saTQjr/C39mBTGXQpzTZRqf6cbpC35V/3/Qrg+Sd7SxqMefZbhut+6XWh35yhlYnFURdiRZ2vWeQ
T9Btn/LH6110rWElzay+Ot5U4jZsn9WjcMpBWf638ROTC63oSuXMHLZG2ewGwLZgF/4+QDmwk0bM
Jxm1C+ahYqos2Qr4EkXBQY8XEDsWrGCg8FkAI+qKObolJTMUbGdXuiGMBvlpAFH/cYE8C9kg/9MB
TgzVCKpEh0xofEEo+i4EXmAw3UG53WdYDWkBZ5yUKqxjwQpBqKnZU2vSBy2OvgbmO7ipuiOtwq0W
SlnRmjlg8RqGZK7LmPhqshyIkv7HHfqIVKftn0bNzBWeDg+qZa1IdPIPUJ7B7cZO+5jWkUDhUkp1
fg8ZyMWhFDY/QGr0HRUvouk2EAkV3ThV1Gwq4n1q+9tm0avhvxjsyLoc8xeCIIR9Xw/3zr2u8FMJ
T8pD0og5EJf0wkmFOEM/KQXLXuxunwObE3PV0nHMRi/vxcCmoYRr3lN9agiVCaIJlvyPPvqWrUxh
aCgtEZooOFdPgnhwOOHhmvqp+5VHwkoA2b3+TvQLb6qc9VnTtzqkMEutnMQv3AcF4LWCq4MCEh5c
iu4Ezbfi0NkNRh4fs2GVUaRLMwQYSG3g7l3nwdHxzaQoXwH/z2kiJeNuJH145H3Bm7pIP7EE4epT
oNliAl4bvg5woJq7+JQjpxgemOdtKoKyzGy9wyz+GXyyoi0nCFoJhrL3ILjUdVZXJWP+s4wNIfle
RfUrvMMxwJRZQBuhpKPlRAOaft/h7w4+8mJ/2izLV0OJifabMmpT/sIsJbJLFLSOZw0M8zlDYk5L
yxxLIbnq3As6pO/YqRz09HjVHe19n7Fn9/2O1d6rm0WeBNHaFVzU965ti2zD/oJGoy1jdgP546Xu
tSguhiQIl0T12rmXTyqv2fN5t34oA7uLc0XPKH2YCpLjS/l6XeCV6MP+RJuXSqsVGStwON7d12zs
zhNmMNvBiC4Tu9s84DU/6DbSD0HllVb1pq+UBzBxP0GOC/xnfvyLC3CZdipZ0uYo344IHfSvssT8
JtYn/li268GpqtQlvhZBUFpAmjKjgKHJOt09lqLj8ZlBqvfuyiOLOaX/x8fo0Eg6G9OdVAFPc0I0
CwiPmDlocxLZF5T8X3LlqvJssKoZM6cdPvfAJ6fi+zqcHIWTQt9LDQrfI0+UsSPXf/Zu/ut6j1q7
um8Xr6nbLtOU3NMTNuQyrOvW4GGFo5K9EGz5clExr7zGHmPsZyNWyqRbJArculu+d7Uv9WW8Xk5m
Bt1Jv4JyvMLzk/c4+DXRfiwYTjrs2iIUfpQ63lq9ii5fvOxqu9GTCWwwuTOoDiFT6uxs6uJToXGs
6flkMiEHuN5P/TElQZn1M1ndz4AqYKhmvAbdJf+xd8IRK4NVAUp6bnLqlfccrYAYKZBep3KgkYLg
ea2zAsskHR4FAwKz2MFiMYqRsiGnveF/hTUUwqXJeEnMhSJeayYrmtkVjG0hascQR0S5ZcXVFpUN
eyw0AvvoZZZkrqqq+kiaY3/iM9lFZSOvwVnGjzEOVwOzZliQ3oZ+xFBgalv2S85+Trtm1otnN3QV
OwqC4wNBbfFCQh7vNkvMrCXjDeWAI0CRmD5AvMYsTQiNiB2/1zU5bej5PUhHJJpqjQJz6JmO3b+N
FgRz/6MckF3va/uLnlR8KAwwbGJHPFPQGGOpVA6ceVnSHMT7ybXyse2Wrw8X+WzOCauI+FAcM8L1
pSRwzLsENn0u9ZRuY6rimB/N4bmg1gNxy3r4zvr1+9gL966abL4MCNtH4YX/kj5c1Eb1tC0WcFRp
Dn+v7XP6voxzrAA+2DBdvAgahhTcHv31ECstvpqBGttHVhoxM4HasOCG/uBX4n1Xo2gzaXY/00KU
6ESxfwv8/tYERjlqEJBppckcI3APhX/N02thgO1iNHzPwL241Dv4MG5/uKygdItH5cVEUL0MUq0A
g6stuTx9JwK3QY5G6yvt/0T2rnxA8KabjNF9NceYDAYXU1zuT8636uFPaQpJYY/ochmzWUJIee/t
m2Ou41acF8/vZMljDOmTnyqmp4lh9QKixVmlRvhtqADX1zYMxwi+EPH5xYoPKC4YoIJe0FGQo7s3
P/3+ZgLpA/aWbwbapcYPQMUNysTqtSodFfIPtODtpgPCpvJQOsII+kxfWZrTW4rrDwI3Ax68zRve
wxzJVwfAKyfTDzsHT4NJECnCoXn/yuINilTWMLSav58JRShOz3v8VBbryaTWfWIlKHUQW0V4VYoP
8suq5JGwJ/aGYCJi5udalyrImpzAiJdqV5jvV8nhTLABsQQp23WVlzerKst5SB5PsBKgygFBdCZy
MRaLxPTTvgQy4XclFjDrpdYk9Hyy5RnzkaSpRJhKUn/DaLq3vdttNx1LUG756UJEyz6VOVYcvCjx
9YuLj2GF/m8StktGdEDwkFgUBXt0ZWyTzW20xaBHEey7MjxgnFptNrcgVc3SDBIP4O9qk5LyMnfy
YtuJcqTgnTvlW4LgQz2nIywPV2hXRxMIw4TZaaB8f7l1ylBm3TJenzYPy7Go2tZS1aiubL2Uaaou
cDAekDj8WiEe+oksMQXUGANSYv9KI/6RPdUi/260JIkFdk+xlr+yMjABo/skZqRIlibW3c0dRx5g
s33JyKCT1O18MOKUSgQlHan+/kqsoG7FgngYO8KUoZvD/6wYXDOFF5jJzxA1iOSQ6sX64ysY3Pc1
6Cal1R8AaMiuv9logoKBUCqlC78/l6MlYSRuRzulWoDicEtMk5NKmqbuFj53Ar94b2JSdxhQyhVA
ndpEeq5eAbGKsvyNd8Zy9HfqUb4BCILMzSQbDI97vOBxaNvJNlyfrCSABlxYEaIM8YC6JtF4P0Zx
tPhJEW7qkQIl1tJvu2cDSFtJs0AmBnRD+XdNmzcydMaIHMzs85UtQBv6fE+FFh3o28uWC+arW8lP
EEN8oIkJHS8+WWgyJD/Zpsj2rl4LsacOZxdSRmvk9BqAzThqrbzdTmlhhiL/lBc+OvQOgEhOss2j
lqpmIYbNDuEmVQThMgDC6Ep/mWqEaVK1xzpxSdkHLj8AHA3mZf+cEol+ZSIfN3NAKQDs73GvlaOv
4ylfuyUyrgrMetEZCmqJfuGoi8l0vulCQb0iwsFtN3Xi1oJ568dBcVQb6Oa2/aJHpVgaXt6/6Ptp
OS55tMq+/svX1t/j+3kczcYYOfaZOLhZxRZpJB5CPlR39gLBMXwBQOiTPw7FAWdwAzRJ8tw8Xw+F
Z6fLHuYb1fXDXwzTOlObGhvzN5xK9nSCcFSzntTjKD+SNA/VVT2K2sFsY3mR2dXZB6d4Scse36P+
afbsazuw1OkvQqT6qGAQ6W6sm9AlqBEccqXS4g3DJym72XSgfCcYsGcPC+LLHWAg9LIJYx/6Bbhu
0gxLjewveE9X0LiIRtC1MGmuaq5YljQKDBR0zsndBdO4+zfzarQEtShPUs+Pv7RwpIPo35tq77gz
32VXD7Q8EA0pkd7FTGVqbph9/+/opHxSf+Ceht6TsMnN41UzPklg2qrcU4ck8G+4u9anzFXz1Q9Y
0m8sfim+AW6Mexy1hkJKnofh7Pia7hEQ9qWLgXUv4U/Us1Dv/U5GA/OhKtJr1ypW+YuRYBbvNXMi
59E6CI109N3dqDxqVxDbIP3uoOU21oyB6+HygWGY999MOkhmfkuV+tXgA7hFFhbyZfwLuOh6mG6G
l26D0zYv42g04joN40ED2uA287GK7taXRzGfTgBaZae8akVyvePhXLoYx9HrqMC0S99Deg8DFRa2
rl7FK0Fk/uNKN+XpqnHItw5zlH3FDwDPupgVAgdWoJRmC6Z4R/5HPjnHCothzWB3O9XEl1PxZiF8
LFzi0V3fr/lwEw631GmQ/xlOemAMx7k0xZOm5ckaxmJm9BVPyKy18cKckg3bKAHELYIMbGhYSaGA
sVmgflQatmwGVgM0tTT6BvQ/BwSJhTrVivhEPnZ38+4vqiJO5Hyc/jP1mADRqr4mOIMgxH6Nk3Ir
V5qS5Y42qjp/az7VLts7llm8YEDqGPioo0HL8J1fP2qz6bD8rXUVDacxKYikUc3yLuLiwPhWPfyA
/DU+CUnez8JrXcufGhSKhEqNUPEv6dAfRubGB9H+Hsd6WZHLX8nrI65F9Mjec2Y4gh8zRvhm9KF2
wxYBvtA5n0pS4PuCPEtMApH4ftZIOHd504uuvSUpIRpMfFCF/Whg7GQqZgslZD1mYwwenj/fEblR
ViFb+1C9Ykpm+nDZTrmNULRu7XTJaXmvUL6MgRCj4UgLJXbcrmgaD5BO+3xJKEziv0mNRF/2yX+b
Xxaary8Mjbh2Fy+5s5AZr6W546kZXN03Fa6ykGdG35+Tn1AaNXBCvXpAVlA8/HZ13iV6ehMIjDMf
I8jx4NluIr0anqu3OUmZZUmipFPuDw5lJwXE0o1VBdBXVybCinQL/RgysXPP4cZFIbyg8UKSrjhk
7MyAEId1mSCem6sZ7/OjZTamt4uhsOZZKWF1s5JJwrCmzWJSok+PGePc3IMNy182h3GIMKdj8tUJ
JuZepnrlMbkRankkRc+C1T8wmudegxzhTw5PP+3wRdSVxp5pjPZT9osyn4FZa4NFDPCFkVgnEEGn
rZjP72qfTs9QG3eCISxWa8t99Hqvzu4QFkHl2mfnfFwus6aaJTOFevMb9NcZ48U6oMl6Yslp7gre
eB4VIZl4jnGxVlz0N9SWhE2QRaCviH2qyoiYlhtx83G5IenBNdf4pMceEQD8RNG554MclvuLMnfB
Ri+By7NNtIRCPycgp8uU8uthV0MsWgA0tz2DQxXyZdXRS4z0jn99rWZI93kV0tT4QtfYZgn5a5/U
339zJME0wYH7UrIDIZtH+qLhtPE6KHktfJHtbpLDiTeW5Hi44n7q+1G26mIEuoM+O2UnriX+7Fus
xwqKh/DiF04X4FDeg5fD/Jnn3bXPlXVOBdSzNeET3jVV83ofsFUEAq/vtx5QAAieM9RIcncFTm7F
N2g2TBXSe/zb0O9UQRliYnJVWbHM+W0ZqHg0sJEWFbUlmaDixjt0AD5YZxqQquPNwjRwU/77OM62
yTehzrU38ZZcQStHzBXcCHnowEvCnPAsjv9zCwOFB7YSrKgS+av8sMCTEOMZTbQZx2n5f7zYj4/E
NH94fehGAQw5ZKLOs5O6OPXxpevTnmhLzVX51vHcQoWXqUBmMmCGPWeL498pP52b1XaZWXvZDwOc
76ZdWhPck/kbMCXKJSTHJEBhWpHZL7x4jvppdPIHUD87JL0YYjIx4/stcp5hnWOKu37rXvLrKhiK
5QU92KsHA7ofP/RIlJtHjZi/EsrvsKS7TjA1mMl64c3vpG/NxCDS0UXNp7KH1wQZA5yfkOyzY7WR
cY0Ix6bbLdXWFxDYvty1WdrOQvlJcUBmfX9YZbtDTQxv0Mzebbc7W0hnZaOdbGVgbJcoqlXST/fj
vQKYvUsK0sDX6EZCfxsKwZcJSe1/wUxXw8/2mIK7JR3AOy5UcRAs+YZX3gS0d/PXEbuCJRC6+nYy
GRXQ/vxlwq8/pmJIUAHPmWgw7YbPanyx2wA+um7dmBPzMGeihLp1cfOZO9ztQZpJt8+DxBAisLdQ
XkLZndtaBUAZT4ggQJ6LJWRSDucT950qYsqGX9/7aeNq5lSzYSC3BLBQrJ7kbSKJu9wg5eaLLKrd
S+CImZMqOgSt3Z3jathVhta1Uy1OAD8jeqyjLWI7l8ENmUe0LO+CDPV6tujT9M9hICpQHsBFhaci
5TG/4/F8x7wgra95z8dmiU23Q6jGOCtSUek+zyYwaQ2QbQO/1LagUSkw86KwunQGw6O98HHU2ZyU
7nJrPazt3dd2CgfmX4GkVLSvDuZIwk8QD+j77WEeW6PhvSYipoOQd319JV/uGY7AdN3Cd77KUIqe
4TcTMAsDmjhbZWt6ZEKcRUfvsBnGSKMMDUnS70n3r/s+PoKrkpS5IYoKKSScVkqg8ENhjiY3mv73
pqW3x2ZBUNb1PnQlWzyZRcLf39AqijQS9iGNM0ztTGrFDnHWdr0nXkP1QnfPCPSpZlW8mVVjDsAb
0ewRYEFKLaF4uxaF3+YG1VZnC4uYqkIhFJLACMMVM9jyk6OO5/4DEUEHHdDe0ix7Z46mOKK7QcLO
tpDY0a+I7c8BBkhspXe3M8CqwegPFyqgtcx14hZ6UQ4Wctkf0Ebl4eldYpjVeSBuC4zL1sg3kHhe
L9yK2psGkijW/c56GeGyHuVyrcK/BeUeCtgiIC68Lye0eK9eWK6FXxKfnO60D5U3MCpClK8+5lU/
HhT09Tmmp/PePtBnQwyxXWVUUNN2l3Bw26VFyTyFMKsPTSy9jcNzXcTqIA1QbgLG0niuvAN1XgeW
TGANW3+0X84jnVaQWxfr8Fb6vGCquGDCSL9nbPrYmJpA7sZ2BVS5UQIquSup3X64LJMAKuPtUK+6
jqatYaT6UfzYrVz7UD3lTFSULlPF6p3j8pNHwGWcQsXf4kA29wGxSfrI0dhOp4ROxomd94li8AJC
WSQoIlPFLbUK3J55n5f4TMy2E8NGL653yyO6U9Jq+ZdjNO8Tt28eTka2zoh/QttGd3b79mO/6x+M
e+KkGHMzzueJTWYmx9VLkYGRs1mWElRhRiI4pc4j4mdBBFdRaLfGDKjoZVFz95BUwAZbZYyRivn1
TVz4K28Psh/Prw+/nym+zV79ImSwYNT4hddKAevW6roYAkbaDKJKLtoNzkPPFYpmEj/0z2f/NVqk
nyFLW32Q7xvpWys8G6AnGOhFvpAXe2EFHk26uiLixdfyRcDsOFChQXImujyWiFF7m45zpvq/R2gD
l9W4P0Hp2ChpAayrUKXkMVudppo3p+29XOf/OG1jkO8yrbZdDhe2x7uPGq+tXPC/pp7uRBkDUc0K
BAMYON9oaPhdTqMIuyWMxAYfsrPn9ulFPqKCMT9BobDOKN6NPgEVKsHTifPXTQGACtV6nuMmG4Jw
uAX34QY1hMTGexYXRlcDPeHNcf1tgMd2VAkm4RFCCsmOSGuhDGzeFEBtS48ec6AkK6coX8njWt8j
5Is3mBs1lw5f3wd8bYf1pfjcvEdrcbam+NfztIAnsZd/NBF0AV1RZPAc+75OETm1LPD3j0Lxt6LY
T4suEC8piFfplqasF9/ARpQ4TlUKA78Jkn8eD4ChuupRA+bVxLxTFS4cdILfj3wcn78tyh8VIYdr
fNPezJ8+VEtEPwoPSXpsBVhayB2DaN5nZnel5LTFt3JKGJ33vUevNhJFvz16x6CENYbBoBp0KZkv
wlGxSgvShJeloyRu6izx+oXWZAiCz8D99Nab3yYq0/rKy64748qErKYe48psfzinWwKkOr39uFQs
6kX9LfpFkQvWSkTTRhT4DJwBVrz+5WC9YxpEI8pudv53Y0RcMNMqdz0rLe0631KymBbF7tUNMRzV
ToKUCNibdBfMerZ/ACfHuvtH3ccBRDJM/Aq5yLW/K6zx8BXoowzHqJveRz7Tg3pVdP7k1cwzwWE5
AJJFZBw4n5V/pGVY4vz8ldrCMpaXqj4s5Lhinw9WUR6ieFh/EXNv7k3WbOaZdKQZY8ig54SN1RYo
CospXVtsPdGtMCCB+4Mqb2bNUqec8uvPGRaIWeROcg7iZsFPO7yde4f+5Otm0flV1lrd0W6LD2KP
2yMY2SOsDFvVjM+jJI1hrUzLbAaINt1HKf/cZrYLZYsXdG8wFzxijqC1J0EhomOhqRY71ek4yhf3
DSueIfVB9eyRHZtS4zGTFn/eEel1nBWdULMjXCKaFy1JsHHGzTIFHpyBt6qQ+dYjmh8Lz68J0AAK
CWPGxUDNPGu+2znYoBhaaunPSQ0lP3ZBCF56pkMtmYJ6FhsBYvCnnCyqC6WRYx3uvp77hUxNZiL5
2oZdA13JKsqdhsZ4Go9qNlrL4RaDM4mPr9JcgD7mQlRdB1GPJ4rpSufK8+Fheb/DOaz4g8duL0tu
QPJRHndgGKN7whz/ViJkT3EC/iDPJYrb8CYW2AMofMTH16Bn/zcXo+SR2BVnMu+2Ft1OdY8UrBOC
RKfDrZ0UoF3pDfQlDx2Kb2Ac8MkCM09QJqnalxIYhLqJTlblxgWkRWtSvkaQj5j/diFox5uvBpK6
SugRkLKTbkwzDWdsHYCAL5HHy7cZ14gdtN1mQOWyCzQeky9n//B666rCFniaiMdh57r8WNuhMdLi
kAHbFKtDRGVOsB+kTK/d5XrJVAc2OzGg/dizW16JmWsA6DfTvJNo8aCPQPVT6DVl1mg0hTVNFbSl
WIreFjNIXuTYSHduT2PShyhQ/Pb7sC0JDCYIYenoQgbpnkwCretaxhZltiL/SclHYDN/Xo2/wirD
+8OoIzMP2+5aq3oWIka4IbYnL4qC4YgLX1S5Cvy63g8tm+NdG/jq29+k9S7VlaXtN9hH1GBBv7rf
P2q6+GVXgK+RrV0wivBxBqfbTLHAQlB7C/sB9R6Dv55IQIagqgg2Dkp9lyBDVSOh9VJp6pOUQqow
r9Ix0BjJ86mWbWS5ckoJDjCjhpqG+o09LkMuG90vPErL3zFSckeQxqwWUC013bI4AzxZlMHHWcKz
43aeaa0TDB13MskiP0ZPNtY6zyiDuXWFoHvaUQvCC0zEMkc8cMKg0LcCRIELR4T2bs7+LrvZdvSB
cauopMEInFa2G2G/Pxe5hNA1vdqSkL/XsfWeunuekeGoOed2hp2tejcGzNpmMbGUlSMkIK+yy46F
naW6gKzBLjSJvOo+hV6ZvLlGcIpuAkKGo2rM3HI28zknRoL3WnSZ4cxUoTJr5oEZb1ajQYia3skz
tIL+uO+8koa+mRaHIUTWoBtgytUtZGnwF/K2vyzYxmpCBdcIcD9xKLbom/YkuIRb+Zm1wYkcTL0O
4tSbKuVpR6WjAAdbQm4tzVpp7OBS69TvYZxah+q2Ng+PrAeRf60GXhKTNK9TBiApcL35wZw53Js8
vK5ZBWrw+qFBm4cqpUAUL2kfakcJBExJnNLrjuOMJvaKw5Lh0jQBtM/JVcjf+ldTClxHQZB3cB8L
noAsGI100g1SnJ3CUR/8iR3R3M1qpK1998c0IzEU4TOO5b6/dyOqVuMzO5oIU45Hr5SvEHx8iZtR
Yts7/JtX61zpW1HiohRxZvgUj/siJNeQ9JemOimixtZWKQQICDEQwOwWC9qaf/V63kkkiwv0goG5
yvrF2SnljasNIhWwUhcXPYqfC9OqDgRVydU+jllZGl3g5X4W/DN1Xp1KeuMaHfNrLaI1u3ufRqTu
BVijB+jVtKMHLxUGshwTMOSh2TlLEPTH+9u0vgboN37MnQS7NuZQCRmfombn0IsIF4DnKcNciu00
lqAaUngYAFyNg4fc+8CxXryA56myd6GU+v4eh4sdp/3GTOY129amP4YspT8mdp6gkMLDGD+Po4ph
83kWspis7fT7o7DPxnRA7QZzcw8V9Nzptm0NgHdi66WF5r7jkLWbGHi0etOpdokYujR5oeiFjEg/
YzJwBCV2b7BrYaX/AVm163nXkgEYivLfV9xAKtzwGSSa080Z0J9L2DRg63oq6MKp2MpgFMm/6SA+
/a+ntF8R+ym7+Pp1CNnpWt5mXPj8fWpyHn6S88xfrsPBaycTlvirm8VvtnXVWtIh77S5ZIps6Ezs
b2ukmTrbcWPOScKUXI+FjdabPi3Rzl967NXimdb4k/vbskaZF6DUTiXPUa6o9tahCs0SB5XbtLzb
Xnx+mv39cHt9h1eASgKcThXGzgaxO2g4m0oIwfbsFdR2HSzZ8RkkX35eAquBVQ4C23M+rKPotkWe
n3XUEzkgSf+BCCaRUYOYfBrOrZQiWsU5zDVHzdsDR2WclyGCr4MtjvyS69BVTpsN/I6+TkzZNaiw
m+kmnFYgoMsbkooha7bAdsyHw00bk+ZRlQHyl91ZGgm9WASy6q10ERlJQcLrOq/VzZoYTAf6uPr9
Hn68t5QIGLXwYof+nQVwRT4Sv9LOnF00fXhBp+BzCH8IyJ9fphy1++c1BonEKhI+2vyWnE2wLcIi
P/rU5s5OrFc93KyTdumnxk0m9/OCBeJRIvy31Pfl8gSM3o8CVqpYVtSnOQlv7dqqctNg/BnoubMN
ApYWeUiUuVnM7Y27EWzudSO6qq9NqLV2a4/vCB+pPSHuuEChZnKgc8XZdWGBz6nbt2inn+bLXL8Y
pEAkibiFW4AZkaF80cXPXkJRmWiI3nzphTzo04vd4z0j7+bUEwNTZvkMPkJmvSSKDJkvixGYmbEw
jtbUHGW9/AHeHaW8ARq2rpNok5N8qZlGkJ9I6I2iDW9zFHvuNkubeZhCZR2GJE2kI+elOBA1L4Eo
EZHesQkMGuDLKWWp6gUdQjq9LmpAUUE0ZV+m9ZkdN/ACztZl3+sJEC62sCPN1UB6zePg3k1EiXO4
T7dhO7vZxVvDMWAncNx7z9GsQ36XmJpnbZwzUvyORfThWumrwPHOwwo9nkz6zgXaJlsAHr9F61r+
NF6RnN88PyoyNoM2zziQAn2cVjxYOr/n533f+RKGzwwcYLtxvm+liB48SBPcX4jZFJlKtLiARk+O
0gAYDZ98MLeDQNCq5QizwPk7tW4zMfqweNe5mHJa1MVlouxVzLSjmu3a9sEWTKSfXXWyC/AnoHMq
7WVibWnx4CGnABE1pevgFcij0+23tAEIz85LPN53+ld0lqmq4kwf/eu8ishmpUX2X1yEC16/xCZ+
uz6j8x95Mcytkbiw+53QKnSQvYMZ9aDD/ODwO2zjW0Q+qlYbAHpE49YB8FEu+rt0llFqlewFSUpn
kLQsQX5IBi7HKSD+74TA19avNbQgM/2FCeZzwE42j+54rtZvmeU/eQveNCEbeicRlXpEvwZrH8Wj
mnmY8swJ0WxWs+MUhIN8XWaYjvwRWpFWLoZUOZY1JPTgZi7KbMlDtxW1WjlnX0OcjEvzXXBgW9M0
GkHI+A081e77P7il3m4RhIJdCM7BnmHDBJW5Y53LMefmKQF39cc2Pp8fCA95hoNEx2xw/j0H+ZiK
c4PoPxO+sJGIfMSNM4oFFKeztx0h/nDctJXkrMNbdZAOCI1wDFl6F3ABEQzWw7fKZI1kO1pl4dH8
FllBS+17492yAvXhOwbGspEqYtqsWFehrLq8kQo3LbkekBL8SNUvXPqgO3oRXArd23ia4SiKEz7q
orL5UpWvIKxO0cYwpcV8tRDErdEikwSOAy4kcilH+PtYPqJNqece1fyYg3Zw+uJ96szIhUHRl5vr
uMC9IaIwg/3jU2jAyzE1DBqrivaOs4hti0fblua6VA0YjgSt+Pe4FdlFOl8jKwwzlZ+BW4Xl4CXb
JY55p7fxFSGI+31i21BPI8dpv0WQFdzT39yG+3gInQNYnVlXy3a3U4mnMTWLZiYT7vl9+FkmzWJo
T5X67xBkXGYudcZYoqCAtcApy/naMbYeA8GOyN2NtadcLqiAlo0RSTTTgXRiITzozBC7bHx2OqF5
qza6078ckiOEEIMByENX3wnUYgqdCy49c8dmEozsGf/ZHQ91yAfTS29DZgnCLFR1a6TgxAWHK1q8
ANr2yrI6CmkuNpfGj344j8tkcPibn4mQvKqNsGj1ngCmMCKUTMXz0YQDjdYLxVM+z+lBEtZAA1Zp
4DqdjWb7j/uyUQBbDtc+zMbrcumBvTMF1pO7/ZunRdXhROtpl+/+xynwa/HRvZ0B1JNLuksCX4ci
LKTqzQYe79S+Ty1+01+hmuUK0sgi/hlU5P9PAb4jgqwrD5qBUQe2GG1E0tnf/M7ngBlOvSa67J+H
gIIwVZ+SvnNbYigb9BnRoQ762dRpSKBxgxc1vk0sQB2PLHUzSTGqYBUji+Rc5np/7nR7Pm9QY/r0
LoPVi2HgtAXsrD/UnoUln/j7aZu8L6SZpGRUCWpLgMxI3ntM2NO5YjwIsDNMJCxvxShR8a/h3XSh
IEuwxzKbe2Njgk/NOOZ9yQ69uFo3kcq3Lir5XAzlKagvQWsyww5OxN/WHIOLiuQoMpA3LaD2anlT
e7my4cRquyHNPN5F3qifCowM6ow3baRT19vU4+yI0KTW8scN6uiUimefVlyG75Eqc4VnfQRm0j/b
hYUPT5bs+XP/UGGRtNEXMC23rmYzP0Xe0Ai5C/KJEw7IQ/reRt+cOp43KuTKHFRwxQFn02PeGSvw
QdFEajW1ZzzKf1H5BgKs6esB6Tx38fQgvsjkZPxGhqXfFco3IHCKJtZRMpO5Xq5WAhe4v4+qL7Kv
4vy0cvVDw9uNmXwMb5pLCzGcRfExhi37A/SOr3GScNULyicoObxQXtoap1MVgizVm9D3iWiVv/6z
Osk5qYoyC7ZAHMvZ+sWhVUJLN5DWfpym+UrKQutBlw8asrj6c1e/z654mmWBq0Q64s0JZ2ncMDhD
0FKdOzBJfUfOSNIZlRc4DmcqkALqigg0tgU5x/Mu7hh60PR9bLATj1xZI1lqhFJ4Rm0KN5WpR/20
Ztzp/Fi2F6GQ/UmHvQz4kd55gcyB0LPwD/ZglorLRb6rzx72C6IbYPh4xtgb7Xqe0NItQ1T+fH1O
jf5L4O2hjxaIN7p4vFoG0C6yOwCAbyf4gretx+LU2KLz03uVVSASXSN3MXlfWsa3gLMDp5MYYfes
xBFaB+z4QVqkVwg/dxGSG0ajvLIGSleXPwRVIkuJPrWA+fokBd43B4FGL/quoFTaMGAk8FU0j73U
Kbd1zFkK/ezdELVmPV6QKvhiWYE+QKRsyZ7GkDliwNnavuX29rB7vbASZwD2dnWYIsj4xRoFRzzc
C0j9+8uuYX9WpC0tga8cWIDH8VKrjWuUC5N954/TDIoomxQPcf0rvUr+AF1+c6z0/ZIesUn4tsh8
7mLuc/emFuDNKWCLsANlD6sPh967TnRkDcWGcTo9sih7NIEvRtnkAhiH2Ea1Q/k+scRA4NcNEV0o
IpKjSpIX5Mj94ZhzlcAYZRmPi/a+trgQ0Lqbkd9sqjW9Pb7EmhTNlxSyEHe3M4w6YUDBuEYrT7EQ
+LRzcvQ0FTJ8oeJyfQss1UqWEnskaiyqXVMy0HkQyY6ZJyKkCx8EyaWUp9pygpucNWgsb6jt8fn6
zens7Gzofnm3YxitOf+n6giXUZv97cpioQOxFlFX/D1tH4p9VgbG/tUVABaswV0fkqHjTeXvpy6Q
PDFaWcAbozlSDDRY/VlB8X3wDLnGISYZUTZNVmEeSSm56cN4h3T5ssNz+o8UkXv1YlmtFX8Olnjs
LtxgaQAsx/Iuy+stjlpJ4H+ZgZi5fG1lhYaVQYebjE8EoRs0W/9rZJhuuibUL11jy5YV+ql1GOwL
mALXZm8Awwea8lo1/6cSJX082QptH8E3TMu4TtrF0AwWMP4abDUK0SCYeZzhrxB/tKOFE9+01Q4S
c2rx4mFRQC/kjSc1i13CEgcNWlyNePiIgODEkKtnhyNQb5+kigovDqErljQXmK8cJB2RU4sBSXr3
KYsH2Q9JCjIwtJ+q1HeunkLGW+37Qrjb2tfIjNaokB0EvnuCzP8Xuu/DrfI5N6h1zBFI98GqbMHd
nQGz+tR4OhoyhW2veOnW/dZau/pwMEzrsNvEMiYX/QZH/UaKYrW5W3KRnDSX4ZOdhKCpda5C7SKm
i3W0obSL6w+NwGKBV9AfLE/O+IjM8OtYI+ng0Nlwxe2+y1A3Q4VmbLGNrlYgATiwVw8nVl1ehS93
SK3mtotAZYYTypqOuH4fC45kKzyTv+pJoMPukDRVTB/QrlT7LlbcTeuncSKhCAVvyibTeleR1c89
CXEovBp8EE0hpbvPmDl/QXsAZeNfV5FTVpM6nvwsOZBPrZs58HHROUL3B9FHw2oYulnh8nt++wg3
+4ufM4yuSNMbe8SbBxsGqVznQcx/K8E2JG5jAec484JVG8hdcPgPVLAbded7UsiPsvyHhUcVdQNW
SFKrarjgz86IxuIzhFGbz7OZ7DP62GlpDAJhWwjHfHUEh1e+N3zh5Z0xf80xbaVcxG8eVrz6bAxZ
d3CZkrtFwIySaghof3XSWNSD/YNvhdBu49P61nPU+MQ6WPST0UksZsIsUyXmdk/9ur3foWAD5XE4
WevHS/rVXylXgym09gLx7z0azK7p+zbPEWztXW76cxgZExYCl7t7mgHtaYnSkhQK0YHs6zzpN1iT
6ukqHgxD3EAdhFPakFOraUbcu4n2ym5UPsXumMVciAUHhu0cy6B6BKscgmxLOW9RHNFMKNuYCbR5
mKXNp8UeI0f2AbGoo6mPGh8snFvrjlCw1NzcgcFGLv31N/vV72xgo6k04plE5a25mtBb5ZuRQuzB
v9+K7TbT2LmC7+MgjUJiU+Y65MejF+GTr5AeDEsefB3f+YWvVT0d39ev+X0Sk7rWPblHnSJ1/DZi
I7qCg8QNcS5+v1EOdJrx2tBEo0rI0nfVcgGrGDYgzeh2PDihXQLZulZKhtmdf2iG6FYggWtB9Nuu
QA6/D34CbwZ0/qK1MDu9Zm4vSJO6IdVPi3nWST6v7O8Zn6g9VmyUTuazxtgX/E8xq4Rjs3/1AV64
1awTKZRX3R73o+Z0ETZoS4xlnnSZB1lFL+47zILvKF3/OGZ1PWgtv+tp8h9P/py2/UOvFuWnVM3B
hi+FrMgq3zXjyahWA3iHM1gZTnN7nF0EIIPL92s0ToqiSwylMqrVxv9NniHLnMrMvRZcV/hH2XrL
4dO6CDxCX1lnAn2IejeT0iVrShMiM8LBqt16SlPxO+3JHGtcD3Ggx6Ao6FAj72yXD5mrhZKT6oyV
wApbWL9Brkkeev+B9SnBFjHEKgU+O/Zg+FIryVt1SiLPnv9W/2vBzwoev+icvIGsz0R3wCMtgszA
8E8TFBhUfM8abcf2pcR4weCujwFR2I9FacP5mDcpFWUG+morFurjIsEY1ZxnD0FEz9se+owMjgmG
5aK/NHJcIUm+3Hjb5dqHkoKaokKJm+wHa+O/8oIv4/pTjUZ4vF/WH7PfZ42Rq9BAoZ3OmTGaWnbC
2wdVgwvWe8Q3RDcQsfKcxIMz9vQbxkQTXec0M2ayftivrpnkw8MajPtDh/54ia9SSVlxBcbm7/CX
IHFxh4R2B7/jkYSco+z/mqDiyhM51G4NDDDYA9xwgtod1nU+tBpqp5AO++5BpLZrAujM9CaoLpLF
TpWiJKj0x0chy7z08cWJBoOt1pHv5GxEq/iCG51/pNClga6s0s+M9G+MKEYujKnKjyGjZnrdZTPB
mdZowLbqxH5KG7NGbH7jo9dgEi3uzqi7UXJ/LTLJHoPhiNFBgMFxK0pbqzveBdNhRYUoeHlOVVpB
vCc0pKtIguiDoi5bvzeYenODw7CWV9rPj7+S1sKD8i/tCzZwtbAvSae2EDv1OAMyp2Uc+TsLsvZ8
y+iieHSJJ6ooxktaIqFQg55PSZFsXpArA8I6ALktj04B9afJaPjbpwlx934/mh7k/mxHZyqORRlI
SIk6cHzYp9Sg3TIUNAAQnpIG487ohjrSbgYGPnpQBgPxpiInLRHJ1f3IdC0EMi8tGoRTiGPOM873
Qo5gAv92LASUai6m7WJcdHhXrT+Olh0/36lM4iVJkMDl5r3sBZLGCXkBu4Ymcb8QqdpHWBtYXy6k
qXzF89iHUPSN9ctpS8RuMUXxvoa3PJY7w0toKBqaQjgbacXq+ntMLkqnLyAD+LYhrO3Un/KjBJDD
OV5kmISMWOklH9G6BIwX39RWo3/U0Z7d50iM85HNaSy814M4Vw1DVuRfcnhBSEqPZlHGvHI/cvdb
hdokAODaWBemZfLDBB6jK8f7760oHdG0vUfmaB/ICVXWb+Mi+zjmpzMZAXmvy+baAvbAkud3CNkD
IK+fzmJkUIGx48dcnIEe2elEbEpJnta1ey46kiQzMEPS7G/WjndthHMoT6nAYhgfE6WpnmR99PmL
exl/+WFr243D0m8cVUMdDtaNL3zE3DBPp35ON9mFsEfcSBHrAaHAQuGGADmeEeMmZ8rhkHraplSv
hSidMohtwK8qRxA3bu3nvzvIoA6pJEeZedd5pXdmFiuQkBUx1udPPHyD6pY4z8UGVFnblrFwWUWA
IiU8S7xOjlOHcJRH/YcGpXPizsVIaqA08lOhAtTP1HvAGIlLzhKUbG9goq9HDn2uklW+WXGI44uQ
LSPV+uviBP79KlAittg+DK40DFVlfEqA7eLWn86yo5958uWZaaNgCwG2hgrSEYLwVt9Ds3AhOYmx
yPCiUbXYRXohosrAzEoBfk1A6GP+j1X0doopy9vunKRA6Iv0NOAIptRjKqTCqLzGmW+WUx8WWBEK
vUB79nlw98BdBGoANnIqVEu3wjSyKJiSMUxULKW1COlRdusOSn5S5IDFyFPi9FJHVmFyPT9g3zlP
NudC/pmKCQYop/QwEDa3z+kCJsvXeyOKAjimMpyxZaZ73KNkxkKTVtvZtemp/nvIQPw7JcSLhdDC
sZgDiemLLnq9bELheoAhXvN2i+JSMhcFNXtpJx7w6ps8SPwURI4vi0heHn6JchqmQyGttOIaPI8G
c8l3eps27KZ7XnUmVjlCQYkEyEs6dCqTaa8XofHWOpLcKsPVpXZ46eaeTHIUSW03cJMgFxXL78gx
MxBlZWl3RDwSJCet2qStv0F9foUumcW7wrCkiZgHu4kLfUsfpZ05MT6Zw98XuHP6tEQY66xj/+7I
67xDcNUo0nZnRXFBIkTgK6uLPW8HTTOTLNi8vu4QyXKfvZZpWckCs/Xrd1Nf6k4Vy8KBh5OaOmfO
GtE0Y+pm3jLmZwaPOeDN7ymOB0w0yNPR9OcGRsBdg+RoDjXVoe0Ryvl2fC1z7H5NSZDEEMrPKPX/
DLbxlz0MZZApWcRGmnzYWNdhsae7EWuKGf8FnQDYVolExvxI7QfQxvV+Kn5JDHAfd2xExtWwn0xa
Ejh0rziDVSM4/vWWmQU9wiRGgfwPvLYDAN01Srb+CP6UbS/HOJLbPTY9ZCBpuWQfEw2FBg2kU3ly
djejD3p0r/+greyk52aPBjws9uq/Fu62q8Yu0Toxjc3UbYfd1794sxv1Q0eGrfOQ19QKJ1/UVpMl
pXVtsfyHjH/zE6qbqnd3eXqp3gHd1WuJyJqxtTXTrCoz1saRRCBnjltukvhNXQ/PY2U4sqI+t/en
TBuSWHL/cWpDjSDX614AwGx2XfGhZ4ovh0+81N4baNkfhX47QotltQXYNFVzWdFgTJQirYdMx9b2
bQmTeg9ienLxUdJyXZ5Wi7X4mmf/gLuN4jiXjhLbeq4OQOmIHr5IqrVBFu1gdN/hr4djBW23z4N5
IAwiU3KQGDpr7a9qG7W04eX087WqnhFv6GbV9v9Tv15azcdMegTSom+vTdD60y4yp207EaFVSGTG
OJcqH+R/LNER2JgpPahZEH3PGtuuHqoAiZu1x7tue3A3Sbe/cOycaKsmEQ1eDXrg0X7MDx1zZqt1
LG3hZGh2Dbf/x/xVvdZUJj1LPltTPxBR1lW1aIvRul1vSHiccM2nL1/LvMCA9gLQ5uZ/k0pkCOYr
C/fvAd1tyFnARIVK3LclFbqejnhfIGd+sM5d/+0VP1r5XV55woqVN/+NIs6sNL3QypQQEbdouZbA
BaSjaqkVc+T2EAKQXWE8wQPu46JIj1I3hKMOOnmIVE9q0iM8GuUXVuj6cuCmz5ZzkvDLI19j+aF+
eTYrHOOdEfwj2Hca8N24Plrl1BYV7QXOg0OZAdl+Hg2QahujfYlC4UCervV/Bh7Vcjw3ayv4OOGU
HVugr9WxYjbHCI+LubPj9fUEXnMPXris4dreQs0xuNkhUIKOXSzWevo0qyn/frpfEFTCa9zFCJA1
5kWU2CG/x0ftkJT4z8zdroFqruGL8gI7HGPMElxDLdSG5FPxodmUOWwNUEwDShNPExNyL4n2d5LU
3wWxI5I+zFVk1V5pvdnCd5KHBBbCapBgjB9ODjd0A4r149kOz3lURkVTRrRwLvQew9OmEKCkLp6c
h0sOmc4AEeC9SJKVldOInK5VSfYhp//1V0jj9BFff2pfscr1JoC6wJN6Rr5cQF8Tq8FdQmY/w/ym
PUBLUyZ15ma+XhopLBxvgGQKW07ofxkgSaQShyDfXUCSySgAa3ca/d/ga1mMWgo7Pa5RopmNP0Mp
tvcLyk/2HWm8I0yTbiMgEs19MTrpAWNjE0sv5EmzA77Uad9185Je+N11pyq03vc9Dq52z/ICamyB
YaAld6uPb+T/tDdVs6wBh15/eDZ9Eky9+PkbggXnp48TrhOtL0Ox4K0S5YE1iTe/GdPUx+Q4Nhw2
81n4i3qo8O1iSHPoDtOR+GCBiwfxPaPx2RzUoT+IPARlqKmeamCRjziCKSIKBEBSoPUHceNZr+ZW
P9QA8M9h13PMVMu46E6N9BU8V8Bx/VgGoYkSmOdtzITUsB3vJcXx0YgxnWF9vph1nhB5HO88PWQj
wCIPHF2d2czgxGpNazC0Ij9wkwkHDG7FIB3ey12HM1WoC3tRcr4WXdJJlmuGOcAw7c4jsFk5+AL5
ZJCWQKZHsDvQnNV4rEqrPSVLT8LP4nHxcHeUvdsJBCY8Jk0jlAQCvDfAh8/TkFEgNkbPeahWdDMM
RQHBqmazXZEgmpKij86cVEGlHBnmPnIbbYe7ASc1Eb6bSY9k89hHCV7MXpm2n6+2idgcffnDXg5q
sOa49EKqk6D6na28NU5bHv0Y5GlnRmb+j4sd/4Y2PVJlggUOCJsingSie7Yi3wktNqX9jEqfJRJ0
9rfViY8lEkmCS2R2LnrAh7SZepQMOO+dNNRPJKCHHmJxwzt7WqW3lOy0rzr+3xtOP6idgnBR9IYk
yha2ggerGmhbZjpAgIoneDXMY0vSBk1FLVulQYOMpVO7CD+94v10i7/1tjREkD5x4lRL2O9n2Lny
6gjKS7LrFKOIL1t9XOSNIOty1ww2PNhDdYxY3xvlP/u5KhGnv4r5ThN3+NV++5OUOB9AdVDTl4dJ
jFmyplrBKMPztvVp696yezKx9RRolCD06B5z2inrHfT8sqMi0JBAGToYOWGH4TBN7YqWZK11kAqW
5DGRl5+ClwTAy+EPjUZeXs0pgaT1bmXvk2MneNLBEYqIIIH8pGn9kQgVU3Xs8+jg5WM4efLbuZ4K
MwHXVTOFgUw75de4j7E18/MxhLTCEO0XGudXi6LJVNZ/NmBZQyf+221CNfjMJMOtTydBqBclLKTA
XhVTrIRyVrzQoEW+6lVRsorJNJOOsJzqHWu+RTitlDJRTQI8k7HNLtgoTTJztJDnNlsM24pkXwYp
GvwApaxUAyRSL4XOSrH4qqtE3AXySY1KEKl59uqGTToUPgdbEtihQuTmPwXZsZfUP7o7wjAVpwIH
/f9Po1M9aHxT7gYFiT6zZQdjJKRWvEdGh7/sbkcjKLOSmvCAXZMJVSMlcdjSsLFRtC5D/eaSh5eI
kSHS8eCat8EfPqug6Gxz6WNe505V6nydMr6QilMf6Cc8UHoZIPDVIqTkiSPgHXG0gFPws9V1hQ89
EZJWeUtLNoBpvys9sm/4bp6cfp7mzxaSRfzoB0YdjHMj2m0lZWl1EFpSXXeh/wkkyTPG7/YvPM05
x7k9KmtvQssdXd3KyNWGqMwriA5chBTVCEM6J1wa6OFxcl/HCE24sTqPKmSUDzvN4VuneYHspi+S
JI1zfMPta4U0fObx5mWBF8B5/8LhVm2z8ivJnQqWz1X7vZg2faCxssqthdPTKxOFcqFTkycWqRKd
vOsnaeIV/r6UNfIGXX5YW4KKc35PA9yPvLg3b2QEWBPDAAzxNCeff2UW2sHGE+h/c0kBXnAG1uJm
dsxpFQpZbXD4sd9xznYWo7n1YxlyuPidJWRJ0mItUzqFu13qefet0/qie9CkncIKm0dccK1tXMc2
JbwzOX2ZgEcmGenzF/ToZ12qRS5eSr2ufWyOHaze++GQPxSS/YEAWgNceIt9LPUHgQ17YOcGs8cE
d7JoHPPxYo887euR2kVKhOH2hwShU0kucWI6hWSFUSUAAGssBg+xJgSH3UohjTF50qogql65174u
ZS8Unh3WKXUE06e9j7Oly7gHjonzfdcSNtBtGNuWxFVVriSLBOpWLacTLMvaGDxqYv8CBMaqP48Q
vzCT3Jha0z1ZS+lrU7tGqi+TiRKe5JTcIXGeIuE0EyYg7QWwLM10hOs/p2V8DdgWnEyZMdoyN1XK
2twCG4XeTcoEJ+ALgkAl+fKYCSp7QCwK2nTZCGQD1pgBBnfleSNbOw7Q/pX1gCSeNjBMW44Sa97l
QmAV9497X3BM+YEkTq/Q0PHGJLF7wapWfN+ZLM4/qwA9i7PcYIi58dHlepAr8SEIBzheP6NOu2Cb
tHbS89E/2NQsepzUN38N/orh8r8AsPNWnFA3QKCl40RQM4JvqPEF84K7G+VgfMlzIJJbEA7u+Hqk
NsYAGHnk1FM1yNgIeh5JZGusrn67E9Xy5FLSWAh08Cs4IeyU2ZbTeXhacuZOm7w73psuWAPNar3D
30x0ukLomVfYQUeXQ/Cp/xDyHAqgoojlvCzF3GdBGjCziAv41683f9OIAHgEXuBMGcHhKe/B72cM
M6YmeFDdQPr10QyoqF8xnGVkQFS98Lnj/uCMO5KDrD1EXFctb4yTfjNEgjkp2+UF1YjTqBBw52wI
avqqz7zm7SoGAT5TWs53gvg+3uvK2ClrILWRdHy5sz1G3Wew0j6LeFXmbtdPTX2HfQxeTw5k18Cg
yoSc2GI2BWaup57RTKirmcpkUQdhmqtDk+W7r3mdlgZL6jHlz5Dd1VfFG9sEtfNQqgb3ceaaj62A
hSRO7cAhBxQLKkdUCi/YYx4Evq4iYZaXR2kfmBVumi4RGjrVPVBow2889c83lGQOPvigi1q+ELiA
BEdOeeqaMdf8gFXzT4t8ij8u+pgTCdPyFhYnNoz5nVrgvh7EdEKs044ZtF4fxjFUgLqMv7K4xkQC
e3L+BQA2hSWCS4OWwkZRRS+j8+sJZswKSa6KqlakAhXqgFDieca6XpLKu2yRxoMPKX4/u7TP+7Bv
3Nn3O7Xpx8io2ZCRZFLqllCiNI3w2KD2PubBdEjUwUAcchvQ9Te4QmuHi1kcE3qvmc67UjgRcpG3
UUOxR6jEakGNAI7VRjPQpfcBhMjdoSpabE7stfvdmH/1smgm7jjbfKSYHXKdj+vSV5EhwdZETNFN
rNQawd3OvEJWvFryU34P993Zcq8qDjN9/6OEzG89pLPfLmSrT6KotVc8YHLamdCcdI66FOSRROZF
m6iR6ZSdGbeh5r+RzFhBubRbfn0FNfCMcHVPPCPednKpU51JY1kL59HFQLe9Pv01VOTCtQZbdtkR
KmEmC2/6aOhJ/LuuqEFTOonPsNvFsygxhYMR9xeAJD/g593zRy7U7CTqB0WDdbyUT9L9VfqETSuF
XkPGAbJxZy8pX3tNWVLgr9edoPSJZ9kUp2ilI/QM+8XQIuLvxgA2Xg4pIyJ7yC1VttAUNjiWtxoA
jH2fZrq9+mnJrFOZ72d0UdnuSmS/4PAj0149KtO+883xGArEaOYXnW9FMuVtmJz6i1KTPqqOnKk3
rXmKygI5Hle3gGNYnYUg9PR5nxo+ohvEYnXR2tRiH6B9Iz78nyAePJEsAK7gD687Nywkxn4nf36C
4VEyPh0/wYRfUH2JhWPRxWMvsR5Ky0iInhkhFsVbe570n8JCLUlRWIBzaDw0V7pYab2GMdCqKNZN
Ui7UjcPEjsso7pWJbxjYMNHe73xRoBAGrHA7ZJTwSB7ptypCkF8Za8w/ebI5xPhIupuM+FXhiybg
Q2We1CDvjsKUwLRQ99UTy2xhoDJ/zaF5RQHW18KXtr7X6N87qm9WyoLzxdxy9gUqg7wF7EEeizmm
BBOWa0qg20fbpXE1P9bs7vdt2d2Uu+2hytpij0d2pmI/EUtG+un585DIrKuUfytthUWjVwA2vbcY
XlmTuAts1TWgPQ2pPBEEt0zBhTGbcJcPusQ7a4pfPPBlB/RYknmax15IRpYFugQdu0v+4NRwMBoY
PJ96xEllhFOyJQT3zboSXi4K6627H3Q/0qV9m7WVETNs3Kx5oouEHvsJNlO6rftW4UNIC5O/OB//
vpM30ChYRYKzq4RSO7+G4YRZCkoGhyn6HxE1LMuekF+px1SwmP/cOMiriDE0osW6mxR37WuRLL7y
pa93+dPEeOo4E2vcU6ytmNWB2s3Dqr2WWO7ziIFpVnigdbClKyQJemq737RHuLdBUivl5zD6u1QZ
ElLTivZCTEoANIVoanRCaMWlIJDZ1g2STAAqjqhyckyMRvTk4wFwWUw5XIKcZL7hLzTpojop6QmX
y478bfYo3Fmctviq0HkE4Vj6z+VZ9Zz5rfkAoMXaX1KAnCshOMWIMFjltcaXtWWstmQmJH/8xUP4
h6j5Z2I82WiCKBWOsXsmw2quP/3vQer4aSlY1C724ZCrFoxAEbFvaOCJLmNJC2ZuTMTW2JV8eQ1f
9Xi/BRSkKRoCJ9Q8XUGgdZgQTzNae0dcVidWsK3fdlSz1CFijaX9gHNm3fQKKV+j/q485R6bhsUT
vCKuSTVUdkH+FuLUmF9I2ZeXCpuYmfTClfqlU3TZMUOGDTdes4fOHqzDa1w0+slkNVXxOw39qeUJ
FQ1WcO/EDdyoiVrbCL9ihVXYFGKR/v+R6bRakcOive6tW6oeXnZpvQDze0rpKA2b3ah6cwxBWNDB
0U98XSJOI/mLNFZ2JD2eCS+WB7yPxaIbl0ct6kSSvzgT7IHPc41d/oI5YVJsCdPZOj0HAPaovMXy
hgew3N9Iv1Dxi02rinAqk6KC3P7zsZNxftNuo6MB21z1sullzZEX7xEz10Q73zQqz/3YqIAz3Y3k
/79m+NiVVhD6JZTMPTI+b107xqmm0dwBcbQBRpi8WY1tmXGy8m2bExEZwHsZoXkXbV6K8i5QK2/k
eeQYmDt1WWEtK+5xpEoFvBtoiHYf+ZmDHLNomCtT+nkO4y8FgCzp+rGsjRb8uO20TFRUdSFsQxe/
ONifchWRc5lNYEnwg5P4/3+8eU899+5t8NrssvnY28x5nnYduyD88Xa5nXcgmhVq2AegVdLFRAii
3p65UlwsJLWLGt0K5/ZGc3XGww3z2E18tLJDCWbTEXzRaC4jB8sfhaTLA1dUoabWuy536qzynScT
LPPFpThniF9WB33s2QbvXxZluSnHSLZoxk/TraeHPpTOdJ+XjA2pUU/92FFGIE4+oSIy4l75K3b1
nwI6ueRZ6N3sR5+bxiO2AhHH3g1o/Dw774o7VdxqpPpKivXN9205LWEtm1tsEnVWIk3FWmzQ40kG
KXl1TIHQZWpVB5Mi1+Drug98IzqZsNhRlLhG6PgF6gi8sypTwveV5/1iEjm/vzotmDXPx5RxK5dX
N2ddrDGl0H70vHWyCYnFT59B4WK0VGTR5/MFCWerMbuwrZS+5Ri0IxvDat2j3K7Ql0QUJuMRuG8V
vz+o215YYPdOZRndKiMiZFbpsklwUfoOphBlNxviyx4NLT4fduRwOz74UfsdR0/h4DRUk3aoEvKa
AHMToA49PjpFczvXa1RTFC9Bxg3EEYzkMcms8CJJvzC+uKbGuMqaPIDJDvhnjz2IYmPzSBF1FNP0
xrray4nMUuWVGacr50CwsXSLAV+oEaqXK13YAS6t1b7daxbrC+9PPdxgrvaAm9f0W0/d/TmZ3pAU
eqYeQ6dMiSiXxLB16sIfZ5HRQxqReMJEiVG3nUQQWpWymyzTTmS+HiKN4MGGQnE4fo38cdiwsWiq
u6FvPlfKIRQXdMFT8YnOho9RlY9Pt5dms9y+1ZFuu/RL/phUrrWSaXfrUQYRTkZCribKG39rW3zo
a1YRbPxA8aZ7r72upXM3JdYkLmJ4KmtYd3MszQAFRw0afTINqmmgdq2c+AkFH+zLrQs5cGe9GJbW
CtYRo237HkaRLoz9BsjLc4WlLaoWOP4fPks/7HQfKDF8gKbduP+kUjMx1igchWFR3Q3AKV1ouvMQ
83f9Rbpnq75HXfL//+mT/ccecDnGpNwLT667gHxU4Qopboi46faPItx4zp0VqrTe6S71nODbh9bn
8rUH1Vkobx0zSF0ycOvsf4K144XT/jrQR+v7keqi2U+cOrMGMLDwbB6eobdIgc2IL0K7ikSTzPp2
E6A0tlTUmNoAfw8cHK6orubvPStWY/EGJPJKHyNgcRqojyaFWipukc6jwp+1VJYhhKIRXDskQTV0
4CoDQLhCFsPIbxmj0xTc/4dXeSgn5fzxuQZiOhGPzuhXqq5yC+vU73ZVdSc0wFEJb+AfdFJsuLK5
crP8Zm1MMasCy4eavuYOjYtJrqScoVHyR+d2RRtqsp9AoVBaM2dDv/uNJoZiRfGngW7A3y09ZzVh
4fLlaiCPQ6njndW670eyugBR4u/U+ekSwLk3XSdfHLUBcwIBjuaDIHFkjI0OIPfBPFPGUQi78dGB
omCwd5I0m+UFlB/2JO8kpvWDjftYv1pXPiN8pRGwUAxX6h1bPqoMpd99EJTfYkNUuubhsdmun/Xr
yxJ2fjFKQ+j15YOql9agHCLZXG3A58jGwuShh9nAA/IYnC5yv7dyYt2r0UK6qZki3rJtwQ+6LF8Z
Vvj7jcGs+UeojaWnDmmP3B1NOd+oIAlizKwr+fpFNBzr0hCutRNFabREsJoPopEXN9n5xfQzzLD/
4bphwKRIx9s8Cg4l17S2oYRcH5uVtoJFugSNwvaaqat5QbP5Fxcz1vk9F1rim0wuWl8PVmwd8FyG
WZjSlBAtcFb45adeTo8X0nJPQgnFtWGZgxI1IA1PA2vFFfDUfJa4b4VA/dPLPZx0IKph3DC1+2jM
UZZJRR/egZDKVvQ2u9pld9gUB/ySP8Nzfa6Hd/5Ln3F5DZui9vE4JY2XJ6U6mtFUEQZ+gVWmQggK
eRYcDinlxdXItQyfL2sqUHuxx+Dm5DTPUeJbdxWytZZ8ZSudOunaX5LGkkXQs62Sh07YLGj233TT
7O4Oy6wEEfxOChWaUNc7s9/4W//tQJ0MgckLb5ahT6Qgovqc3xO4hONKEJQp7c3cyiI3F3d4UeR5
MCjF8nHsmuy+d+POePrqJbwuF7HTkrmlrbnLQw6j935O5ABi+1x1Wt/Q5CIZmATvdC9s2h5We4D1
u0eZQjwGnQRNOb53FvY3XdWDvXHWUHBDPxUsRHqNRVsg2s/3RpPlR4w7N93qZI49Pe0lw3G9PAGM
emjeMZNN1qDwzdVQdAfvIa6IROL+7ahbLID7iWAiHfaGqad3JBznYY1mCLczFABlaCNnNWf9cZkr
nwibIVoE3lK9YqqZo/LoOQagPj+e/KKMBXwH6T+5V/PoxTa+bgG9UL3iSAu8OQ3RA+2QfloZ7VFV
byVKvE/81pSVm0GnJi8voRy46In1MgrZLfbVQF4sEtCYYf5IMNJHbH5GEOZpVLWLGkuQrOKs9QOw
QjHA20y83NiHxDGVoS4t0Zq3P64F8MtXlMBf3uYlxPyo4HXRTPk9QyzCN3RO8xSxF7HI5wtmaeS2
QLB/SHkGrfmkYogaESXhg/lV4Kfic1ncJ9r9x82h06muCApa0C/tGEyNI8FCgZuBCtHRHbTj2cYH
ULfG+cP4rbXJdgqJ7YDMvaNCBr60jTer1/BdIWH7CSjdyjZWTuQXSG+G3tRicSZuR6fVj7sVTUKV
YvXE7sQL+UNZq2uSL1HmB4aAqY4Mw0PM/3D+4D1niAYHZBz/BW6s27508jYq4v2hsRWAYocYr3Is
LcMxTQo6BFBdXPUeO0qgo5fU+AV8hJvEP7sCUnKsPDQRUk3y7lV5Mk4W+1O1YblSViErrqK8S00C
ZbLihXLMazU1CfS7GspZNkK9LrbKb6ulAiL+iCxRaMHVr1hDfsvIKB9iFVdAyNw4dMX2k2lOI6aB
lMwnbmJ8hDPKIYDsIApoqqTk1EGl4ibhPNk0aIXoRrDNxQJQYf2aVZEzrCJxmtoVdjbduKCT94Ad
TerlNuQ6W2KupyH77MUCAQO+J3YzIs6CxFqCrNN138lqAp1mj7hXooupzqqID9hb0hLXnVCE4f0Y
7VkefUcqsvd0siECWMCMxYPMc1EWMfnKnErQ0ScSuYkujSJZG2hx9SSGMdB0w79lQwC3VIqE1m88
DhrzVoq2Eqlnd4J2hVug8UNM+ceNcN0mNQS0LX3sD4y5cCs9LfM+rASN6HjRt0EJHXG3DkL6QOXX
MIjUzCDGnsSWJRfG8TnEAe+/HsF9bk9mA1lOJRW02Ds3xWBHbj5FNdH2cbjVSbOxBJ16bFbddHkL
SpXARXvv6ek/5PL3CZJSriqR9LZaAOQBLl8Y8TETSFSsEeSI/kQxqUBQ1eHlZRaHaMpJ3Ear2U6g
PoISi1e6jHP2Z+2TxWud7FfGrYF+YcDGVEOmpCnsfv6HfwPKC1nwnkY7iM/S8w3g+UQDgvmZQ4d1
QFraV6tvMeFFb7QJbZupiA8cUeEtigt9o9SmKI0ewuCKpwP4TqrTdBHF7DuLQPCsLb+edrq3oQIZ
LrVyoT3tpSV4bDbaYED6E9/uFmzNpBBTQQ19LlmZFuQv4kRVHH58Edrwz8ahlj7Y1Ihzn66y5UXb
62f+VDJzl9MQR9ZOxCInM87uaU/6lJvWT+G9dKAwQQaIiJYkUOnVb5cShgqKNzxA3zeWlwXXNcVS
uCrHhgOe2uIqbNHx8rXlAnEeUHOYYAYEF9ADFCY7qajwVsyCraW5wc0a4vjPOj3KdGIHTpgEvAwa
7xQZneUVfdukWGrIPYBfATrZwnVg4wDd2qOCENWDmrdGaku4dlYUyxGKLjqhq1SLqlJDvQ8auXE5
p3xTeOpxVW29U6aIBsUlEDU8OsJbM+0QziEALiSsYl2CBeHeEXXWh3tHjp+e3f4uPprgvH2MO5NR
i09rUcl/9WzA9y9wSXzFiwwbB7BdmfPl+03Nch/s7vht6/rby/ReAFherzx8NDhrlY2eIyWz4mQz
Qn5cPeh0wTpISFKPM9nt/3YZK3wEOzKw7KwZfTdFdpMu9WzcNXIbFqbcMLVWsy4Soml4daI9Kd0a
nFy9F7thuP5zV9/X/zr5NCbOwNAKuACKcZJKbTasRB8MDULXChlZYHtTKBLtmI1zDucCVjd7ft61
SDDk9nkh2n45I9UO9i8yH8GoLSltm969kGhLKK+T0Hek2vggxl+3dSsDirB3QIJjtzZGMY1Ule8p
dF/MxSHOwmZYwgyCIHbHKwBSmtY/RKRC+e4iauMetbCo+AlO2KsUpMHjA9IeHXMoIMjrAgwrlRUe
N1mFgCtXb4/9E6SwkEKwHo23ZrSBQpdQBarNBdwUvihY9UFYva2AvZgMz2UUseR/VAHicKM/qTf2
HaqfnqjZPaSrYHnNfJdkCMvhiEEzYOBoZoShn9zAB20MrMJBr2hNkeLLl8Rv0aU+0AUSGe7W6p8e
4vdkJY4FXEvOdwSXq5lwX+jCdDkdbxwVglSPX0BEY9N8KMnZI6SebdRIvVPvIq4OHTNTN0f/w3so
D0Qib/U0w87/haF1oX8ShrbrHKnVA9leBB2Yvu3szHu+xZYwsK8dQCjDkmvL/zN7OfQvcMOJ8keF
MHE5Oi6sDm28a8828HWOVPSbSMpT90F0zRi+tt7ASDAxF0dlj7PTEgXHMagmPQegj5qwt/4dv6rd
3g0LKvtem5hSd4qL563gseU5vjMIim1t6GFDkR9vG1gwpSfKzLvUym1syA9l7YIR+WoBswUBsgai
o58l58C/MSKlI5/HE6JgJPyhI72DpDJw69thx00fwIx9KGeSfP1+2kyl4qk3at3QHpCl/DU2cX1D
iHtvRymJ+VkqeZkg3xN21RuE6qDFgciNILUTZNDVkS14qAOF5ZQ5OvweoXQZmMjTP/mFWCfMl174
kVJnec/jle2+v5i8XYmrrrxYPU6YINe1wp2UC6rAfUv7NJua1EYrBTG2ng7Od7SW9j0CepW2vXks
YUoOd0ubG3jfdZOhr4Ey+e/r3AuQMtnCFd86BZknX2Cc04+YeO1BiXMSx6zNFNBDnIP07Eulb5xn
BF2Z70sPXCHY9TIP0IJS34JYOBk5DQetQTqJHWsWHvaxtlp3bBsYEZCbMHVh8ay0zAfVry2N1YQj
jDQAF69jOiWr1YhZMW9rJZ0+afAmbeWYNAU8Yzs7UVdef3u0sc7jdpLZkz/TwQPISLsC4bfwyetE
z5GgrgGQLXmxhK9Bzjft51PKQc+vZuN51kDz211YrKfZ1oyQJz+CT1j6mQ5C1fzL0mxKNuomEi9o
mZbx7y2nVhg/LjPHRXjc97FZKgUC5YCORZ1+P3UtDC7N4qIcdRiqsCuHkL7/cZTzByNh32K5Bmae
ISPGaEhWDV1QWdonSIkM4vvo/V3iKUB7FY0+3Ybo0VXJRsIllZOvWXstMEhXQ4Fn7EiKTHPeXKvC
t6vQgzHTOQcEhg+Z5hclzC1DtuQkPbaw7smJNfZd8R46YxHSX4gAWArfc7WNIsDgAQ0+ByR5Y3ae
GAFZUFR9kOnVO06Eo+/X+FCp/QYVMshT/6gGXQje40Maa4pateE4L8S2LeK6Ou+dxbybt5qjeInX
5byc885/LbOajaWfdnGpC8uXDZQY1ALIcRfPTr7sZnSHJeWvTwi3kcYhVKM6UqjIrsBp01k3vB5S
Ttfc741SdTUBr3PDBigZUPj5ixForicaasjARESsRWmpaR+Uu1YWOdQbWDRHJrQXWUoirRbzv4tc
51dlIEcjF0rhWFptdd/XBbhhYU2PJmLq8jdIX0Id5QcDkcsvAE0W6LotaxIbRyXVY3feSb3gWvz6
eHqXMbigqF+aQi97dAKGdhdchTc0A80/oaLZupId5CgJJIgaJuaeohd2Zb2JhOx87USlsbdi4q+5
G1OVnq5OCWv/JNTkuAejqIrpGmRPuf2m59Xxj65yvUPv8lvG/4EeyDFILVXJD6bY9mw8W1uLHBft
SGiW7zvhCgSnlmu8WWulwgCWn5VlFxBgKoPngcRQxkgbE/lI5ZqeqHCJsXRP7bmTajySMJMo/w3A
fkDnHGUuA9Z+1pY4WubGl0V3POGT0kezDAU1iOWqDdJsd+IwgNcxIBCimqeGLQRoMO3D7soOnDXo
cS4BJNTwhFHKECzMfk8NbiXUS8D2hyxNauIIRFJdsIEq2EAo8EgAmlTvm4E4wAefCE2cXn8tDE7J
pAxwM0sP4F0TARmJsrw9varGklhO7Lq7yBMFjNEPSw+OS2EJtzVT3FWtzVyTEWK4BCREIR5GUzl7
gFEFNOtsThSJ56xkUy2PcA6V/XadQEwexBHThgH1sHLTNa4uDeH9o5sTNU9bl4VmkmIYZDrQ26Oq
GlFSTsCDuq1dR3ZqqotqqrVP40MQStrJLVcKD5/LLLEUdrrquNErkhZOmbATMGHzgZsSq0EjiUh7
T6t2+VGvB9DGiG1pJV4qpSHXVuGTf6jSuO9lVzU11IqFOk53h0vgFSem40Lki6W9bRec+BMZHxHZ
tKdjHE6DW+wtHmlaYulkPybfSE26yDyzgmnurU1WhFhmXf4FYjrmeIFaIoTxFIqLT5j3CpeJ1UeP
wn7tPgjkxLK6dOMv3+yM7KUCDJRw0EUu/6m9Et4HlBpwgAIbXbxc0WN9J61bNPCedMskkovGS1Ka
P2lyjL1xzj3k+M7Fq43UoLCbEffkW69bdMn2+Mp7UEVNKPPNdYM+TI7JN7Ana80pvG4X6McWS+1Q
n9djw8csKujuNmSarKOmwX8qJlfmHWMsL67i3nXyYGTUexfXLJKC9mbtr9oJun5BSbo8+LYHVK+p
3n+UEVkFTlEZhkd/bzQdDiM0YzU6gaOz5xfAym4QO0gRRjyrZ0nVHwG81A7yLptA1ecOjwC8Uvu9
LQ0E78Sd3gePqvCp3mdLSwarjbfJ+oTBTINVG/iguBx0JozFMCkm4XQPJH1mcgR4/5H2eymF9nWo
znetyTwqV98URqsmSrm6ZanEMI7XkAbDmtF9eHSxszYRcQW109wflOYAxz5e2CAnXkdhshMnlTmi
I+0yeLkeTHKOVzapgsOfRBsao/LxgeNwadzxYyKESiPYSl3wpg6mJTZ5P/I6SR5nMUww2+DsecQ0
DPCO/jqJI3TjazR+MC3gGUP+R97LDVgT+xJ0iX5FDkgcEmnuT0+Pyn70K1gwr2ft7AcVGvY59IJu
CQzuiG30ZZX3RTEtKdrQkE+kreN5VwyEHuBJzV9Ex2v6sObP1rMNOiz1Bf+DnsKgVGn/gOT7netm
hdKC5W74v5ljrQiLtlxpqBypc8y/RnJPwzhnOZNEk6AIQz0PP3yHlq1VzWEkH/MGNGZU++ShWEMA
tg3NwKBpJhs49HPXY4ph2cJSvDDpHaRmTebr7BbUYGa/e8tGa0nvNujlh3yPVnis5Z2//PVJ3nNU
8RfucAnMRRX+TA3uMHykdhpYagROTwvPCk+YpiZ20ZXKmSUdkXbLdz779YR8bhFWgjao8XKtutii
5LiuHzpzhHhKeYW8IAgS2TBo0BCSB3lUIYm2bES/xOknx9Xt0ozsJOrNYT4KEPi1nyneLWjU+RnD
2BZcHCapgwXSfPyaHvL+98fpMrZBbr2D4nvliOdUM1nv5KEMtTsOdRgaHHPrYf8rSTgtfguubqyS
E9CZZvoR/LlLha416WyXqW699D7bseHKppNmyWDyjYCIj5GH1ZDRtLkQlkaa7uKyBNe/Kyrw9tpR
01nqNJSJjaVFtGmN916ubQT0J5XvuYDJa097lWw6nLnkKi+/2vMLXNQ8BjUFpYdeBrKF7OWfRrOO
TCnSKGhiO33lJPWTKWVLBVa94H02B2qBcRRp7GdT1iHyXp/zNbQd0o1ZJn3Ti1J0y7lsUoCwjkRa
k8N8c7VhJe+q5AMInsYMu9lGYCO+9zsrVumIipjK/jfRwALvb4DuKPdySSgzLcD8iBMugUrxxd30
ucCHDgqyJkpmlywr41bVxGily/RjMb6cpJNifapxa3AKETGM5nwyzQURc2grQS8hIB5bxOcsJTZT
/CenvgwEe0FKy0D1hRBLJOvH7pNjM4WapohUuRRNNw7zkHEkGo5nzgj8B1ilhWBCrbND7QLYHE+g
Ueyj8J1wuMyEo2sYYl7lRgHDhz1672AkBeSdzBYIR0UsQhYX/14nPl9A1SaGwTYd/irxxmLqRpfk
p9UgQ2b7nfyrdLW5YAV6skm5KXjMe4DMJ5TRN4pwGYks+wmL9dE4UrOqUDasXDL09owOa+m5O+iZ
V02Zv2fg6FA4wm4Gk5fVLbVXJ0/WWwJGbKPIhNIbfHwdn+L+BEUuQ2FRspVOaXDYhLWi9bbBiIM5
tKefoa+/ugOCAsUEjI47cONZ+WM4Jja3ed7xK1Mri6i7sn2mfzCNH4ScbGkwUMVVum7r7ER4C3w2
f+erBFkxCT2mt1RSmEpGUV2F/ZNQIkgtwHf8SOVRz5mOVQ6fFVbAdy1hK6BtkhUXxesqXR66EBbI
2BzXGXM1rk4HT+YctKkmeOmdE1hmEO1IdVezRZPVTJaJh1MGhiqmveqAcoLnVaUbYPRmpWofGXzD
aZcobBwGbQ11wSBPQMWHwyLbkztrQd0ImmEZV5GC3Usrtb/XmDfjpWGODaenbrS0i6UClzsKVdpj
6YIzn52Px7vM1w19y0cdF43cdskIwOevx1i4Ic0bCr1oo6+VaJiBcg9U5IYD99zCPkZY4cnSR2nw
VIlXA0rTb6TyUoIgLr011s30y5A3MG912WkH4LG6ohL7ZccXHXn/Gkmp4IPAoxi/jO4B8wmYV95Q
L5mkbfzajyauRJEOy1RxOyoovRopKLIzK4JDd8IqCc/9xjahuinAoKCCc8uaF9uiQAjkrbGTyS1C
yrff19u9DFoTR9iGldN0SDD8zQQo7rmYCfKm/EZg5BnkGMBtqoncJRNiygHnk3ibSglR4KuxEQr+
BQDgYfTNB2M3JKZ0C1lTnfFgK5Z0sXqi053mWk8lYeP6sS/FC7IxaN3McDPJl+ANToizCyBKdFlM
gvvuLlvHPB1WNouZY9kwN0Nm06QNq6xXeDNvP4YSAQ4k9Ebs1P6R46yvrSMyn7KoNoH04Ts5A3uy
NcZ2wnC7tJeNtBkQDT5fx6dq/rnI1BSIXnvU3skMiIUoI+6XvrCcyxUe0cHZqijgCeGwmjW523UW
PUC8xfAjTbnyQKUOdthTtQIDnNwtP4ZyNkfw50tESgo2mpGP+LthopAhPUsm1gq4JcG9I4/MhB24
KfzRgGxA6amheCrMhRNiYg/cGkuFCI27UX+ZDYGcWI5DvvzKSgZmG4ki+BPo1S2dz6mSagC0p8A0
f/jsyW52pDCshi7F2mvrUKOrhz9fdRYofPZUdIWahqRAXpAdFOjFUujlj/GrmxL3PK+pwYo53wvP
X9NCvf7VK03zSwAEPz4K5k89jYoWT537jg84XBS3d/5lgMuWq47M8FsQM/rn8sVIAjHBX3bPw7Cw
FfavxLUs5aOs+faChKdvgGff0zAI3maO9vQv2/IpplnKKTLXtcCLTH9Nuf4WPaQqaXYMwGYAUpSL
41jJEu6vLUYIcje7B8Qho4mYCb854z+TaAW0+ScqIKQPWZ7Uxnt/pcaTCxREijuF34rb/FpBD7Gd
TfWrXAY5jwl/vlKAfM7bao0pMQIGCJWZyhJaiA66nSFlyq8ibyF5CM1CS1o69dHuNWuwvtIzhhZk
oArzdKagZ9J5fuhum1HG9tt3lNvXEwxmyjHKPkOLi7SYMf6fyhtaFv9VKeNJOaO0ujj4yTP7Xb3O
O7OefVPAD6YInP5nwI78bq5R5wj6E+YYAD+0wcMGB9F21aMY5yBx5Yptd2ZuFcD2sAjq/NmlwTUq
qvW2BxNeiyeP+ixZeuRzSwkWNOFqlyYuIJ0fxoQdgPPWqQx6lH1UIZi7O7iCkEmhvKdqm3zUXk0r
wub21XiuNHsMPfXfYzGxBnBi9EcT1teKg8dC8VEw6tvMNNN+msNvac5jF1d5nuyf8sGhCjONeM8l
lTEu384GOOL/kevm/+eITHtrsB8RscRnJdJFxoR/2G6kpe9kS2d8QiqYVOdBckRZ26QUYuvj8/Bu
EF6UBwsWKxDPVO3MnFb+wMjQTUBZQW4FwqWm4FtxjhRlP/M4Ma9eaAYOzkANeztUcjjCqIXg435U
Q/omR90eBfO3njJo0xGiw/uiyrAT7AXxHqtUgLBTA8+X84jilxm/Z41rqT7aoN45RLT8xQ1LJlmi
6SSJLSHlvecloVw6UtorE1mIaujtD4YEGFtsFpu2Mi7GnCMPRPuQ4DhRNJVftyE8VYmD4tAcLWtY
W00ZTnLVd9aTff8RyN7YiAQQuV6RTxBxcU0lfKbXs6n4704AZG/iGXkzH2pAG4pF5WB9FYrvH3t6
M84+WdyRp8sq/egpyFCVZKVi8lPz38jD5uTviRHrMd0Tnnw2VkWKOZ81aPWstR6WKFvSc2GyPA/l
uQMUSkRE4qNBg6VDK59Dhzj7dsU/2K2lLtCtENOwkes0iSRejVqkDaUgNalY17n31LaX86/Fe/I/
y+sOFtN/UB/+SdK8zymkb52hip3rRF0nFVLyXS/7djiMNNS12cBkb8AWTOSHQBSorv5RplZeC7tE
UeF76VyB/76KNTXn1M6hzvXlvRGhz+6shRplzVYdXWyW39wOMxuMYt4tjL7iwD46xFEnwtC1Cu/7
lSXkYcc9nFCE0F5Du8x/kqzGBjsjiMJKMI8bfObliC1VzhP6EFN1bdKYOnqtg3R50UzsEDnh9Y1+
ZBRv2Uw9IGIDx/q4+G1D2Cskqhek9xUSra4ulyG1FEyYEERkgP20m57brf4LJattMEx6EZprfkAd
Ndft7OfNY+mQZ5jyyBYDGuPpO7mX+JPYplwnvE0/7MGwrmJ9tUao7NZIUPlmfrY7t85DTdho8D7C
njtdrCOHDXFtPyIQiFYhgM7TVGDY7UgorIF5d0Ap8AQIt6/WKwPnBmh+YX9eie9hjjCmnbXtJC9V
nIc5BYvZwHHG2791Z2Abw+JrCghdLwcpYWTbb5OSqp37VloIG4wQ3VAgUsgdbU30byDGIBxEkNfa
GI6+ifLRhjh3jERHoRcpYnQQFft+XTwIgh/+CHUb5j9SVOTT/yuYsL0ekoFblogLqrsrsPS/VJLD
PUwQCkE83fn6D8z8J2hlpyGYC0E2SeoyLOfGUr0CJuTQ043cQN2339JbLIKp686J/Yf8aA6rN7a3
amCwt4qJpj9XkJlhubRwBbUwG41lCiz9OlM4LPZo9QmReTKd/v9kFLcB7DkLSm4HuytVL+mHD3RR
04cJYU+RmpmQTEuEBnL6C6ct027lTWmrecKsvI1se1esYk/RGze+br7w0i/UWTrtj449251fGAOm
t5/jazuc/LEj9TUpghFU4wrlwp/BAgGD3z7RiaKD1AdHxeoIBIqem382Xbe9zSNEUGdhLePnSBD5
m1T/GcD+zSq+4vSObVN8UwfJIP6KK61ey2RqckhBXp1IG2hJJM0to/XIX0vaw60yyPF6i4fSOsSz
e7any4onPM2lJUbJ/URKqoUYR4+yk0GVF+Ud8fwA+FmNlTTU103VnmjzWOV9NdsvCfhQs12bCcc6
wCszy/vLM1ndI4S8Qz36cJqO8jWmIOXMm5I6OmikLmVSfZWszfg/1I+OwrwY2sBEEloI973/UrNl
ze8ikr2O0I1O21b0Gt+KMy/nRqgLj95TgN1YACm2XoK3zih8cFCFi+qKwRDmwHCdc3WNWUWDRZEn
t/q9ZQFIoV2TOYNwtlC6Ootzy9XjCJRfd3ZpumD9Z5gEnb8a30HaljEJ2TfgCf0Wck6qUqkxWotn
GApuQVIaIOrb2ogoeabgJw9/pMEFfGfiQuljjlg5ZRwbcVNSLF2FR64vNGwPh3BFutfz8p5Ju5Cb
KnSceGB2/Lkk6jPRbPlBSn7gyh+tOpgY2LSygzOif3TN/vve4v4+H2LPZyVwunEdEfA0/t1yWi0e
jT+2jFN58L9ILAJ+WDvDNzFMHslWcMKMdPoDMg6tptx8loGUKrgLBvpxtCZHMiDBClkkLMTeZtwj
C7iUDIxQlLGUK7qRmje7lznKascvLQy8hrd8SOcGJcZKoEzz6J5g6P5Cnw9b4/OpYTLq9D4+mMSL
rYhgBBmk667xJy6Kvs/aeLgSzIFgkAiOE3YCRiPDZl+pyLAFSwDb04sAgwDL/lOeGT3gZeO735cq
1knzfzSzv9HgERF2PayUltk1CWHwet/DfkkD6BTC7w7aGkV57UYqCeLBYEhXAicOVnFundABOHkF
zNsv6HkmPmhsLfrlhQ68GabXlaHnC/wxY0TCgMygl6mTCDOb7YyCbJzQHoTsPvA5qw7D+CQpj1s9
2fe3MjLHfKU40jwms2y0D/POuOk6mGiEHk7X/wWDMBfmOKI/qplmHyRhrd+X0jQRTW8a7kV1iz82
goqUitP+88C4BpFBVA6OaHKX1ejKQ72MlGT+rvIDteKYVcgQB1ulfaIW4r4A3KwCpisYPaRCqmLd
rF4Kr5zEtllAnHyO45Dwm7cK9yNk2WUZdGe/5kcbZJu/eh3qjDmmFXs4Pa3uo0i8eg2NXhMIucMm
yTlRrMUsm3qTNBgB4ovNwxZTg6axihV3CpOL1ljTvF/0emRQXItiqG3GimAOZzzDjhDobplz/vy4
6MM/EUleFSByB9o5z3XPhfR1yx/YLwKKAMoXM2QSI0sEmWuMIoSAhSGj8MzuuCM4Iko2dJicEASk
NfckyS8Ujo4ISN0tKAl6l4R/xkHMG1+kLijlf/l5HgQq2jVuZ1kja7eFJrk6L0hMW45YOuO9iL66
P2hEHoogyNmGhJhcek6XPfJpvRi9vjDjPLaemdbdwTuAwD6SvjRj3g6oDt98v63XdkpWi3ATl3N0
xJv5CveEY/e9DCXb2l1PZJTsHWSFUTV/Nk1sPY8YJDUUsILvfJ4cHymK4kveP7ETrFVgVMcaMpuw
IDFuso3XJH+9eEzuLB+KKbveiFIC/P3U6gfuI/fy43T2TgJchLDxEKrl4SGyiyqFmhBhHVCC+s4q
RGBeDnmOcz7xBRgJrsrvNDkW99JJrPbJ0UV4o0746n3QEfaphbWQrXTKpJPQO6H8117xfrSTyy9A
CwChqTcQ5KCn8FK9WkYMX9Q1CLGLCM5gg3/E/WKCcTXRz/jrDc3x9cera5feuCjRJxGFm6U8aLBJ
gMVdca/iUQ1ny0rAMoMq6P+EkMUlxYny5AbJLAft7nXO4kMNBcnBk2EAog2q5TlVQ+C4YuVLD9Pu
m2e1MRs+O/8cjLqT+H/IDoh9pdI/eRjlJ10Cq30/8OmYlR/2jmVPZdFjzsYxR70lNkI5bFxpRZTR
UEae+nFrFS7kmBRcdWxE4zTakTNe68GcTjEV9BImmytLzLqNYG4AbLeOC2Wa7Ek+ts7BG4QbOvSi
OvRf9ri35NyOsVmI/yZDVeeNpWuoPh5zRnjSk6ZsLwCpA/98npapB/hpwxjL8+1rPE/dIMg3rFp/
py+rnS73vH8eyoP5Ua7uvy8nh4ecRcAY5BiRhZBvRxdDbkOh0LUHGLoh3usyEAAUP265C7mnJSrg
R4WDvSZKWDQ8SOb3ycFF4JbPyqe8Yc5WqPyxCiFxMgSmEAFnLEAFkDu/keLi+9i8r4Zs9g6PWrnK
SudTCMMx4qSyPgLKxV6JS3/QuzzeJBRAndUZ5b2WZD885E33bRaX9zkxpc5fJErKZKL4DkxjzIaR
0864WZVOGLtwjcUjinatKHLGZtyy8k5Z0O+nZqwWbdosC5K2PUxh/8taWsmgevjfq6cX+SBZib/i
VqGtJEzhNCxR1GoXiC3oY6gAPQnZvRKeMd7e0iMa9NErFDPR4ec/gyLXtEmVKnJ93zKJScF734zx
1yticFzaFbW2qT0BrjtcPtrWVoit5bUtGC7XbHP8GQk4TVZ/Ssf05jRNN4muGlBtTK1P0f4vBxY5
XGEmtjLHEMEqTDHnFGCfnYlKt4cVgwq6spVIh4J6rdkAOCqF73hAO7Bz/dQHn1fEC+RgG8T+hdE+
AlboJP+deToYW/A9S9/M2dW+1Gc+auB8lVVbem6s3Tuueg6i1UHI9cZWiv8tcEIyoGWZE2IL32CO
qCKMHQ7MSEea47UQ6CiExbqVGk2r+krUEKU9vSDYpqUQRK1i4jdIV+bU8vjc0B5Arxf7F9ktmTgk
L2POsj0NI2rLsmPniWBTcLdy6UFEDeDnL4EsM+R0eJkWsRiMd79PIu0OgSxoey3kPug+ZdGr0KfM
IfjcDppMTbLTMw1WXvmYtLJOMKxgnJzSKJRFnQS9Sct85NqbfArt4KvyR+EVRmfEAYy57vh96/2+
jLiT8NTQ3FW+NLMIt23utI6zGcT+MQqOPysc3VtL/Y1E8pkm3RQO7X2SZG167K+vn8NwOkau6jqu
LMxFNGlXTBljGZwwCvaMHIE6ZULmkX6Jm4B+zUsgSFw5+P5udO2TzBEKTSgE+Z3jtwFPWts0Pc7I
qj1D/bGdPwT3O565jj0fNqCnbj7b7rJk7j3UKytvRnI1Fba8FYQAc0imUF7POJH0ikojX2NI5tRc
Oi8dT6VpzZQ1kx7W2JAxV3B/NW2kUsEb8G0kAWL6nzeTCCAHzdKR+wNRpV+0iZM52fkcWWoMrQpW
+tiY/nrr10krjGnEwR7RIOaqygZgsAD62OqWAIvvH7Co/JTvKPVVxlGrw108x34fmVl5cxpLNfDE
1t+uD9V8TGtZO8CDuk/gFOn/7zMM0YjpUiDZNOUtD6nYhxB66Fo0n8CnYBxCJD+UO93x0HDkIca4
mU6yvXRCh0tVCwtO07BCUjeE++a5FMTbOXpXdG2+nhhg2Js8nJ3Y52s4VlUDac7OztCdqFr9Su9y
oYFyoco+cVtG7temWQeEXaHKDEELgMyvWES+ap7veu/opShC4dae57Dwiut8lMZT1KH7hNOaTSbV
7EkVjFnUVG8ZM1Z5lHX8Yv+zUduehyrViU5RlkPGiPWS7E3U9rN5DwiK9F07sRwsnRR+uUbFnCGr
E8j5tC7fxNO69kAbWVb0liWYJpTg+UKuVeIpQB4U71t9EAlEa9nZRR+Bw31dqCoxkBrI4qYYTLbd
JQyns0Jq6wT4nu6qZfdvHTxbdsHM1+HfUsDg+oDRqx9pRuXgQqAtFagaK4tRnSQCkuyfrvVJV7lq
tAvJip2fg/jUn904ds8FgzIzjgJUOdtcaTFu2xhC7u3BkzQ7ZxJGK15rswPVFldZQPOE5TZFzMJO
ckHjKSwS8I465O8cxl46awMPOsA80nK0P/6TgEYbDlSZsESNlL1WuXLwCq7tVwMBz+eqm3QCaGiq
KzQRl0h1KMhX0emxkFo27Jd49kYnaStqMSEYwdFCfG8yZfmTWTyHYdnhr/Zdc4ZBS9Xh3ftp20FT
lqHRukSlkvVfmbQgjP7YjTCgM1DUZsNkxMbM9fYYopLFaRr7bxaLU4uM59aZo/q2Qg9FLm9vVUZ0
2IOJ3CFzPmnKM9LG4Fm72igideJMxgdg60LvhjqBw9KP6Bob0mnCixxs4nr6Q9bqEQAXZ3UZYWEx
3fiEZ3YBjEkN49yrkF4zsjnXZrULVeAwoa+sMfNY8kXC/qpxsdzpjuQsa4/rF6JFU3+ifoMD+/Gf
xntjdHwLBqx15EbNXX5SV29AlzdAsM7uB1D/DWt7VMSCBa5Wh5a8p6+BryEUBBqk57iIN8zJTqdj
n0OHM/WJ0AC2qn4Kicoih5///NYThkArQvVYu7kcnWLEMAcYGYEjW9KGhVQKwKy0ITT6VHOYunIh
Vgfui12fdAVTg+INx/rpHqjjAOCo7sMTVw+Bb5msq6nByU2huG7wOiiciUhE11O/Gp3iPXCMYQdb
z0hwR0Cn1ISfuXC3pjrxFMbiqK+UA7ICR3p42xYzDSfOSuvYxcZxSG44SRR4EqdHz1R0zFL7/BQD
mDKaU7ep2BrQacijzBx76ZcDYyoxX79jDVFJDgp+fTCZQu1xPaT06rikel2ROwmRl/RYX/srLxTu
RD9AUYcFunJKKw+8tkQy0OLCSNnMMM2Pq9+WoXmSk4xq8Z24torUbmpUJnWHDDjyM4Pq4g2WoxIA
x1tZ9pi9rWhUB66kI4FfeTYFxR6aPY+W18p9wkRUQB+BP3iyKipRmO2cPbH8AWv6lGOsdkmZ2tuS
GEXp0hb1MukibBOg+UFAZuCbjAiK9Fhc+odLxQKuK4mlfl76JNqweiV2nw4dkzW8ytE+4n+oV+dR
Q7ohmf4h3SS+aa2Zuxo5po884D/RDqqxMMKNqFcDqBVXHrYds5h0oMwXfAChiTeeH3DMtMpWhUGC
pFQX8kv4tUNuriT/Is0N/rO4ATf0tiLuRULvYQrI9+HunLqx4OitHbR7Jpn1ceQs+B3PihVq7HPd
m2hgUsP5KFfUcUY9HWvgIRk2H/Syij6LFOdH3yn+QjgbQW5tW9EWiKpgdtOcvWgTCI0v/QDoJ99o
x3e2iBTWUuqTo5qkeFLi6E0HReTvcazzxgMddtdQASn/yeQUzJzYQPLc530QbopjF4PZf4GfV/aA
t3GeFfDMbvyt4FJnwU9NZ0fUy0ZmGIfMWIUd+IJweatoyP6mOSmPECOANs7jXg1/AhGHxDUo9Y74
wSqAD6hHBO94W3ackyfN3Rua4VgiXRRthxoSwh40O7pLPyva4MSIckEHEvIVCdkF01wfGYDYtznY
QRHbbjdtJJhI3MT1sXwkvpfilO7/IqiUsqVOl6qFR2CzE/eON0fhWjmEoMEr8yCsAAO/HyNry3VI
jMmqj6dZJq6MBxX1IceXNXzuG7mYmziMk+8wTcScw2hoKeXIpuxxEWDIPF7i0dmnznH6FXqZJGip
8ci9iqiFnsCCucZzUF7g2WYrxDk+iDRjDbmR/uPF+WknKshfY4yWEdcwVXK0pU6P7Ga/X3bu4iXz
IcnA+/d1M7eBXRXSWlKvI67GR4dD7G+lP2JzgtHY5H05/BM+oKZ8oF92AH5XNN9A/Dwv8IDk2LGm
vDKkmy9GcGn1m3O3JsZyQf/b9yqmZPqilOyG7Y18UFjk+ix+GLqyeLmCPF044qQ1nWxGKXuOA1RE
uzjc/TMnvO0d8yq+8ItfDeR9Hc+4+CAw8/ffT6rppqomdfUhQrG3mq3cDVnt5Ju020nRHaFiIrIj
TQZsER/JpBL2gsjRZoItkOYeLePXusxZoovJJpHi9tfcdSDxF8hvvb8NFbeK/Ss8lVZaqDk9SpQm
GTi4Jmird5f25siISp6Jf8ttTqWwLwkqM/dcKGDX4HvD17H6HHv+/QlluBT3HlD6EMiPspqCvMFo
89b27PnY9ZdXVvqWp+93itkqh0ppBQ5uDwsLABwRW5bEGBfFyXsEkxhw0aTCQVtMjokJhHq9gQy1
gYHvV5w9RaMMBWmRmhE+xrpngZ9MsL8AE9qrenNkC32QBE58P4FhOdQ8jK7SsU7eu0SMQYNNAjyp
QRhuc+/mMwFQbiGs6RQXN7AOKidyZa6AIw9DtwzmrAwei0WhPRZ6oxI6acyzs7WLj3lPCxDbtTOa
9/o51udX6Ly4pZTfvI50Ij6M6uluMe51EvCuTrMVhc7DES/WS3GKUzAoLUCxbsV9nLy/PcpZA+Bk
Pi+08FcnfS6ToWvWKxyux4Bb4ukK5xJlHX9qX+79IcChb6ah2InVmCO3cCx0D1gS2ugkP0vwUStB
xEgDUTSaKqzNVYtCDrr46PlBuMbLNjP1ycwI59Q7E/YpWFaRBY7wuw1dhjnO+IazIqrACFvyHo39
v6BLqjGTszVJUzqQjgjPxgDKIszRTFl5RWAjj3s5LZfK4M0fXv7rIANR6sT6P9kOjxrPDsvzUNlN
PjOhHMtuNiiX18QyWn+25ZasiT8R6wmOa77mXoNRnvg+50rtAaFwqH6aBl9hiK4mduRHu005W5lM
bQw9+91Vc+Vk28GjmCxul/1TDWxbR/QDuXJ7U9jGUGungjYM+K6C6K5QlOj8FU8HXq6a6xAWq9I/
OZWkWZ06ourhc4GtOrBJGgJwtnb2k3WZRYZSJayMS1VF05zyiG25yvmr+4kw7exy/J5o+v1ToI75
9gg08O2Zaik+qXvPefxMi89HkRqKm7aWeiLZK9EpgtlhWUy3SmqH0hGac+MMebh+ifRQxHQknb9L
gb4VbUZ3iVVuD3xZjVZWHWRQ29MBxI6onTKeXtrZXzGrnoLcr4mSOmcfCEwJfMTNquIgynEd4P2X
qbtjk1wrn31d7WPtwyuvle7Gp8luQwGChbOL5qjkvtgCJx1OByzsgkfLmCG5eBjU86ZWHsJxqyTv
yQgnOTgIx8P938w1sUScfoxQuRRsqLqt69jfUIKm9s98qlagWazwib3Z3bWfYYeHRB0LVJLmQ9Cl
7ZMktolG6pnKsHzx6u26PYMYEuKmxamXua0X76nnWF22dPmD5SKThdP7RV2Wr2u8XDaA0wcd8UeC
5i8s8vG2emGaGyndUpg/fhHBGhkx6eTUdNibcfVeCuZgluhSfNxWXU27Fpv2OU9eDYbF+WzmIw+W
ta1b1feDwjkN7mOytmQfVAJfOpFxri+iRJsNiEg1i8VYZtoW+u5KiQqkyVvx+U7dkN1DH3jgkmYG
m0cDNC6Vz5WbXehfWiDOLUV0B7GZjvsbXNXkDHvfiPSo+HLOfegGXTXFZ2psE54AzYYzb/eqfAcu
vDWjSY9Tsr7IAdShrQ6fYXpAnabprrV0w2NpmbjG0TYOJBFCmtNs64LABx5NzdiW7dt2I0GV//cQ
Wc5VKIsh8DLcDzoqn5hPIuHjOzxaCC5P9Uhjrj0YIiOpb4LajBvsx3I3Bg//pEXJjBassMwni0Ie
t8zIynfaYdfwFTx4ViCSg0/uiQIq+YN5/XHno8m4N0iowQuzU186S9Im5y9yiLPANTz8LnnqHFkf
yMKdhWzLwkjQ2BdC/nxVjBojx1fCcTPYqMI5zcccYveTuEUSZ/DNkBkmKz6Y2bGhLGedo3kSyRwy
Mrpe4xpBmVZR1MoqArVuiY0GnZq2f7EXhAA6M9UihrpM3RBI7EljpPx53PhA8uY62zn/bkQfasbm
tDRC/H2Zm4lGH2XHyfJG8G+jhB8ZrKtySDWY6RuvW+UKYMithVRKwQfFFbocLcG13T26GPqUoh0N
6LAE7ND/X/20auhY61rg3g9Oy2W3NfIIRJvX83IAGYbzVs9Nffhmyy42mqWNfWdzAstYwLRXmomH
p4GHNLYOI3Zm7g7s+Y7HhT9ZLEmwdlfFhtoEneojs89UoZStbbCHXuRAFIWrh5iTOmEys8ijyIk4
3grkeW4RDW0BAQOO2G+V9oJhXnt9q+nKnamKafFK3W4efkge0RiCoEj9XTw33I61Wg+XbspxzmTo
FiJrp1rQpfH6OXryMVfkFfllbBxx8F3xV1NqYb/z5wCK8SkKS8az++0CSYlyVJ9hjG2iOYhJuAg1
2MxFR3T/+DINtTvuQeDTR6z+wM5o1+hwyBhI0dB2023ZXfy5sMyfuuPs/eZpPItF30Q91Xkeczyy
upTHBNCDb4orDiQy1PkUmqOcxBDeZ1iONDnKkByV0+Sx4H6Wn61XhO5T3Y2uIH91AmYXWgXsXv4W
Ovk60D1datWngejBk5Ek1SKtwHZMMAfT2cvtaWBJKkvakjOuLScDFMJvlP0S9mGipBVTTPCTyJ7t
1Jc/ZMrw+eoLhUGgX7y7KidavviDn2Zv+lK1oF3DWqwNjLPvJo2+DC3uotC9hltK+sHrWu5ysI5m
b01cphjROXIzrcj68DybJ3F32bVUZ56uZaU7xwVx1t1Su36XwAWr3yXe5VWCqqXToPbAf6JserQH
YbRbh91h0Pf7d9kf7Q+TGjDc1TA5NzPqVKO49vIIc/gSILqJjw2KkMQkwqJfvrS8cQ6St3o5czux
0xeS5/8M4o2KoOk7ZX1KBNLsm75vsCDLrBouHgsv000UJYer/aTBErfJm2B6r2no42wCCEWig1oY
G9RBnZbZh4RDG2Mn0O8c2dRAzALJcYe31WwIMGmOTOQtDFAObArk7KcgfatgSe8FGWXCug6VJPZg
Y1S1GhF85Tybxf6YSwP2YImmNr9DS1XnCUgb/9PGtVq47SVI833AMAgpzzzuZDcBbiTTD8Ua6N9G
1dIeILQp2GuPIvz0sd8v09xuK9aaLMeoQ1UZ7eOIMZ2seiEhbDUciLNIm9AC216GS5Jv47FhSN6Q
mi5CzU1dR5t0V+yZvO6K7EHYOsNYlWIpGTIY4seeOfyoGZGCVe66pP2EtpLlejeIJBOhQmvKZZtC
IxsGBwEEV7OpzwVmt+zJXexwjPNAYz0bhyWUMyvhlghIp79l/dD+9m5jfEi0xuv0XG8Jz1gg2COH
F6n8OyiJ0RZUR1QBMfIzVJ2gGOZL0JRgNAphz57E4qbC+JGSRLwTBTReQpPBOZeq2+XWsSIfpU2r
yMCHI2xLoEvx7v+ccSrgZAFk472K+VwAAc3Iwmd4AlrFPUBI+8yuTMBaSMx2qRD4MYTGBot+8k51
HFU1LIO+TKY3OMKvddVbWm2IIbM3vfVv71gFo/OS0Roc+ejNiOxOpZRx1PJtOFeKaNNi8xhzWFn1
QFcJCY2A6kRRgo95doecoieQjkDp7XRXygS7J+lBLH5a7lNR2K74RUfHgSikol2vOmYCTVMJdSik
CFxyUJ3AhT/3FBhzllHq4J+C8v7FMcs8MRdJfCfT+ttu8q+RR0cEmFihom7FbrbaboUBek/q2aPu
9hAj8gvwXtHmTfcXzsMb2k9s1a+nbX0qu5T8ybYPbth8AmpJFYOFlMETCiYiqiZYV66NQH5ie0gs
RcRC9rIp3Mxvg1Xfy4obYZRqRlLDwNg1xC/xTm84tPfMHFurAQJooqp4M8RwRT4HxPApca1WAiuY
sdu9EKOExSJDIBbyENk8PtScA7q+I83EeG2dc3iTcs1elWTZE99PhL4HN49z5ANJZ+KzgGgVJa/q
BSFARPA3Sragdza4f9OvJ0DZl18OMnaiUndk50wX8qy2myrtpuAC1SsqIaG9XJ4jCc7a2NJf/Imf
fwysRkOM6UVgOoctMtjYLcJRXajLAAPGWpvJ5WU9T0f0cise4Fog6a7EWxQj8OmxnmGAWU7JVWwb
vBPPkBL7fb3cHXKV82NZ00Rs0JQHQKKe+M4blTXVU0/rDT0PERLbnFsxO3Ab3NLgRwPitFUDYGdn
z43GfBqhAvJ0SGIX/Gahv4RZEoFwmvoo9MBQfLl5o1CDQw6UaZ2Tx+P4sbh2AXb2kgOsrdaKIwvb
aD7pUto/Mf5lFcCsNTVlU8cOVTO7wwUQW/OZi1bY588VeYEiQsvHH4LR8Mj+K9gIxleJUy13rckW
yCOfds0uqEuJMwJJfTWMGKaY0uAIaolLAdE7mu3uR0taOLrzFUKaCz1ZP8MfMEMDuySIWnbgzNZW
i/E0TelvP4KD+oPEJi1ur6QaaSLpA7okbw6Up45z1Sncf9ke4LTk4Nui5WE5Do+E1LajyZXbUknp
PVS9MiUs13giRd5MKee0Z/frbJvg7wzPsUP3Lu3JdDifKuDiav5lP8LSmlfIw4aHvgdlETNzXWZ3
skC8LL+bwDJ8wHjBGhFjFhEsIsh0XagGzE0Aq+ZvXR6KdxpQ3BtEvWNYFnIFpa7qnBBizMuBPcBh
DIxXX/rXgX0vzP/2+u+lojxq+GP0tF3SWe2364MqY+2DsdX3b/0hLvyC4a/sweLOIb+Ci9UdejGD
fjpeTyxUX1CNUW+aUwJcsxLqs5xl1udnFtecgzdxrjWouq7jrt+0pSIGsg+PJ6jqgX4tdqzK38K4
puKiYRAxYXXg8WgoQNC2u5yT3djRC0AI68Ok5Hqz5W/adPXpyvhSTrlO1jIEJMBbf9a8TPYGeYgI
glXTUSb9xDTODBt3u78+AXp9Xpe+CTi03JxEHE8soYr5AaWIbO6c5rQ27Q2ixUWXmlI0Ocy+tNKb
Hed+whszfTZar8IehvyM+eRFEqlqbgMQkZm4jcq6O053rN057iGV8OEmaaHsI0cVP28bSDi6JX5y
Zwy5qn1inj19RjDA7Xkq7sJRDsSnzwCyGlI7+ACOjOAfObzuuGB5WviyxWGzHJc1aXohPklNJd/7
WdigVCtGY9qYUhki8dhRqEqH2sRhffCgPDFZYOmzVz/j5FKUswGBvxRTrgjphwIxCpjcoclPu3En
NPP0lMaQW+RYtFpO4p28X20RmZsBeokWIwWOAmgAZOdMFO4C1wDG9uh+AWuz/khpu1vNoOg7otVc
Q+dtoOzNDWRZYYJn0akgUw3P6q61vjQB3N8fcdC2kn/pVt5Q7m2QzSKnnWDPblnO0WpkFWxV+mME
Mh7BPt0b47Hzbqqi1zrDNB101ZyUUmebTE0EkvsuX93Vtr4qRz8DbSGOgXadE9tLAB1jyDbcCnOE
7itTza8Yd5WPdCTlEAF7rTmPICkDmFxYKRbHkbbh0snAkKAJSe8KiabtgArbY4QJGUyEM7p5Sqi+
18krH2Uj7usqcpne7YZCGaUxMNHGf8iNuvgUqwDqoEY4/7ZMMEkPC4vWx3irWd9UtkTtxiuBkEmy
9q2/Estnab7CO+rW5QEU6MLbE5XPO0B93NYz3fI/Gr2W42nQ1aNmOZhxAwCI+X3lkm78SaIBFl05
Bk5+PrIU1oLrQunpNSoo4uGQfro+OCs4HRxQGlv8Nscm6/32dZRHGoKPcFGy0VuzPyCvP2LPe1HF
93ad/pZQ/LKi6y+cR255rP2yCTXxmIjUcGg6O4GY3FDNvnk51cmzdjsql8YkxPbCvnvIyP64JxJ0
2VpHtrh/NgS5++Aq1u6pUXqKjpriU86wZ2E+350JbuJpxeIEx9sio80ZJ8dUfaJH83cj006Y97u8
WIR4Gx1Zi1VbbEQfMgQvxspk8JNaP6WwmNGXG3bhi1ngzMabj49lbmeZ3/nAx4Orq8XC7TySu5jn
vJTHSLRh6zEob2NWo1a7k8YvswUiT9tvBwyUOcJEMuOC1igf+BRgf4Wg4jDDUKVhF0J68vuiN9fz
OPX05IXjhVaMWva4SWkMPXilknkDY0XM/7rfTMcnvb1uQNeGOpRPl7aaAP+XC2R7ks4rn/ut5bEz
80M2kxSHPm2iYmZnnZAEqNqu5+oPjowANKmGp9SAfsdf4QA40XxqL39H3q9nw6OfZnZJNZW5osdJ
FiTQJ4tLx+Oh5/AD/mwvo0VQLZ9j2qMs0wLEuBVjSe+RHhc2fMI4hdfsiHwmjxHNBlqN5Ur5iqir
zH9s27N3p4MCvXerhICr3kG1vnuGfDSoPFVIzTRsuAZfBmFfJLGL4Ei+LmY/p1Nfy9T7s/BKz27N
3SA7cT8FJ15dpfcvbENkFSHvnMBK/02/lHccjRLRb8LhHikd8yhsyfhfWiFCCBiilFncdnPFl4xL
HyuBd18G173GIfbtKDxK9BChSJHcMII0ZyrP1cZgvWlEWo7x7smXVv7tmMMxR4u9qxKlPyXQtw7X
5wFQ3Ta9hik21cry1MDOnCb3TNwvcaAPtUERbRmH/qQclEItepHtbHCVhkAYo9Opy+I0JEufvQM9
CiqlNh3IwAuIj8mI0E7mMta7+Hv5NL3oc0YehjxCVPeu92OFVsGdS30n6HbsS0NZuiGvlp6WgT1q
wNxW6QWZ4vmO2UdECXhh5BbAg5E9zta5EnFOR10VtRC3b0o5tdOSRbPvO0/mujs8whD9mfqu5CYm
P/FbyiKXuEdx82S67+H+g23AnbBQm/TpmZH0IiNs/vxzzmoFKV/0t++lq2plK/YclmKg05xCZJGc
rjIZv5q9ZA9khJpyvtvJfZB4cQrSvKAz4va8NvmnsiZw2sVaAHQw/Fd/3ikB/tscLDxHA9l+dyHM
rhekSwU7m7qizIHSq7Na44IF69AD9AjU9S3rN2T1MV/ojeCHIZIxPqbaOVTe4+zFnJba9VsRrTlY
KGchDjEibxrqg+IUzKMtU5HykTP5dtSxzGXC75Cu2f1A4xqGSsV/TBvRVodcpmVUbO3OC4cnCCMp
VciuTuiXXPWnIdKw7fFRY/SeohC/mZJCfJ9I7qaZvOQJrtty5onI+GbjwZjQz+UnwJU0WJOw8BOG
G2Rrp/loj+B5UJObJ4IdaM1g6YqOx9a7zBBc9xBMwaae2YKa9K3LD/+mgxIXOvd/aH0Zz4o6zo8x
EaBO/jxRBlAOL9T8FinyeFe/VS0ki1cKZUQ/bHfzGzpEKk8Dd2A6Ey0n5915YHLz5mpCAUg5H+lB
rOI/4jxxKul2aqD44pvwQ22yXlRSUpLjtq39Qf1uWVGJ1Nh0dt2RDeLP0L9EZygBl2DPGqZL1YIg
Ds0BP1OQNydXR/Bz9wXWCrWrVUAkmq1UcC9Rep9LR1F4C/6bn5mztLRg9tIu8WgYUoeDaUKcs01K
Bo2Z/LpZV9J/iLzozmD0WQ9JL+FeqPgJ3vG/f4NJpE9wdu11CF6OMN9e5Qp1AaHOxXLH+uq6WkeN
xgxtiwoO7htBL36ZRUdT3UG+3cLwegzVDw9kk8FbSWC9QCWzgLvquUblHeC+GS7SXxRBOV/qd5+B
cNBEUc7U3Egwxecoz1e9x+e/gBu5PYsbf3JwhX8jd+LL8e3ADy5NvK//MzbsvUaJsl/k+ZKR9B/H
vsCrJzTad14oRt7KvwOtJTZtfaEHJVMMrLrJfgXtV9rV909epvTJcoaneeQRjs+H9F9KOrcb5ZzL
KTJRhXLDz4ThuUEX6y/uou8jKxDqLNDr8IWbcn37HkUqlINkskAZQTKNl9q6G7FyufYTUIqi3Bv2
v5ZNpwfoMQ7rcU87VAk3aVhPrg9o8C7bR+VEIQ5Tw8TRq6tAq3ZbBLhEhahr6mHTLWc5DbcZ9nFz
6Cy6Ysz3fTk/hrhVVl4I/ouEuxA+1liOCDP17Y/1ImM/iHZZz783QeDweh0ZuzyNjy5NYaMtvuwj
6Rx9QyZsWdjmolfXcj5HR1GjupN1GFAlgXJZb7xi7MDjPyuKrKXmc/FJkRZ7OfdwO0oOIvqUaYdq
/T1+Ey0hXruvzw5zoEoQ+2qlHKYIOQpO+BeQuKB1V9QCBI+I23UbRsR3b5NFr3zBvCFr8tpBZmqu
QZdYBR985VnuRlx4I0P8Cs/p48nW9LAG5G/929dycHio0SCqhiW2UALC+zlDUQVAwH86pWGs4c6T
qPc62nYCNhKOe8hxwpx5HWc0TRxqzVl2LhSFft4B7HhMwzqYgRgSXnBXzVHBtBH2rMq7E20Ef/ot
G1OgfeoEq8rv/wC7Tw7Xfe6Y4CTE/f7AUwF1Zx6t0ejOPvb7W7qyy9+zkx78uVP9+SVG2DZARXIw
M5jo30Uv2ey3yVo/DL49O1IpnpqEcpuuZF6o0PW77nULXZDm226lLLjryWuy5vap0oNDxBoGPRUi
xSkbiTRBmrNYrmc1Cj+29cZBEZ1yD4HSNlYGBq5Tc0cd2hvhgiwrxqyD2OealyMhWbHDAWybZ4kB
TKCOwC+zRjBQJlRTa6mQUqamFC/pzs0hXhLA2zIgfRiW3xqUYSepN4U2+eT025ODmw865Fx1ttH3
cPV4RoscIpHMYUcLlKzdfFEKKepsT65x2U5F9oo4yZhfAY5cmLuJthEYCmXWRtGF8kKkjff0iBg4
VntAYNBI2eDhPlb6GqW9t9U2dZdjahU4dykfQc9RONJyGP6QQJDYSrSS45g6kW0SrCNtIQFgtOpj
6zpcDpI51S2XxqZIolJK4L/TiuzC7lemZkGwmQOBNcgAiuAXSdQ2HDj2nbl7OEPXhkil7OO9hoze
QLFkg5IGnYdexfK87dZS8/6Fhbj9BW64JjEEBtR9ESMX0CGt+dK/udOiX7Fk0cyoFlKqEJmx52T+
ObJHxPlUnLLiyK9bMzjt5W5DHzo/dq6sfE5DPHA2Va0uF8VZfjaThu6LzjRUjz2QSQgb7M70Td3R
tt443i5MaMcC7q+g+49JJQGHG6mn1Or5qAgBuGqLmndlymhGLQ13phNtyOn3YA0GB6me5LzENNUo
3Ab+CSuWng/udbqLPEm2W0Ki1zNWvpdCpb3Hn7jADJejT21BfT958635ipRsgKRHZKh2z5sefw0L
HZyWDKLlOicAT55YRNGtKfvfMUqNXRK2ypI6LkQO5RkgelOpw0ImqCqWIqy33SiFdOXDpKXD5xRf
95j/aF4Omd1508hJdQt3gLrNdlE04fP87/rscE4tnk3bKwMCwqeLp4IED5dffdurUWfo1+kNR8ZK
uxVgHLEuuDPmP5EErAVTPKbicUcKKxvoHmC0ALyRaAPSx6/fcrX1pfzYQl28bVXgC2oz7VNYfGl5
f3JBCI9Vc1JbmJxQMfUtUYh9q07oovFsKPOSzX97S1pSa8Wm1sNWuGEtvh9PQIKOjnaocy2N7gHf
nkf28exExLl2j0UuqcsLJEtZMqa4jleK0KlgSCK20JwspnzdAQ84xPU7jL9wFGB6eRj7Lx94ljCo
WQEid1rzSUlVt2oHYk5pf2TYf3NVB4QiXuzweUnMRLxDpJZOmQEFv98b53+8XhYTnuVqrhJg/Sg+
lqzZ/FRq53aVAVnOg0S/L0hcAvztrHOphNaHyEPLKUtV98FbtwmhflmWY0m3SyYU1XNAccAMqwX+
5L8hywHQHNwWk9rN6+NVjselbqOFlmwgGf4A0lg8apC3KbtKD7U7iQKW3Yu7kyaMm2ybsn5a3ezb
kltw+5jmkmecojG1odemEkeri39fJ5hrQFcWcJFhuzFnijwbmJSXxaaWidHRu2iu5ZNuDweO2Od0
qEIvVu4Lg5ClWGcRz0qvZW2kBRqeFBipuMKvCxsdaMuVDVPLErEzySdjq8Odg026Xj247fkzXoU7
M4rD+QKcZY4P8aM4C7jw/dYqli9jHPlmip8ZsTaI0VWh5uI/sIqLC2dg3MvXP+23zrmNU5dSOf0R
NS3Uu04AbHHJtMtz4ZptOBtdj5YjEevWDORnyYaR2osBokD9eXLpqq5Hh8BbRuTOkF6yP/Zx2frX
W8vmBgWlsTz3oOOd15CDiJ0enu3nIr2X8vY+qMwU9kgb6FG0S3hLZYVHA6l3A2+4suztIlzT/DNx
LiBFoBy2SkczoL+d90cDsVaV/abZKUXSQqjwdpYoqE/y2gwFgMPZ7OiFoW7yahh/cRjIffUn7VP1
f3ZaMLr2noPbLgsftPy4RIyYLReh+sEdmuQqyyB2J4qROTgV773hayJrXEEYTnJBtOlI4dxVwBwh
7oiYAlXeR7AJ3bNMaFUtM2FN4SzCVCKdQUF1BPmBWvprIrUb0ALgmlm1KRo31bZzGgZnEGatRBho
7NX1RHys2qzz+pZl4VhtPDFWZYqbVFBAGgEO3cXtcYw8u/Iaxhvm75fz0J73tWtk6aY/dP3XxdlE
WsfdPBmG/3PejNX37ELieAehZKBJU6L8VGwLbWInfjgRToEpLvUcxOzxaLhhwttGoNBqcdSgG5sa
RsIPlzzFvOKJSloy6vCJWbSB31J7GaG1Apr8mLMtXcaiBBg1SBgiGO+3BNbMy3BVUNXqQWTacDB+
TAxR6HXRNAOQGbuBIgL/ZmcLyvQd3j3XVpmb/fO8akfK0oA3YDUs7nq7T82hua4lRzjy7RaL+7aI
mzndpaPq+QJTMJLF0Cdf9KA3CJvAFn3kZKHP98FHikMYsnnUgpj5hfpjEab7Hth4a/t6Q1KSiCBU
djoXUyQUizFX4UIHXjer287P7FRNm1R5Zftm8+swxF5u/dVq8DdYLeAc0k8R4Ow3VanFS0cMNI7z
tn67xN/qZGB0Bm2TDeMamn0c3g5eBg/y5zGE6/XL8GG0uRlTQxAkovUaV6qthYsXFKwsX96arDUA
YeLj49/CCawA2b7BG1iLBz2O3lvgGQ8zo1sZNHCyWPln9ylg1bLP2Dss4SCzqGnIw/Zm/bt3dg6c
kIECxdSQtQBR1eQOLVertRdz1opbG6VNIuAEEgapAYUM5HLftiJQtfilx6Id97ProbPu8O5XfLPW
YDwjCezPmjjNM0eKLrfPzZD0+p9BSsaxedwTwVOw4tm8/x3fE3Cjno1rKgIq3lXVq1/P8hiPMFXT
xe3VSTK9OZifOv6J/lg7aa9tjpdIl38bnt9wZInaIsNkBTnJhpf0ppOT6f53Ci/h++yC1hoAQWqv
UUfAMw7TxrakjdSRplDcSkMdyHpXT4Mae+gpp+rozbDaadEqhoxGxUyrgLuQS0ylwQrQQI7s6uJ/
zrqsWuqWO5Who7sjXEd2ZB3T2cd2QcZUxXQhuuNYQBZSDd5zMkrvkoDOaPX1ql4MGpUS/xXAw7YL
naD+MII2OctT00PgZA2XAq/W+2nAEuaGquPQkzx3euG9cnI4NSym+8RD+iD7kwTyBwxXvK/7E9mR
2U7DKJI5XecW5Mvz30EnDaXtCRxI0rDtTnDvFMrUC4EfEoSQeKD93bAH2ysgnkF2qVk1lzGhlaQN
PLS9Xmm2J0Dy++EdQsU9PX2asrzn10GtiKsaSMWKoPlILcqPbK6ZudaqvGjDv33+Ex5RBeSyRSVk
ORgWNO33+2P60Nla1qihYqsb6wzmtbvFsaeWIG4saEhWxrFsW+0I+eXWjbaIvOIjpbNIkz0EJsIE
mKPsh36jZrXpepZUm4QCEGCa4NvLbm8jdMJjbcMZMgod995vX+mzwzccAcclbiJysIwamORHCx2s
H1sTUjtobhkexFBHdS0xSHrVumXT82Xu7mg7wAwq5UFCkIxsP5RufQj1WImAmshXBNQSV82hqaC1
SEn3IyUav4eUo7ML1YDq4BErwW9GAWEwVvumbwWcYFJU41azGHfBGmXv+4UjzC2KQBRdM7n7mvUU
ojsgGP9XF0n3ruTqjg6F1LLv44MeiAhD/rPa6/r5DaXZDwSyY2MncL55A4ErAGfg7K71Jqr788uR
/2Zo5srSW6xTIcL/xkGyALgpdA+PNjlGAZhEGIrfUdYwPKN3XiN7ryURpJ+fxDpr9PgHVYVkOHxE
7HH5ZVB8lltcF1iYIblcoFpXpCrRNN2CL9gk2zLM93y+jESlXzQtsxq2IeO3iq50zsXaZf1v5JZv
7f9MrXSWOsGAfzKBeqhODQqDEXv0hxY3gmK8ztH/pHwSK/75LkY74B2Q3YGpUag6E1hRgdCDG3Gz
u69RvL0J59yYm0gH6Q6eSOTNrBlzs2sv2L0WRNb9HT2G20yvn7hpkogRQ9OY1fNKGUf9WSr2Ex/N
HPP9ZD5uRKiyEKsr+xJL5N9kM9Gnd7vuy4+1p+RDBEgD/dg63B48oZqlZgxN+YRnXE0qMTFkCMsy
GBeRObfyUCVxnqEcULH7A15m9p/iXDWB5khI8QBYuKTNjJLIsu3KNkDwR1k7vjU9yyi6lMHV/iID
IlBVp5B6Ut5bgHLP1CzIAaFJAofAK3Hh/9XdHbVLKa3mU3QSE89sL0ZyPsTD5xBNGrv/T6qc1u0W
ylwVIG4gHdG7l1jeGIZe0Acxzs/y9mrWz5AK2me1Eb62j7BMpysR64Xic4znkyAzuD9YeeIiS2Ou
RNDd/XD9Err7hBT5KwW1dbCUpbJtraDlXCrOBn2pOHdoBJaE6sF1vcvTCWxiR6OMs+6DqAfc9TCB
kVDU7Zt9lqEeepdDbYNeWktJAfs3r0duY0RC6qtjTFnsxpxekl/qyVhdGUFs5q7EmdgcFAKe3vJE
smuXiGt+uW1XOrNb7GQSo4CWwE16zat7GgNqkE92r8dtuGTDpWjAbml066sPbvSfnL4JsehywtmT
HQzSsOo7BGDz8x0K00rUj5IaQxvjnMBlOUCHrcoKAqVkANjGSD7toc+fwk9USfbGVrKhNVsYt0YB
SYGQZAO72YTRcsQYAJiVC16T+zmTBCjw4z3PFGL61iZb1DiewvGZsRpAfCkjLiCrxnC/hSA+nUpj
NyfqLmRTCCOELqdIBhodEuWJgmP+nNKgjIq0pYbqfFJHunuCXnIdbbD9LnakhvIAQ5zO/dV37PS9
0xd+hBNjk3FZTCYDOPaJ8EUAE7jrBHzTiZwmzb9SFROVCo8GFz8Ka88X6BSznBPMUDYfxnt7wwu7
dJabfAbK3KnLrNSAi3XruqEUtocNdUfv9Ftu0Pe6JMQxnEKm8W630sngFZF347sAgQCYnwaalW7x
I+QAFj11mma6/tR7h0DvjPva2vFLivj+TJurEjvGHT/pV71TKKmB6VIZTRnJHPOE2V/ffjBcQsM6
a89M+BnX8dQfv7eUD/GtxEYG8dsd+vPuNJMpIGCOFmqDJQ7LWPjnmhz91lwUlYfVH7IwHWBk9y3g
PFc3UeCOAi2KlbcqZ3IIjjn7Uo/dtOPxYi7t3iaUp/B9HQ5scsMT/n1yjaqsVQvmUfWW8Xn6GsHE
SI/VbNxoEzkEy7+tRD+7GfP8tgybSr6tAJR4GPWhnZQ+uWq/XPq/JOwh/kLNay9LSEq5z1vVeRJ2
qzm3FPG4SSu6P3QppE6A0fHW0rHYwZRkVUIvkgfLiSLyFVywyFUDO1sEvI0CGX+X1tkX+vGasx0n
57bN2/R8yEJe++nfybvMiip2DqEM42k9k6ZDakWsATPGbpQwQOCTbXzVMCcw/U34GOZpEh9b/NsS
8a0Yhtsx3tgdichYy9p7NIBi+MN85JizfgtVe6UudlZ6ZY7nuRa/ypoo7Qe4wVjb15c/lFNGdyxR
dOsBYSj28SCoJy4j3jRNga+tR1gH8XSRpxW2Bs6RgCLLJ28W52JbtFNcxk/TbhqULDGHivB8kclC
GnkDWxHzzQQ31FKled6wix7IAlsy3hd21NltXlIAniGc8NKHGs7CCOoklSDwzuYSAO6vyrSxNHWE
Y9RZyOxuQGcNbsu2uJRe2CYSKiu7USUN5NsgtvA4csPVMMAuD+atzQnweNRZcs/SXjv0cy7L40s8
elO3Fxm3OzLSG1LphxZ/6fc+/diSj02ff8eB6Bno9fNg8rZKPKo9833iSOpCoZOGj978N5idH0tB
h31un6reTkAV50zWpuAJW0SHYA5T4gCL1HZyYJQDJt6J4uDBrcFGEhv23oDBUSt262K5bXqpLte9
Lttfjjx+2EqCiTLawnOnTFKJaFcpmDZ3xdqHMhYDCo0M7BktxJZf5XwFm0KpDrMQkoUWJ00rzi7A
JlqOUTj62ApM/acWRSERKSvZyIEwNBOdZb678hWuv8h5kTtkZaEXwuRaJHSRfPMZv+TrYSs3geGJ
jRFAMaRkBYJdC/nwo3HVb2MzYWWPbxCjKOy2g9W1O+8C+x93TG4frkkvogtBqIhzOyiE4PtIHvKY
K3xQD+3tCQR+0Y6SOG1M1Ltx5IHY9YCQJuDjad6vMpBHsopm+XoYNT7hZaLS4dcoNz6O1oQs77dT
24yNGpMZ6m03gveiF4rFUHGGnELk0YrDiQu1KJTouEbNZsMziJixxv13PNCkBC8eEI2Kkhqp9CIV
KeMxfeVLJZRGrn733RXBlvOIIl/uR7pKcXDXPlblb125emhY+YYuCuwCT+Y3gtwmqUbBe7IjWeG4
h2fijfB7orxXhZYO/COGiEH5KnMUhGY/xFeaiddSmo4ikACtWpYzo5oEj8YbN2/xSCnYid1ZYx/z
3uLLus7c7xTbkGkn5P0SK62p+zddoYvDY7Xgime1M9Yq2dT5fzPGzDpby8CPtrLtct1yvj0gNgod
Uo4W7YDPs4S18Mvfe6Tgg7by7w6PYzZ+km0KYFSw1n5dgYxZzmOWVX/3gBnr+9QtpZvqP8WdLqJx
WMG/8NmDUiGSaRpf7P7swpz1O+fP0xdxs8if14i0LVcojag54O7CL2B83XFLp3qFvx9/+Ji+UQ+P
s3ug1NUBKgZpGRVhu0icjWgSLlds279cZbFRP0gbJm4WSR3D3IfvHzJXGJ0bsHXxTf00PJqKTYfh
tOPQzm2pk59PaUTyGuI/Bdn1I19/ljW5AH134cLwH8hbOqavztIhn6pmZthD+VSiy+z+bHYUZFRE
faNO3tPpr95Ml+cCgcp4DdYd/XiduNZGIz358/XVVo2FVW0XzglOdDnxZWKdYPpFWrz2CqR3OcQt
0deahGsURHU7B0vE3EZ5D2dphPHKtHccFeH3MgmxA7vsPSrwJ5hsK3mzfZgRrKnOUxLyRyhxcATx
1TPZSwn9Ogur5qwvW+UhhVro/ZPKvXArQi3hKNi5F774+NQ9FwUPEg5oPfuVBZ0PVsIQx52gtq3o
Fg3xqxtUJ5U5r7A1DP8NN4E0h5HYcPymk1BaHfOplR44nnxOgatQ5ZXD3hhCQhY50PhsCRWD+zHN
j5p9sirLu0NmaM5VvyeOS/dXU6Hk6s5PK52fkrwpWBiQ03OtZ9UHARgSMbWYPu/3us7Z/+BICgBw
wouRIwHy8mZZwMPLyomH134XIHGLAzMIB4j9QUzIDqFixuB+6G1LVJjRVva4Og6ZVOp40GyByx/N
s43xHb0MEkZ32KxesVNCGDjMThMs9dtBtjyT2+mNroFR4x4Nu5LvEo+wKHKli1b9rzSSzsFgC2Vr
uuxr4rHdna5n2/3LSgOvL0Ax9ZPBCXYHDEU+Xt8eF6FV/Xt+l60H3kznXSO3FRrh/nNZTYGbB+sd
/RUCqlDCzI9F69Dz2mM0lh6XFDB3+cQjlo2SH+SbaKjFEiNDox+cyIRDB3S/Y/DKdCRdJ7Rbvnib
RJIGjcOvECi5VN+lRr6sza55cGyL5mCmYmdlYFcwfNZFLo+0+vq6qyuAzafS8Ct1HXK2nLJTKBRI
P2iZ/89yqiuISYM3sl9w31r7s3Vln63diBvWdpgCYxiwRF6zkEd1u18I3iZIK0NzDUoJoDFIkBhk
/LAjdVLIIwKZGGyHqxk45V0Ix+FmroHV53rT3+5i0Exh965QxeUCLUZTxBsYGn3xm+9Aat4QhQAd
a4oBbuEGGx2EBXeplZImMD9F6FkHPHz+umHGrYrDCqwsEhKRcUeSkrFHXkQQejQmiUGBRZqdtdzl
K6GOO4siU5DkyKn33MsYqriBh9Wyhvh0PKB2h5Wy2au5EVDDSJcqQuj5BwG33Aj87u70ETP9G5Yd
nV32nMwuimeGAlF13AkQEXkc5Sw6Nk+o6Jme2GL+0oB91rQA2erYZJW5SSl5l40sj2ZCHm10QvRB
QtUsrxegcpYTDtlzQwLgMgmE66sgCVpG+W2aqS7zZqjjEfds1P1GQRjuXp0Mb0k0pSydcKm4V/PD
3+gUB7Gzg7ijNg1ZGsV40gMjt3VL5l1y+t4SJqhsr380YOpEfqKTt4WcM1LMRThxAKeZDiMqqsDD
briT7XLFNq6Gqnd5gebsGzTy2it3yDr9GntPnqR8kqXDTYmh5GTjDMDsISABcq0pe1iOLrcjy6aU
XVuprm3EJ1+x/bi9zo7402Mry1XbIKe/459QszYJZiA/gS8KOQvOCaVla9Oyhi55nJUBQf1tUkMV
D2h79PbR6m3lLW248tNKIyb5/2YoULCrDECl1CpkHnErjAjI1YiDWTW0GfRhX18sQCcn01LG7xdp
yEZijL0efivJx982/c+K+ZTyq3yRFpZyiVOUCaUVXerxlaIhjf7KxGyugiSu+KEN618n4yxv7pus
FVpUIa/h+X6YTza3rr24EK6TYw4F5eodTfNQW0/cIr99cKqyudemNez02X6ujcDr/L/C57xVI1Pl
I09KY7jyVFM7JUWV5fDHE1Dk2ibKVLnEwEQqXBKHAJlVwIOZ4jLJbySfsJYmClCGYwKr1HyRzS2M
6zw3/l8iqXkMYYEEORhT3DaqgSKNOtnEojnx4/9FsGbXeL0KiJi7OfgddnAjwHVmE3r7Ahddbm0a
2XVk1Xir7UJc8bCMp4Hl6Ya+t+4UnBOANuh8eKmcthsNym96697/fxphi6rjXiR7yxWWqtSCFYsk
EM+3U4RDojvAnKNscFBDp/by62DLc4C9yz0cYjFqLoSqXUEgk5MlTgwYgvQz9frqq2CO/6DTfLRs
fmGxdiaJhkdGVZk1ENaprnpP/KF/bzOxwnjZbvH02cqYijw0kpi2yqnKI3eHMxI5FwvlMTHUPFir
Oe6Q0jdwf129nOboZ8/D+9LPSdpydD+0nL6MOncvhGpns/HlxPg+DBwV3SjrPF7V6NjI+DxaYBsu
37A61lwEyH47b3gPegpdgY7kRewNzd1aBbEiAg6qfoZ2eRndQYLWnMfe3NQC5V0RZjeJhQy62+06
5qBw4T5pszGrZmXIIBMS1utwFIuUuk/Jv4N9R1CRsXk1sgIt/5RSU1QsytByYmLhS/KSqhSV0CS7
AQThf15MMLM094hb4drY+E4os0V4fOnhji2X848AvwzNT2BfUhda0XR8V+uchgX17VkmgovCudY8
1atlY8gufk16uwj5CpE4QfUCSaU9W1cFFE5QPeoLKQFBVI9kuVEkrAXbZg+xr3pN2HvOp8DpzZsO
W+M99X7IttdCrvl3i48sErKlNx4s+vu+KAwJo+mn9yEuui/qTCwV5PnfBI9f50tPzX8nSUPAYprL
k8gKEOakwBW0vzm2HhmI5qjVGSB77XxspTZWT6xNx9TLkEjsk0A0sqGajZbhWhtcg4CRvtaMLwl+
8fgrjwjZK3yRa6JAIhduZzBBiHDfwEqSeXOtoPJ1WJ0Po/FbyPOhFk4lAlP1OrKMgHld9CyKAnvB
/41ucgZ/aEHExJptY9Dyhbezfx7KtvhuVQWRD/ZiDFCwdRciCoVnZGYGP9q4w99/iyrJz0rqrfDz
CtakrFl+hfRQFl3mDyh0EdhQLXctxW7BToTOQIWCsPEffBs9b9Q73BfkZTKgFiPtAg+tCYM7gYIx
5XfKQINBXCLvrouAtP51Pl/xfP4pkg6RO083zKfNrMmU1E4afuXTPA28QzaujKARPDy++inrbVeB
YU4tmA1hHFbaMmuMV9K9O+V5b6psVIrv1Q74/b2WQgRzNBldCC5HPNVMBmmTIqK/Fb1RonQgriRb
9HUXiDkabw1cZ1Q4Tw04bGyok+LxvJeDueBcFXoo7kKFdwqnH5hpJ3GDyrLRczmbm5bsU1UDXsGC
09fEJxCa8i7G0H6Dt/Afakl3sM18Bw75fEvmOSAJkzeGtoeqrb+oCHWhG2XGQi+wQwefjuibo5pu
5oVuUZ1rZPa+b8RUe85DKg6tcIZuttEJj6HwxB36aqx+u/QVrUt3hXe2xECCSiSwIk56kXQ2NhIC
ZHnKRHDHweJzdLX+FEZMNHYNauZ6h6EOqZAxuCJXrXCE4fOBnQHrGpT5lvYmvjjp0ne77hTyIn3q
OXV4HheR1/3KV2LHuKdi2+iU3IGe/xL6ygdu2WLzEj+OUzUYjCuOINcc0/+B+vNI30IhSnqtIJsI
VZcplglY44yHW7h3gr8M2F/DO/kGEysUW3+z44uxyZ1T/ObDgNVF8afS207pbWMGedEK/2xuMR/g
WPfaQqCk9ae+VbqNw/OjEqrJKihMVeShP5q4gikPzgRnP8rwz6RnzBq+AkJD1R5pRh481I8r5ksx
RaiB44+AQijQBFLFSfJmmyHUCJHkoQ60bpWsJb891sm+o5tEZYjRJQdoxSd8u5OtEkI8AKF5Ji9c
GJXINQtJbK0I4l0iGyMMlk3+Dh8p/Oqq/yz9NMRKwgf4fXsanK31gZclQcLmCaHOYykzd0zE+HhJ
Pl8aisXARFiaTN95Ne6cS17b+DCoRhrSe5HxB1Bym/xsGgLTPo6TUhc9AseiL9dCdEcEW82RJMbf
5RKzMr1DtISh/J4xp4Ck1jX+OA/FpPYKraEFHQxOtU9Qggq1NXlH/bfKzeCIfPAMTdqZkm4VMRWK
ITr2YZgONAoi/PJx5t3OngKoQFnGfeN8hpQHwyQpYRG6t6iRiz4+t8pmzo5/54M8cl12HWMY8Zq7
p73jGwJ/B9x1ZIRmNUq0+qBVknIrfAA30I4BUmZcCs6ecB8eWW8TUir2bfRVLyHqAgzKvnAY4rWj
axu+DBqyDLjJKs8aFQeYxvZ/cmlqMUHTrr3OElVRfAFIB3jVjerGrhfjC/kfL9JimpOrWzpSZ/Xt
gAQ1FItRFoJ1bJfsrAi67wmnHD9hYvdWJqMgiNc9VEEtjA5BAY3QqDwJqV/WYtLXP1TwOufPia9Q
KM7lZOFKxoyWqEljy86LBiTQtlYP4x8fsRA+HsWCBT3/idql81Cudfz6A85uNjkJWKlDI93fSqDH
O/Guce1ZRsZpI3GimU6QqN91Au43+evIchi54P0RLjvRbc+ga6yU/B4cezzjTCCbvchuA5N6T4JS
WmxcJJ8BIw+qbduTE+h8fiCFry3UbB82ODXornzjbcCAPcTK+ytzBRIc/WP6jild4rLj4e8BHoiQ
2ywAkVO+u+qsVK/R/5GXTcHDf9CO6Pj9sFkRzy4JroTYtThAlM+cTzmKoeYqbpqej33TBAR1rLLI
FTW8/ztyZ4a4lYi5Y9RUXS4zSCN5iGrkqcEE1bMIvLBGnAeXNGgrITots4wwyhO/IS9zxg9KYJ+A
1zpfd8mHjiwL6KBk1rzqFGDl0uJI9fTLEgjnYFS9tsW/fm1HoCllm7r6HIv9IVb2qtkkGwKJPPnJ
j4Il3KHfLuNNW/MCeqv9VvcSfWvAeAXTd7MyWq+0N8bo6Esx9+7Z5odVxJyvmAEtETYSgq8gc+BU
hVQiQj8IQBaOpOIXbwPG/hiy9HHXJPAV+CCWFcn1So0atIng6ZWAzijf3+EZojwTkaP+O2Jp9Wk8
/zLKZV8LqzhkDVOuaHDe0k4VhDK9v5M9XYlwVuF4k/2q81OZbb9Ydvjvfzt1oL1nqXvu0nFukrlt
RIv5kxr7dTOp3426izgznivmrvZxksD4wj+NhcRtMbuHOjQOy920dkpRsr50VZsBRhE4lt2t7Dck
V38B3ncxjhwnEVCCxGEqkHuoJyQMeS4KZ7SpdE23tRLiTdHj3aByPwqKeXDbXBAiNQeGocaqP/5m
OYj1LJv6v6MxICgAIaHtiId7P+CMNj3UBEWb1PNKt9mRelrQ1km8yPNLImNoGqXIOux+xtAyifX4
aWSEhoEB1cssxc7Nq7dEm2V9jV0GEcGvpkM4joeWmOMS73T1h5KCJ6VdRXgP14ToJhZeToZh8K1n
EkdBe4pCtRh26zDnSk4Qb3T4D2R+S6/xqnfHPPSZrSj7RAqaJJ9cX6W5F4+cl7bzuTt6pq89BSSI
+m3MslLfSMMAQhkmbuNlq3G1B0GdK0bEEzpv4PHHbvyfp50ZqyifLYdkHj+VWcRZv8SDZEmXdCxZ
NFZz6l8HMXpEBXzrZplOO8kW5ycH6WH31vfhMeYZnYbew9JaLYp6BiTkP+ATMo7tKZulcR2oFRHf
AmD8oJlgXzNrBTBktGmxm5YosWsNxajYHaXXCM8rhwbAQWTjwuIxmXuD8/DctQWNVkdnkAsn+gdA
9xL+aRL2nNLWVxVEuHPD1nd6gW6CQAXVM5A7gQHV6D20RLpFxd7FK4vZw90S+XlyXDJtate4NFT3
xdG+CYCT/DDf27voPy/LLCxmjUz4teRvSEwzpUeAt7mcO6BDRx8tzB+30AZGLfQPEPCIankr13Oj
ZK9AS0yPLmrX/Yn3Huly8DurYef4QqyYKhU9QD8PTYkfdxkKfvKxQJS3NVIuh1gUFeS+/zY4pIxC
XHEYtwCZzp4yBQSUQgz0Yx6Pp/J8WB+4CJJqR2Lsgv3hsddxZXWNh5NiBO7FNkEyYCmm7qcIKqE2
i9s4uF4ERqdkQSOtWumYH7T9jXEzhcxj+A959VhAK0x+7Iji4T6DZUWZMJCzfrwMZWhYoy5oRJXK
768+1Nvrb0P+djJ2xa5lmpOe5aBIFHo6vaqDaBe53rwbVYeQOuxD8ge0wh6RlBPkDn+HMejmPzG9
4vTjoEcFqvDxzoLNcw7c9UCT9T1XTfCykrTfrU3pak+bf5CGwvZH5DBBi3zhQuU2I4YFmyzDhHNj
1S5qismfu8+MdUx76sa2QUDLSVYfnn9QTZUKbrEBH+8xr6COxjz7w7sxRJNC90LWdlreoTn/+d9T
YCHwy4B63q42rpDLEaggHevov2gLTHUzE4qdlSuj+S/mUdOfqHsxzu+HyF+RNAgbtgyQvMDpIlmy
txzxQuNXW4oKRF6emhCUMimVCEUa6J6QyRW79PNwxy5ZyN/X5/r7P1eB+XNxHkEQTx9EIvHZnGA1
wLEXQu78Hmur7jKG+mWrLv2TsprFWXR5goJbmVD5Q3NJhrOKZYT7Dyeex04SfiPADR3CkAScJD3v
Es/m6SskOcJo7UJ1kAUDFxYmmaec5GhUcap/VGyoFUdTZMRU32WrC3ptRM18lSc9RyTiNchIXiTb
CRAV+ZQP8fBLW8ywa/pGga8UQQSYWlljQUR6hz1WtPUW2AZzT6s58pvTEJyfyA2+OaVDdQWZebcN
wwjTXwJmdeWUlJaWzQEnhHB464GZ8C9waJjZihziySlbE2BoiJOqKb0yIroh16CjcxCydz7z6kkv
19UaaP5/ThFQg5rrlWPRSojnRm3RfUWstxSsddqNkaGZVMN6jOAqOW39TMI2DRvLFiQ/V1g5qBuV
R0/Qvt4626u10IAnfKA+BgazQeHsx8zLgr0ULKGKfeHLU5+lw5jZotyOMPGZSzPALlz0iQS/oeLb
KKTg19sL39q6PcBk4BV/u8xGM17wUqidv5etnp/hkRg+aRN38vhRvsB9HAk+0EO6MJnX0PUzNX5W
gRtTBwq4bIMzYPSylH7bsJJoDRSEQ3SVxwfRxJ9lEe/RiO7aMQYI5Tl439YJt+2l8zW/Olgy6aZS
5kpHLkc2BtbRoreE5PcNvWwaHxtCASzWOq54slbdHaSQpIDCM88hvBVLuf+9eiZzS9CgMT3qye+L
beHf6v4stV7XeglNbPj+svkiDUsk8oOsqxCFYezXV0EDJEgEDQL7fozUUzFfP9yqHZI73Qm6pp1j
u1+836hyeMXHY4qcSh0A+18hD819psBXJNE/IVK9P/7oIPgJPErxIX7ifTxU9sKdK1ZqGwVl7VcG
2eJMx91UAqefXcUpQR+CAOi57mdifX2tRsMWmPKwIHyuCTM5MYaAD07s3wpRbCL8wF4f/rZhubwz
IFZJTUk61Xrmo/yekjX/xQNTNUqYs1O9OeI/YVHnNjHGXT84pHgP/1eVE/Vi+f+xRDj5ilKZA3ot
NAYYVnqM1ydbAW1QPNvGBTM2wT6ikNQuVVhL6CmTCxCUhZ2gLI27QHUA5Gg2Fo5VaNI0ghgMSu0A
4ILEfap18+xlnKMdqnMfiQNAyYAI03Wvi+PaKmgNoYit8gHNA1u0yfAAk7+HxTIxkVg8H1t/X5mt
7WWXQr8IQ4te49qYB4cGOIh2MHYlAMCUDaR5cty/K/G0WjR7CjaTiqPKMp3ZfBeSSxEruZU7vEor
CZaIZe/zi+tSo7THWLIcHCuJrAdvENOGchyOqXps/HaU6oBZo1zQa5cOTRozCfzIy/Sr3Cd+eC2e
wOtd8CbAa3lYLxtSjgjzrlQAQhydndoWqjEnF+wRj4XwY/AsIMb+CQWk0fgB74AKOMozhQSn5I4O
9tm+3TZuXsjZIuQgl9PYqA8ySHqxSGrIyXmszn8yFfCfQ+dDJz0qm3s8sSOZzoJeZ2mPiRS/mAUI
eZnO0W+W9wo07R5k0FxP25XRpycTjPR4eI+rNSVrW/dFB89QdrbJh+zO9PIzRldQ4afDjvl3YSto
QTbB7GmzchVjb5vbUctyUuhIXla/hwmMm/JFwas+yE1u75L1U66neHb8dWg2p4PqZTBwfxqY03ke
pwo/u6y3n1f7zH3CpJ0vCvR9a3DrZFlnifMAl5QSV7xpt63i9ghtBUiPH3zIkbxxyfxK0HYqgmeY
NF/C1j2SLwk+D2nh7EypGpENvp2jilWN/kDKk/8LgtELWWUBLNLgp8qTD0a9vQxOMGEoHhxITiQP
OPHOAtXYWLbWRLUsg2pYza8SJU/ar/9btDFVzF/3B+fuxFjL5/fLSPTXKfTftx8Dk6DunewYkiDy
e/EbGF9L+NFDc3CudZaamDdgviOsbUfpXfXpL7RWVEYUiqUCPtyGBbKuWfOGj6OKzjlD/Y/QPkFg
ng+YsChuf+qL3fb9ggDtR2tIl3scz5Bmfvn96aWn0u1EbFAPAcTNdEXYrq2XunXyencb4Hzb9fOD
VokBZADFNu8bsf7PaBc4F9qcQDGZAmT+EA/F4m67d2t3cLLAYeI5Qar9WENB6QCsVHPGWoyRhs8L
7f61JLqpl6b6y8/27jiEKpEKvmR2anhp/Ub3TRLJ/lxOZEOfmly3x37QSz717kMVBBVfZWpY1L+7
f7sOBQWuymN/cH/Qb/TUerrqvDKzHQpTEu95oSPfyO5UqIY8m3LxXCsfwQNyRNn0k+0QKb49oly5
9GXJ5CaZl+5hMeV5+pRuavZ6PcvlZGiD/lyDm3KUxCl9EwocuvgFyvROMlqsQre3j8R/yiPj7WKp
TpWyNgygUONvRfw62TIP3LDAKIU6RIBF1RhGXp+i5y/D4AtM0/ZL+048Qbh4fP19Eq7o/C4CUw6I
GyzoC93ricWrhkSssHLXXLybbuSusmP261ylPq2iFERPStQ9EMThSmpzMCyZE+gSRi5kzk3QVe+x
eG/F7ywwCTYB0p/lykRFJIxopLqyOTTFvEuTsT/3bHNfhfx/i488wNN7kdFdA02TA9mjEXTmZsUV
w3lGhaCpgvwsnwiYpjGCK0k6u5xLNNEvVjU7wWgYVCyi/heFkI/rof585c+DubtL2qJWpZwQG5QW
i0nDBGelVTIjsKyA1jiZTyrJSPZFC0lee2iYFdCPu5wwmJaW51bvH93k0/mFyXqcr8Z7pnyPpFIn
asZHT0XMt991n4IlgqgtVaqUBiWlEozhXF2NjBi6NYGb6RR/XUB3Y5GGCei+zDPkC6il5iM8l/+D
OPtdSX3BBeBzTnrbInFyzFvAIP4EObETmp+AfnRvQEwMUfhHPwQ4i6GucKWyfk/brb2rIYtneUoP
6FzA3QKk0JPbvY8uJDPuHL90wZJlvCqbqTzTPV9JsZuGjtJrVW+nF3rI12naurRWTHSW4xECeK7s
KYjFeU5ZbvYc5qUBBLrEPgMrPc1esZ8eJg0fDbp9QQaIVIFllO48qRE+SZwgujsTGIyRmfRzJzkz
Kd3X8WHWvRtN9TbKssthoEb0fk+2p32oOiipvWqto3RguWliaMaSpf3SVdpM1wmirw/dzKLzhYAh
0w1cZlbndXo1tpgIyOMmGHHBpFajP3pE24zuGvN7ylZTXseD2ZukymWIRtuWiROZJk4M+YL2OiVD
IaC/2qXRERhhx8f8c61c1EEflEda9nG/K3sloajTwLIurcAgYsotG+zUuBNiJnsjMS/CqHWKn32c
o7ARzpCk16aRFgwuhALwBmC8gEAIRsCxN9tMTkTD0FcxOXaF3JpRdM0nCIRLFTjIyyzXIGYf9rgs
2JAXcEJgVj0EwiDMjJ7+jaPE3JjXyhDq6XscqEoPEFq6LryDBfsq9tzWCq1TbWWLI0Rxl2lQPhnC
1o+BZCWOf13Mxbb3aDvxPZL95zPxlNfi/kU5DhGKDMLh/el9pOKx5K+D2P/8ZDUql8685sAGIgsK
3ed4rc/DIiT+Fqqaco8atMaiTJHeiL9krBs8pn6tlDg5R4VowiEyi7y4Q0e3W2WQxNs5u1W5beWK
u8iAW6qYnNMvtebWxvgr3Mp0S9Guk3JoJdlYTVoGGKhy4Yznex0RnvgN8i9MWVZj0I6g936LO2rs
8sKhr9B4eNmzkYO0d7F9X6lhQ/oKpbbFTOcOyyRlJn1dLl25axFKnndRp1Pasbhw/rPtPXdMqITI
sbLM3AcNly7VHxPR8M9uOzirhOukeg1zJOVRG3c2geA8HbE/d8xRiI1XkhW0dkFICm62YlzXtkPC
KH0USUX9Ys+gFQPV0+SJyZbhhhKDTqOM87teyMiYAKGgZ5p5XIebpP5FQX1NYb6WJsOXJxmlzOMb
If0bPe18nMYXQFjqeYsz/xwA5/9/pBeTaQzAGy0ibkFhQo65xOnemaaoC5g185QA7cyctHSmv3Cv
Z5zF7QWo7xY6OrhhKRyHYQ+rXLC74CS/hiwUR0S8e214XJQBQQClCVGNxLRuG5CH9y6SkDq7DgtX
KOcgFezpQP/1nG2KSSFauTutFwpTpG2yM6XA8Isum1Ac96jdkOgXfk+EctYmpowHU8ID21IymnOr
CcgAZDIvSysNOaOqaUVZTeWcQq04bLELQkUuWtjB4y7mxtnu0QikFr1eAS5o0AlBOZuluWy92YsE
DOGe802dfLYPfuzUvywo2RBAmuJgFCXearE/IW09zqpYqQcsGvWncy2HOcMbn5j7jnvRNfwWRODw
lqHu61D9HoSMAPUb+SiCNAYR+xZoCGuSnZyW/Th2octze8bbxAzbvnzBJ7yvov5JTs9un2YeKiDp
CkvgFNyOQ1RwPHoA1FjXEpwjsSvxRGK2V0uGznefgDByGdVdoppb6y5MxqHowV8Ug1hRJ1ajRPEx
8wwoLmmgRw0ppk3qGCxBN1KndxN/LdUHl5TOmKJuggku7rpxium/6yPyRmWO3IPN6TXwLjAVQR3a
F9gCOxIjWkcGG5lPPkmLtQ6Gfr3ZseGCTFc9BbWzAM+opkN3ShloHxLW8oHXpnfgEb99+pd9xg5P
g+Q86CzU0c0CmWP3UxNrGhw+BY+y1JIhpVzl5x7kyYMHkuyJLQUupDyLPywNboOq/8ajVuKFLTt5
OT1uu2o3GaMFkxJS+9RQjAbgj2AMHADdOtso/NyOVoIM5o01YoZnaxZIaMLjuUnC5Yp4V0mbuwKi
jPzHqqNabrUcMUhdJFPbJm7UpNkJW77y128yT0XwZrq6gtpSsRM6+BJhLoWZt5U9ZI/bOY73ly/e
Kyal51s0ky7H7fhYqgjDE9MWYRYkmYnFm+/mTPdm0KfFvnaI3b6K4voos5ae/YK4yluVuMss35vD
RPmEA/ymBOZIR0jxmXnL4YEPCwpEcUR+7nFEAWJbu/OXnBfZZBIpEIIc/R7HeefnAb8fdBLF+icM
eKBle1qjZ8kcWj5TFCswOCXmAUCdK7S/+2ypJZahpGqUWKrpkJHd0b2kd7pxWjUM2ZAeb2rwvgSS
IE/9PDJH15sgYEZFNDulWcx+fpB/LtdWxNlm1qkdp70qSeb9cvSqbVnZMWI7wY70aDTweTfk8Yae
kA9AbEWj4RgV3mEpMI/OJ06LhKPF4ciEJ5jPq+/jPSx2OLva512kUU5/cQJtlJG55GzxWji5/96a
Y7/9CdCZHuHdazIcy81H0f3PKC6dd1iMN36iHxHe2ajjUz0c5u+kxNVn1IaUV5VotuzF68XAKSwG
xgIrLSUIYF7KMdzYxG7ao2Dc1JaATBjMk+4luxN6RV0xcD2NacZo1zEv0JxCrh2UwEeBGYjc1zpE
nFJl3/RHx/mqmrnGwiWv4Ipgo7gcV9ZA+WPu6OH1ResK6BRFvcKoI3Nzs98ebf3tpGnUj3rWCYr1
VeiW8cn8oGZiwliCLsQZsojZQQH52HtFmGyy+xQO5hTwgKbGP29SLNe5/loSq2yf6m2PMQFAWF4T
HV95dgvZUXV7sNnBY0vi4I7yoRDAAd/Jb0R3LP2n0wmG9CiPiXmEHTYIPf6U2v/si3Cm2KCPsNCM
ZxdIRVIK0SzZZcnGPo3WDB5Vywu0ClQHfCqDx4vpOiUCidp7amJUbaVNqPsW1DxfST6ZCZLYvidq
441nUxzCbmZqoj9AmWps4tGBdkiEs/C86VVACgv6MPRNes8p6H7yXj94eAQ/e1ReTn6h82xdpJlW
zJFGsJGUyqmyf4xNavkzC6MONXjQd26OBRzr4dGhLBtHzGfdW1GcgdPkuf7MA6z+5VQm3n/y296r
mynhvypIJ5xdodQ3t2GETRpbMBTP49tRMbuCujUgsCx/UHV1MKHCNhA7qQ7G7MVsoaUPyrsw4vUA
qgZU6FagtCwd5FOSBDjYrjGxVkwhvO4UKNEx6GppFCYkexZQOeRHJrU47ccAyVKtzn34HRIMrXVa
gHyvEftT4/p49mIGevBpcAvMRjr83Y9HsdHYOHPQHyPPkIuSTSCrQtiqQDcnZluRArCX0Ckvuqdv
IBVAFP3kQB/stYZ7qH7dUBk5BKxVfcj6steiC7vbLT2PaCNxCmOlh4EVzdnqSLrhOQVQL0ztJBDC
fuIhaqE2+Asic2v6nqgXoEmUybS2EWO9Sl7XzGcbWXGYmXK98q+Af9AbrMBCZ2WGo/vKy/WpesE2
rYQbP3bQHa0nv4gz81PMYk03gmm4UsdtDVYmfvkM49kwOQnloQgP9JdDu4Q0wUrYqi82aHATPZad
hO8QNYYWSaIcR3j5TWIeD9e7F3Smpi2/znrffP96gjmnQIoSXJ8l6lbvUdcxRG7Twiv9XmvEbR+i
xq97TF5uyEsT3lY1FD4YVx+KhGGSx5MwnxvXKgBSl3lvCbYWtNZb5eJFiRLnJMQg40U+K1nqgghM
VqBkSsnD4440Mww6QFM2rl275GqL9GDCAuXHCU5E5zlkRcN9f5WAH5wE4Oq4hhucC8YSrZbyrOyU
VbpzUdkFaUhJCOY4dznpPYNfVEXMP0C7T9hK71gSu+dzS71GzEbCY0Ru4PK+DdMW75FtE7d0nlnr
xx7VjRqUzbW20wGctXbXkuAGz1qtJakhib2kVvPbOAcDDGxr+qUP2LhVV8poxzgX1WDZMada8YWL
LSIUJy3Bt6gYK+e8ouPHFdoHnftuNd6LFbT/hztcANFNxaFVJJtyuZVHvyJnQ/EZEyMavGGuOFxc
MVvLLC4iw/ZHr+oRJq5cRYjYeggC04If34lqFQo8+F+PlWi6vQVY4TUIx713OfPFLdot7enuNIa9
djE7CKde8HBMeIQ74dexRbkIE+mVQF+pjIhcn1GYIiKPZpxLIVGFITUfcfjBpFhUr+LkwPhaZ4c4
BCPXAUrrDPVk1qcR/9cQHScVFJF0VVyWvISeHDcNCvPfGJxJPvhlMpG1IU+qs1MpgKxF5Xng7fQW
iJpIEMkMrqyhbHZ647LJc10AzNE8XzOBaaa9NeGLx+ksl44KcZ79KXTBywj4Yz0wGnWjSBqp2+sw
568IsnmF5ibqhFCLuBd/uSTiXQxV7r9dYR4YKuq8mVK0pvIQ8tMD41Gi0h1n8BQu+SjN5yejSIKq
5W6syCkB6SIzO89XK3ykyYyGCna2Y+lwXjv5Xlee6WYrYThCDyZ4MWZVrqfiy7GR+CQCq5le7d03
AmKQob/QjI8e/9TOYZf5PV4Yh+ZsFM2CBmtHa1oLLUX0JUbLx73DzM/bSnF9gMFYad+W/4KSL2Nv
MChTX5VLqJAMu8ZFoBIs+4KAfmGopygjH2U8fktqzHU44qNaML86/5+tv+m3sgjUF8P7yrYZSAxy
MOCGnRtptPn+NeGwD2St7HcTiOUC+2U1ehQgkuNxCgSxgNs6vomLaqh3jdhnIk8RtiU1bpvbW/FG
Vy3hlBsY7Tayvoe3NxmzmAcM5+PCBl7Q/bXpxADrKe5B9tDtoqoJTkVwx6GSZnbW7Qq2QnPlpA3c
z6z82tC4sSd46dMYqqYcUCvF98OtJSfMSO9Zv8VqxBCka3LFfffuzImOevwF+aftYheuRwZw/IqT
/3rf9AwUlGOGAb8bzTmBHdHspA/f8Ieaje0DbOfIPmaKt1/lzrWbyl1jl6uYTMIuO99RDkVvglwn
nlrWNqTd15NGKWD5jmALvBENVNfv8xjLo0Ndc40otb+wHbo8KhACG2LJSK6IC2iT7FiruwylC/mj
LRIM6FgJQSBqvPBySgISFiklR0GrHGMsBsp/kjrNB6ECi5I6nXlUzEZpX2D/5w0NNpowRrm5dyWS
fLTnR2D3p77IwCpVk4G7byNjot8S3xHuBZ/+g5uI81CL8ExY97lNDKfcFBZ13/KTCz8UHF/ZkUbG
LwcL9WP19Wf32wuz8zwGv5WoH9nS6lxyG7fXPS7lOym5yQJBUzDoOsbDwljf2xj2pWghoVFqU67a
ne0erqZKRqBWPDbGXPMa6T1n85swBmMKNllVPhmgDQwn6YH5CL82JFklMr+ha4v9h10BLahmxuAy
6cmR2BbbtATSRTmGo3xQQTXc2q1sOe+OvmHHobsHyFE08Ne9X355PQFJZJ14fbqRjkSgUADALmqH
P9IChbBSCdTKzUbkTE77xYP4Dz0iu9FW4AtnFPu/okspVaeNflPn9WK4PhytgTb1hF6BJj+OELKQ
BBvB5N5c6Fx31l0MJIuak5lCfE3UfCkP+b8U4U8ceaxn7qwpNlSdFyZbUtlmXeh1QlJqIobOs8XJ
Nya18cf+jYic0UXZpXYH2FtrGGcXQo4gxnf5syP2jO7hr8FUWLQs0moDSVGZAmeRKB3ZngUcSWmJ
yYcJOnhoDhafegIUbdKP7owtmYtSqtAeerpTBhucEBKomXsrmtziovDIHl7qLYh3FCMyQmKSsFqI
R4mAhyoKMYfewUB6FuI7O/pJBiCRD51YIV7h89KX6EWO9buUAx9xdlEjw4qyeSsDwynWhz3bfWxO
atJTOZEqPk1p2spqINpW+QK2T9JHZclMgWwQFqJfKRsuV2ho8rrx2M5SNesR7yGdO78w0FWNCVS4
/VR9F1fXQkUj7KTsl2I2morHHiyagW13Wwko28qarAcpgl2Kg6JqWUKS8SFmZIjUeJ95kX1a1Pjg
RE+rLZN37wpboAcwin1TM28cXrGRD00kUDw3s7vui3K1qnwz9wpZbb0EbqMAEe1hzyHvxrKA3CGw
Bd8Si3R7gp8i2mDCxWQREDdniIi3lf1L56FRU50szeBsaC/t5NgYrwDX339vbTIQJFRUpG2gLlZz
XnZ2yCl/EbknRHvkg7OOkfcL7fXWZ9hGlW0AVBrNO/6co/qDeV7WkRnthIBVIkppI8Rkyt5CNY+x
leGQdJsnVUj8Oxm+RVrPoeDooFxcxQx+QHI5ydbVQ6PajjxV6kpBLDbj1o+OcMwY4P45ddUWWRar
nHpaoK9yMIHZhDii1dCd31/O9H1dCWbZNU6A0Wxrp0OfilBOvSBpMoCQzbtK2w0+3MunMxl6u05s
yPQ6GYdOb0SnW4W6/rcxOFESHNgUm+PdeaUv6Z1S70WHndqEmVsb53AC71QaepHFRv8BssVG8mbX
izfY0JKI4L3pmpoA6wCganVh9/8BoLkvL/NywwiAAasMa+E7Dm/ohw0OsK2jO2qD1cXkAOZwG9xM
ULU1fqhVQ83qoMGY0cwnFu3IBdGRmU484w1cGzJQ1mjtryvnVE6ZHkRI2KCd7JgUx9ROQ6ENNWcR
9XxASZYJVE2JEefNiisBhiUhyJVWY5yincVZbkDZhd4HkwsYPXGgDbioaUlMHUk0ybV373O86UoH
K+j02+rw04N259nbr8HD48FMKbGGf7EkvZF8gt46aQcYL42RZy/cLEnlm9gOA0Sw/o4vCES1wuzk
DTOQac+zv01jFDo3J4JfZJSm3gNLV+SosySPtsEuZxsWR9N22BtQvuRMt/vDQd3HqjtcozxP4v1Z
DJ11nNrGsbnoZoiv/vOvHnOF97uLvwkyLBmjzMRV7PqSFiY3itj/Opg8Zr8lrpMwRziLP16FE194
Q+MCgF9v8BlqbXIwJda8E6qm4Cz5LwAOPASYCQQxyMKx22TLAtFV/HU2kPUOWMVHskoXD4wuzbzy
2xJEyxDfHnUnRnb4IL95SPvQidGFqC487LD/oKtMqIyftTUoB+F5sJ6PUUrXxBLFCWqsbCrJ12dL
PujnphWaorAyPHYn48yeD2oLEZL0IIj2v3s9y6IxnAfhrxCDc0MwcDy9x5aT4ZYZpboUdjWCOAJo
+q7IKAwjQHRBv50YYfsCa0nGFeL3Pm/cGsSGE2UHissLaodqq0yplCKun8zrtKZ9bFv/iQ2yaDba
iASn7G1nQaAkenPIVKbqRN/zoOS0yr45tMpDoND9NHy53r9hSbkHo6itDmcZ/Ov6sbMU+A80ZSLb
DY8ArKtBi8aog9yrxY6bWdAKIqsvxA+FBJoCxBP+mr2PWuxcGsllAA6b7W4IpXM7rFIS4Bqi4VMu
ii8DH8SzAmYEaTLVdrsAHw0Pv9cswjjf6VefOAO3wbpINr2JHJMJ67o3L9SHhAqgFiZ/qr73KGXe
0CNpG7G10MAtFN8RH5fi4fx9ytDQQmVE2pV487/ggvAL7vnUHQK7wZ27B9/hWVyAAUW1YT2mynjs
iTe13vJE/rxBl3O62t7D0lQ77k8yxtEdQhnCvzt1xwgmlyp9TcWitNriz8MvQ0N/Bzn3bIAHe7c4
08Fyppmvrgr6ppcLOza1I8Sw1ZLQqpayC33cyHPG6XQQOUODWOMZ+E/ADzt3nZh+m65y92D3GNkG
2X2Nr4QplsIf4/N5tppLXXfWA6iXyVYgXEGcNzyZQrHzH3Y4LxSDQ+Iyz8mv4zJbhQIxcBzcibTN
Og21BPGjrllsts0svuQLWKOoPQjSte/UfI1o/nRJ01gDNgPXNfJSHK11+B2XXuEwffCM9U735+S3
BINHpH8dfwX/VSx7ULuEQjozym0TKcNFTntseRssVXzrtzXrFxFKMspZ3ru1n75PIfMpji9ZrKSq
v8X4dldwZ+AppGWWqRfIeZyoQCGKA8b64S3etYdHZVKw+oisGMlMcfiT9humQdDdxVGqqpu2Krqi
JFLml0hfHyUB1Gd/lqxs7pndMA39Oystj4aug8cBDeJ9V/6cB1IoavqUyXCYd+Ie0QNbhnfJtd5V
zMkon+wBnI4DLK7tmHlOhyWJtB5uzsGUOjaI6DPFEiHWVu1IBlF9IyI/7WoGRoEUBm7UK4wMnu/u
kRTuY6IL7bSDQuLHtjR4A7Yh8ueUVkxth+LOEq9NPe5gpfeJ5KoOzmLuiySNAYBsr1e0aidxrs/W
AjQRBcR/Epx6OvDQbWFbQIHagkDS3Ppp2eNiQdiCBiUes9wYfWsUSc7BCR4dvL/QZkTBXVE3NyE/
0EM/ILbTFBC+CVKhz39UdXcGJ7h5xjQENiZoBWt/5JYlsVPxjg8XH59NaiNr1q6sVShd/LJ3RoJ7
x+rEKeEO66LKoOikE6kD0zC1CXz4mmVNpu4wY/T8wR7INsssmmyRGC9U9DDwH8FuDn5PWeuqxKEJ
9T6v7CK1Z04guEN57UW5nSQ2+EihaskPvC5iLnnlqda33MiSjMkokf30xtaLqxXJGyb5FKP2Mv2e
hwxeaHDXPx0+rxAhwLUBGWz00dZkxECYefDWB/JTYemLsJrNtU26oFXFzQtYj9ZSNxoD0MRPF82i
5K3oB/3O+esm83xX31XokJrFSnTb0d9rmelYL8l15EbyUegvY7XnUbUCW6eLSOiqm8ttCrAlXnAM
p6FbwNKJW+wRhglMlGdbnorigqdN3NiLWmWRLrd/W1PIVZsopidZx4UjaLMufq7ePOB6PqubKvCd
jr36EA5/NG8PsyAZMACFOcwGLRqKLNtDv7P646BDMY2aG4JEqQ1AloyetljoJHSO95ZyekNBlWys
8+G2LcKabRekrtyM6bLQFtZMqFpvSL5CF9bA0tMnWB3cvLMu8VemblJ/8HUXS7pgEz2WAqbTYR7O
jUbzEzVibUxKdIH3LAJto7RUTGi158m1WRidjYRpnCMDk1WHHjQiK7EmEAFGN+LY5+eQAp9mgk04
FLguA4L3HWfgVw/ShIvdGYUBxX+OP6FiDcHQZKIOYtR/GK7nsMQ0mdAPk6Ujib24HP0aD/j4giou
vTL9p5gH5cSE7uFzDrtL/KqmgVo5hdvrhhK74N3prYNI6fFWOZdNpNXTX+NiDtD1ztwXSXhVwA7P
FRI8k8qs1LbEI/yMiZmynDs/xUTJgJ14u4So4gzBPjL7TjUTKS0Qf0tFp8qHBOoMkx2JiPN61SQS
rMyKpsc/Ox41/SWyOBj8V4o7xj9aDa8WUsIwKjIQPrZW+hCOCoAuQAJwfP9k3H6agRuZDIwP1xrM
d7Cf+KfDUk4C6xCPGGBGPc1Y/N6j+zfjS3FxNsMM/RhA4pXlDceaN6Po/Hmx4PpBR1W8kHrJNsq1
MRtNy+xmgz86tSRHlFZTlYvLgE4wqUzOuGG4IO9n4ymptmrKO9MSGLjCJ2vNc92jvwga67VkHrzH
m8QKK9GNV28fyQ4f3MMI5uGRgLSzk96G1w7+vDrm//+pTyiywn4LaYJFP7yV/I/bcgMMfmbATgii
kWsqXI3R+Zu8xXZBITEq1bp5sGftmFFial9iz0G9tMl7K6HZSx24F0xKCSdHo0ozBUxGiGjs3xIo
P29EnjwQCyNX4wTThOWvcYn8zztxelS0HrOHRsQaC7PrYeQw7yW0XGDhP8ngRVnrERv2WZqT5U3s
A9SRr2xXe5f9pe0Q8+n/QaUp7K2mgGkyYnIUaSlQUTde8/ve3joDRWtSkgvx6g7Kh+oiitnR8UWg
z7E5tAoat1Z/OUE0t9Gpp16lMVKn1yQFb4O7T9rRX84ktzR3z6Zd5KMb9YkpLJMa5+A9F8s0MvdM
MiEblBoM3QEYlfgzdQZvsEmT792X7pzvA2h/PaWr5n94E8qEND+mGYijdNtcIJOAZxTCpWHYvSkD
kp4O4phZ2oyS4Q7zM7+wC03nbUjjXGop7NXhjkfk7yhDOkvK8OqH31SyARjkEuHyX7IRY0BY3ihM
E4I6YwXA2IyVTSJ2HKxiO0gW1j8zr9L5MIDF31t1nnwWaOgcnWIaV5Ydcv4W6iN2F+dovPImV/CY
V93lWzyXiwxfA+2Ng2jI9WMuDQUcfZbjAR2ivO+c4+9cwUiNScBrv+J8aqAmT2hVG4WomPOYDAB7
BpPO8GVmzmcwD78Xki46hr14yTGShKBtrcvG8/aJH/cb1rujP1stZNZ0VwU3OyUqOFh/sEhiZyNN
fyCOEP+51ElUL+2OMM6r9H3sXbrrPASZTANuYJKB0Csub5WhJgdL7UMLAi5Lh+0XBq7JkkSHcyGE
zIehKdWhpejIoUxzdjPCb8Skce5BUrrEKjJKfJht/q10CoEzrJDYcBcnaqdajeaBog7Cf28EWvp0
xTowrXqdb0ENr0Yyf5DkJMirnlP4BgxlCC5bjCjBXwMnvfMo5ABlEEj2SGLuqJizrY/cckNzMzpA
7mA2l7h4e2rXvvVhjXzUl+3HRnpqUq66oLQpvEtEQ1kbb8hDVN44mk0YsJROIE39Sy+Tknv/q7B8
HkC7oQoBzE0TjIB30o6lVnsxZZAmWypn0CixLjnqImlXhufZRA7eHNaKL0geM9Sc+WgonefxyTW+
igKZJJh7OP8gB+5hpvNdggQFJMNqWVY4470UeGYDqtdPj8Pr76xDG/aehsqh4q+sIDOfRTTsQ4OR
i/X8c3Pun2sQH6QdqG65vhsDknN8mtlCR4fzIPLOeohln7hEE6ESHplig58k5/ShGICTFJtzz+u6
OqjaGLvxQLBcLO1MZ0XiXFOz/dE3QCv9OETUKB/2lw0SVaI3Bove8ij3dCBfsUjcXAwKMq1aCAj3
2Ha3cSuHtmqp6iAvwuXzQTBPwNWMFVZ7tL6oa6y44Mg7uYfnaUmdDpzYTbXpsH+9t4Vttz6OIRJ1
9GLvl/JLdh85TA5O3Xn0YpKu0ROGBe31llwtoVJoClbtatnUXuOJsr0OQJwdLdFXcn7FmTXAsGMe
h1vjHG/zaYG7ZIYGdwjs9PisZLF7ov7wkRoQGEmWmh08KZREHdqBAF5Ven14AQW4jwD4/J+gSZF+
PQxcrodNMvcANBZbZrIndrhZvQ7jpHOpWcXjUzXlYtbql5YoWnWqdvagF35Vy8MiUek6TVMEH6tc
jE2mJY7sCo/GRpoLxkaXn3AWRoCLrf5mQE1agOBcnmQQVmRt/efipMZ4bn25DaxIbGS+K2Pf9UFv
6IPWDMuKAbrdEhOU+HGVsq9HIFkr8lzenvV/bkrrvR3u8Z7v6bfznE6wv5bkWXafuxXFF7l7Ky1j
ZTbNMgD82Y4iPXkAfj1yNnp/aglfX90hQpuI0gqi3lUjw5R740LXvd/ekiOYwRWt+4axa42sBL8N
etjifvypREO+NA4gv9PlnLFNVg5QTzdkIOKjiQJp8ouy9HAAGH64+YscDLLxwy9P7tZZSUBEBdLC
LTQprwMc+eaF1EWHRkeOKmstO6yCojQraJu3E38OPfd3gkC2CSnDuJt89Si28QtTq0QHsfUDCMtQ
7FhOqi8f5jZeqbuq8OFvLd2sWNEK53AhT8JbJ6lGpr4g3cj7aqZLs3hwWm/2EA48YkG7V/0fuNUb
YvliM7hRbtl7soG7OyXv0GxWQjUAONbAhKwN+/G4ihVKrDeCdLEu1VO6Ry8Xlf2zP2ErR7Fu5GJk
layloZ8hKLkibZRq6fsJ70yARBZPHn6Ujlg0KbIyB1yUYnNBXbYI98OmmunGOW20xU1z5LTClf5t
lh39RlbLHpfdEzqSwk3gDNL1Pw1Pfy+/mwGG+z43fGbMMumuulxc67QIL20CEoReQ+eADeeZklGi
ssyQuAK+jExWTO3vQxD5RnMMCWTsOPzLRWx4UArBA6pTY/tMjBNrJwS2QC33dVEEXRb544eGnFbq
YF6/E/MVtywUZqO+jMn9ftyUKSj95Gfm9dE/5zwK9IzgCA5ZxoZ2MVo43VRGLZ6TNuOEd0/t5jQS
/rKz5834BtBsPL8pxJZ/GGCMbvzS2SBE7M4Kq3t3EGrkT64i5WxpSJQxpJThB/VqNCsDsYNUlTlT
rUfMDHWwVLgRAh43r96dtPDrSCa/6pz6rQbFJseemhUXHqnz/nzExKREL+ScvN3AuGadjoDUpt02
ysFRuhV3YUg0mpaJ9oQrlkRrfuDS66e2fgRXdDytryNEh7YC7blqOPnGxhVJJPLW1ToqSXxSPsPe
9Z37jeAury5o24hefKKm8hEkOjbN6zWfBWqdlFdBve7xIayR+1A5PpKpZCoqGZsJwcLHKzC+Iqov
w7nU3vJzHvpTQtqOOPWtp11hE26IyjZJfIdY00naf12t6YhcHlJf1H0HxnmaOpVjbMK5TI8lP8ZL
Y/WV1VKLD/q8OQOlOXWSTQhLNsnx5yF1e+aApG5cyBV8ewhhquob1c1vTMljuYHPjjfpvhNbdd7e
ujwqfqhFCsi2DpUswJN7QENEYNqh+h41hv+2MrDA+rZYjJXAlr2ipQzvu1ppa9XUHfZhsxCcd0+Q
IwtMTSFxH6659Z+qjez8hs+eQ4ZCIBauyMtzfZ3sZ3ZJiRRgb7TD02myrKoxSChSW0R/OwKuNGSc
DahJdRtfqF/FPJ1efRh6I/rBh5znCeqCJZQBlf5YCFvH7NFnbZcU2oRtmSnSKcWqESfZvx/8aDYd
QRjb4bzj9Md78aO0ImLIDeHeCl6aL+SOcCjyNBf44y0tzyyohrNY5DICHmwuXEa/LBdW9H6uK7Ti
dcTHee+skBWwh3OMiFXJqhhg6Crj8s9fD2gfCKe2fIaDrQf0NFuaSRKFJnxcrXzN5vwNbZjJQ1Mb
VbQuKafKEwh36FN4xpH5vPp0dv1x+MrMmNWVsNQXDzj9zyXp1evKLRRxmrqlTPqOh+KYuJ45w+19
Z6urrc8y0cXYtO/02jKZr0E1peKUKtcmVwSV5YWzMw4TDnveOrc7ylCni9mbdbfg1ArYJoRg1WxE
6fqtGdm2VNvaZiCfvIPAVvAinpuIAEC2BC86AVCiTRCpLRWociJe3PVWWSEnZZfgvdMeNoJ5earj
UfWuFLUKyPZc5VSqDd+r0yPQsyzhzIKdjH5bAAnv+ao890QUBGKb0MgCI/oKBVz6BYYbPI5oPT0S
qjwYcC/7dGp+RaD1Wc35fR3OQd7rrSMD3XCkgXwi0L9gapLT5ShKzCKneGDCcNklhdcOHIcDNMG7
QAT3i82154Dp3foGv4dcpOHMIzFdAQjN1XXQeVsZNkMS3GFeYU0zcJJv8DO6o5m5QdFSFGbbEgsZ
at9HyKMHHFCQsU9fkssBQBW6OzbXSx9M1lI8ycle2dta1CcHsK95d43g6e8lE9oIGXJGv+Y91EtV
StculIhj1eiIGNJJyqggm2B+KXNhn2OPetKnnbGJA1sPkAeEJONAzuJDdPbAWpcKldwF2S0i0YMW
17dVdmQXgjltadhP9HhEKbTYl9xl9Q5H8GuBpvzL+l4G1Y5SDLwHmS/rUgxq2KOo7WkmlVguprAI
3UJKeqx93n3QAPbQozPUSnqg/ZK1woBs0MZ1fW87nUjWdNEUIKhJmZ+PxmZvApob5dvuOCagAXgs
K6vO/KVgvOEcErmkfQfIEfpSRiGUEtHPOVttV1lMpK7AUSJC7+VT1XLi93coZn3VNG6Z+w54EEQw
0fLXKb8hlTlkfGP8HdmGdPExYuIWrAAzpbnzgtTKEaKuZ+IEe5dOWZX6ZdAEx+AehbLSjAm71hm+
DzFpqMjTeFk01YGJ2kMgKxMIOSJwGmjt1yN1KAjCJJ7s8V9lz6z/Wxsan6xat2j+X8znkLLfhRTD
PWwgeZ7X5wdEOfxM7kLgXUUmDhE3/wT8jHzgVP9D64MdhC6OPAUREvDbUxAbhqLmJfyZvaAJDHNI
nyFsh7iW2lyOCJVtfEfWO4m6t3geHBHHUjAy2dLcuiGk3TepnqQIkzxuCZirJaM4QSncd7HUfBB1
ghE399Va7deNnedWFiQf50YBfdOCxhFHlQ03cLT1s50Rzo3UHPJt6nK63yrjPKMruotKkkuVo/HM
KujL8oy3jjPN3uoE6YC+f9V/KK3b0+RIjABJnQE7E4cBVyAgalhHlZwxWpbnhat+SoGlbFxKJGnC
IUdbe6iaKGObJBBYFu+N8iKMcigtYdkBd4cwZosiBKVoVl9laRWcePepx303TnXuXIfrgsOymbDP
ojMXFj3Mu5KTLcbtjS8+Fd/yy/gywzzWrRvHMTvDTAoD5E/weBZaXE0TycedMQC3Dk0J2/OBojjr
2VwT/TzEJeImPA+Z7MyPC7L5UaOYSlnFJD9nlFoblem0f8dfYp3qkFxFonKOLKqXzl8K+S4v+Ei8
efH/JMm0yH/iCQhl/g+Kvygd+AFfWfstKWozwTnXbrmtwsrfURwKV1Yeum3Ft3tJW6tlpLo1Kqc/
aBLR0u8mdeQ76Yw7wQCCXwA8Mopk0BXGo/ZIzQBbaHCPXIL3RR+zKLWy/3jw7Mly/y7f89EXNYny
AoBBiE4D2Zs+lbPPeHgppzglVoeoi1hVWqqOxurvRZz0pJnYbeMErARWtqp62ODStELfi7X7w63s
zrvg/GumsR1XufRutq1dX3QLkbII0dTOvhSbD2+mGx5whSQ71wZ3vjrRFSr55LN4EGrSJflI6YEV
8iuyJAPr1U/KHNZqfYD+OGH635ppLsKlXFiGcK4sEaFCh+qZGR2eUMs3mBvi8Rv59sWaiCJpl79r
qdFFSuSHA/En9HjHTdl295yIIDwA4I53r9PKrA0m7nnx/ChFORdAFrPiW18bL+YGdW+9cAuSXW1V
d/kWMQDqZ9KgGknHEO+wQUbjKSGeGeQdL+lU1/zfzjM19mN+34dk/ZyB49DIzQEudyyQXD1Pa0FJ
necbrFoyERQMMBGWtVcWAxrGRoCmS+PizKVMyv+kmm+DdTr5HaT/UFpBIQB/lmFPB2SnaCDWY5v6
qJShRBUGpk+R2LwTC4XYzqjgn0LntGSqj3QJeW136UI6q13cb1eG3MBxjBnlDv/RwGaIUZsNesCZ
2xd3ikCYOpCeWqslcIsX9oSBZ6P9AAAV/5dS67YreQxUzz7kkrfFsfyk856DhVus8pW3AAFeA0zs
e6p+BwniQQSapxCvxUHgQhjhopmwCQnW78qYvtAQSmnpv3hKfbGW9hKpFHAca2nP9j13qVyEOLL2
Pz6dQXVnBYHtY73kLbdt5oNme9H9SprGnV5l0K6PVi77mHtGi2/hxY+Rw0xLExvPmKbt6X9nkEwN
gBBlvTZalHCsNIs8UA8GkFAic7i8VxQOX6lm6BMuqTEI93UZJoClWinZcPnmaF22F7e1J2PvOMum
vQEB9vokCpHeYDCt1WPPHyz0ebvnjPVsmRR/++AKEAHsBKVTDSQL/j7TFE8ZZSrKe7xQjEdB/Hw6
mnYN8d6EboBaYbLbhmb+Ymjh8LEd1xVxDQLebPeRFY/95rIT10tG9W6sfEaYLQHNnP7J9bYBw945
SV8726Rj/TJvP4AhcwAOn4A1ql7WxJ9xXz9rUW/yu9tFkgJ8tVqGpiVlc1HB+LjJdkX59uth9Zzg
CzAodxdwPZw03RfenSrWsaetx3MT3d+NSf3phk1wKeTltEBqcvt6CvmH9Rk6hraAQvBPpioIexXW
BiNHZi+z6Z7AsbmsjalxDTmUheroklMJ/jeg7QlQQBuWCsyxVizzs7fAoAZWYAVXaBZ2FRyYvz37
v0t040AIANnIu/Mnk0dSEm0hNbqlJISvA4TLaByPTylLUtfQ6pthZjSd/la4uZbiwy25wU261i+m
3LV/RQDZlUUcjCLcMcgxQ3pg6WRVp3EGUB/OHYS0BwGOUSQQi8o8zLGCy4YQ6lrQnMqMONUV7VCH
JNg0SwkrYjyi9PmVevVwwm9YbMHTgt9IKQeypjuhaqJGy8wBQUDODnA6QexQ4Xn+DewJUNUEypYd
7EZCImG+GQpthYhJYmnHx8juseTC8Wavbz58TN8lxT8S7ko49hcnzxgTmzuYDBobYp2B1OCZ65Ss
LbPhCZpDMJAgRlFh8An3gwTkcRe+3eRxwTnt6TTCYMLuxdQnqJE66s7Jm9S00qu8hac9tUds4tJi
cKgXVTr1rABVgD07d3lv2CGjDnzbeYmUye6R5HkWhe4c8t47L9lmxflLMRghGWzAVzgHEc0mJQ0K
/b9kVNn8wGHOjptmOvs4bOEbcUtDsIdTXcjCszyVSdRRYxAljVjrl+lmhJZE4Onvi8z+DwetX+k4
rdqQjKmhawVy/mYZ2iMXNbUkEwAvsjh0RYuqR0iM1Bd404hEjvThx6STwC9XYJXERrNNf8JOBaMK
S1A+B5U3tvzpR1TcKCyLDW2HfF8fT+8drla5ezCRShjgJSP/qMmTeraQL2awl999jegZ408ZovUM
kRcoAsOOysZrZiZ8FZJoN1OrDQUCieQcs2wuOH5aOjBnAdPRb8sZOshV4obeMTCP7Gpl7nHJjwan
cRzZlQ46Hpj9W13zUF3qMO7lKiMPoBgjxPBmgnhsLEfsI+CZNFUMvi8NzZmKnLtBjgpwjPexfhCp
gdHMq39F/iRVllP6k8z2l2o7OCwXbQxwiWizatADx95K8UUjutvB1gFONTW7jFuVR/RpB1Iext+4
TRfausR+d/017UTfJBhxxKzUAalVIWHyI2QSM8RC9+1WqC97VZAyVet2pw9O0sb9VtpVgVcE1T29
qQntR8XqeUxF3RRPImR+mLF0xY6epO/4Juba90QUkOORJPYrMoOl9ijyvsDI+NiRtI7lVDE/Npwr
UTlvCNAx3H1nf19L2RnDf2hp4hVor/wCmqG9ok+SaiBK95NW1WyxAAyqDrpsc647E9oADtfWqw/r
dLjYIHjJMiwaSDiSrQcGjLhI7LiSgEne1kxQFxMUpbLSPviwjF+dNWrbxN56qLgeLogOhxoaOFyG
jlqbilVnUThMqOh91TOj8nSm68aq2UI/Gka5PFP2CiTH+kYqlTaHs8vvLXeiuiYFVMLkIREgQ4Vm
cAifiAZoO7A70Y1pAZWqTF60Y2GaoREX2QLe4/Ng6vMP1C5fWBamhooiQq42Z1vAhX1U2StmO7xp
uaK6V2gldY6kXwVkbPwTAXw05zFyJEdMKswAEwxQbp8bwIdub8F9yz/taZP+tqJ46rPe2yMb6v3e
VkC/hXqjfNfSIEIDHqwtSgnwkeQSu2zBu6in168SD9RvHZGxJsN4N739o6m7vo4/QfQSQrcXMlec
piQeN5OEV4EGEsjm8wKqYQaNyNJBqY3FjoFQfxVfgFxGcfByrhcyZT83Ed2c4zyQiujoPTcOx8T9
cQczfJAMCMw9VFz05KCUY/9He4ZKdLfW71xSMQspXvZJVZ6AESat5FtsEbXVpJsVZZvEm0MUokM9
LDRuSJy4shb4maNp3aSFpYvLW1X81dhWxAUNJwpzsFMJybSEUFHOH8dV91q5XOUHaimUPK12R31S
2Vvo2XbRkP56188IgxVmYgCq1h6NqQD3gaFZrG7XC9w1A9bfPZIidkPYToI6Ci9nmHGVH4QGPKjq
t59oIWxGXIjipmOuldOeAUChu0nNm71/WP2ZXOGljO4dHzLkOXBExmJ4PQYvEE56kM6BGaAzEj8F
p5U5iqUmuAHnBsVqHL16/L8UHjmVsXswuRP06+aIhI5xVqAPndCtMZTjEDyr7uJNbw5uiFJe2hYS
/Eh4++55tKxDCvT2CxUJ3qpCdfuwIjAtdFntJE+AHoOKK66Ew8VH+NoNBjcUY7U302wE8iV8UCOE
RTamIa+hTEza/Ea2M2qY6tMMfz+Cxjio81z14+krmMDIsfzQW+ALy+j0xINIZgPPHjpRKI3yoEl5
eX8Z79dF9cjYjK4tVjK6HQqVIUTYmbG3kUtdj2pWhPHAYa+8c9UcFbNqxtTu8GUam+Ly3hk3gTIj
0900FJVmw7d/yxGBO0kt+9cjXapHcXoHZl1KJXghHy5Ks2IJCvw+kOgIhcf8WxQYw13Qps3EnM1J
J6dYG4Azro4rj4zCcjzpEHGeuEAKjDVhhaWwjjtrdlF3khYNuzyreMvrCKlDTCMhfZD0WaVsJpfW
1K1ZTW8nmAe6BQM1UuYY1oyc+Wr8ROsB1R2YUBox62Fxhv2/ZdmbHM/SHG2wsMW3dOtATcWI7cJh
nOiR1lw6QbeND6Y1o0Pnbgbrj7ZKtQgklUgC0mTewYaVTcukeOXLAalp7EK7TbY/heCBibSlNvOw
qz4DBt445kQQo64fDGRfEH46MhToYvGk3FM9hGTDKO2nT+33l92W7X1SU9l7bFvj1F41igjmH+1D
C5cRXy/hGnK6YftcvW28MFVBlSonndHkJfN18qpnolAivBzpbUAlfpCbOE8lTNUTMZOIvBoSxJ8X
cpvgwYY7GhZEojx6p0T/IupasBQTObnlexuuquRkm8iLgF6+4TbaUzfikdlh+llpYwNQ0+7iYmw9
sPxAe/9tKwp8FtBcuO6r8Xw2ODUpcmcsbp1CujwnJYcrl9mRxNc8Ym7zgTp1d1Y4v5xz9fK3G85S
TQuL5+27ghIQ3ZMgcKSi4nOsdUCBA60JRl1abk2OFMRkeanQKMT9tE3pFVpqcLd22s+ZN8NOzMPw
H3W477ib+IG+TAs+TRc4BPpZWlWO47FWoRHnXHK7DSM0RTgTbZwhRWeQTzRk7ljoa4WKGRYUMz/A
QSjMbJUwSIyb6Nd6iAJ0C1/tYpYt5By/eQTL++FW/yvJMDF5ZwqXUQ6a9EKtfe17ZM0NnH1y59Wn
+bzGLCkJT3fjyu+VChO4JIHjDBuPxSpRoSRaELs5g7DIBCjgT3WAoK4gh5A2iNN4ria0l78HelIb
JXLRRgegYWePiQhdvL25xy6VgjIwWVnUyYp2DXpVkM0cEPBTVCDrZP056T1r8ROJ3ed1WYjjo+oz
BFjMLf9TeiQWejbK+J0dqi3qycUCn31LjQfib92y/iJO7CqKFrEJ4//KOJthEb8xlw6EUiE3HUv9
11PDzi+Yty3V9hjO6p+yg9m1S8mgHsNIbKpIOthSx1oxstsBJjmtQV/QCdRtaBpDJL7Mrqe5IBnR
9DveFauxwbPLzwv6BMaNSVVNBNmjw3g661WZXb7TuuMk+UIGL7VTPcrGdF5PB8US+RRhB8z8F8+A
9G9W+EZdEGqfe2avCNa7utRewUKJ1ZeqGWUV7nWoE7zQAvA/fDTTD+4C+GRazFbC6bfAehvrKPCz
bYfcz5CYpfVlzDTLTm848ssM+7zd+0CWRNtxyN4+Dl79MRyo6n7GX830OfL2TF/2WxO8a4DOCXkr
pTtfhArY+1TYNZNxt1QGYYrkwP4+/oofKF35wORZ6lM+qeal71nm04rQ+2lddArBctomRvNOASHF
Ql57KemXi4ux+zqbqklOAVGjX3zhyjyKcIv119e+3mIJ1lqvMnfoFOAj3brN5uUAQLSk/HZt24HR
L1Lx0qhhh4TLTVsfb6VRYl+Tsei2YFcMCcTRFiW8uo+c8znrrxWOcPXIGqZkGSzKRjnjQoNRjuoj
2YL8/yt71SaRS6RmFXqeW6dNYH451pwPFJ893fEDHztaMh8KutC8xT8pltle6gYw3teSdRGP1ll4
8Fl5rjzPNYyM1TH2/k/SNZ6VuIBpfDTJ3HlAtyqLxYiCgAQ8icGD9g2Yu4OGM2/Z6vqZCoaASlG4
cRkPB71YtjYLo9seb0IjX6TfMfh6vdfSEjV27JQmHnOm2cv3qt6Daoa1EMckSKRUdOCBAS7wmhXM
I6KtW46iffzEWLwojvhAcFzSAev8KxGlZyqmGYebH4ZOWqFjNLmPydGctqRs2wdQe5647Ps6hh1Z
xPySdt5EVzFI3ALLkncq045Ow5XB4mdKPDtiAzaO6IiXq05uWpyaCSS5hCRFwIngYQE2LLJ5U1a+
CfUhTcuQgMWDR/NIjLH++q+Doa3h13fzFzxZMSJgcr34nW/bEK3Q2BMOCR4GZvNqkLXWc3b6zXI+
uf2ntwRJe/cM3qCrcJ84eksxIJOsCmAqxaqgHx4L02y/ooD9ydmUYFO4Lio3h2weRbmJJwQ5mH4M
Sockdiv81MSF+8FlG9BuA0KaEXp6L2e+TRQhOYi/kLLXOld5Q86AfwRoedchbJ/H1l//QgScufVC
YPIW08CtfayskDKM24U4M977Ygbd2Mzuaic6j5n/JAEYoWehsAbqhkbFXH8LmHF9rNsE4DlTEpan
CldtxcNQP5pk2/HUCoBYMOQyRH6oytWkIJ9nPysjuht/XtOwc7jfEAryZRJPsXnJ3Ju4B6R3+IiM
80Y1Frqwc+w/PD8RceyISrNwbBPZf+GJNrv78lk7syAZLgJ7dLNURElrb0KaJIwFng4DXIZOAM46
kibr5VI+vKJWRBaDmTS3rfgtk/Y2WR5mo5bORQQSq5W45nycqhgMknBStSlfc7WN/ss4dNg/a4oY
jdAh9AUfI7c4BUBIt1HtEXUqp9Fv2QorK2C7FaxwM3pf6vp2aYVGsCpL6Jj7M5ztTw/AVoMMBXYV
3WaexGGevGdrYVFrcKPwYgKTRrr2kBT6JXj1CrZatqo0KTJqDbDUncjbwexXCi/wqD67j4+ERKFP
Cyr9EGA1T0q1JqoxeSrKtX9AU24u+7nXz/k/qKM3DuWAixKVB0JYLXDYsxMPHM31SdZnz52MAhFZ
6d2188HkYjgIjIQx1a8VhARY1BTpMQCbyeJJoZmVanC6ie4u2ueB6bziG3VDVTHiK8N8g2iz2rkP
RajOKihALMblNIMpcdFTzCHInRrZ3pQan9n+16aEJ5DdKBpXzYhmFW+UWRVtGqtJ/YWzCvFLM8WO
bIYvaRrbeNbC+78a+JvF8kp/hoKTwcIGJZvwKkm0+vXbosuKW0HkHpfOixbG93gpeL2zP+ANhqf1
5YkRYv5YM7I3XSEwc6iyWTlFvJUtUKDi9CsdyXQxqlqhbn1k/EJS9oXdcpQdRhUK1ECyjgDSw6Zy
nl5MrwSYdRxrEAUVbdhOiTrbCPmMJEGidAF8NCMibYUsHAxBfeTnkljn19sw2AVvzbB5X0UdQngS
lAe+gh7VNX0eKuW5mGPGbHD4N/lxoLaSQ+boeCnkqmU1pW3YbJqyEzTOVXvLtFnrzFceXjPZ5o/Z
6/An+53Rx4phf7u0tpeLqfJhnFYlGpYCqEOo8LhuZOIuOygPGTDeqmbcjNI/jzscxpoPK1qbTT51
VTPZE3ZvYrUSe1smO8S85dQ9Q3iY8yZg1sHeG1vi6oZWYq9TPbaRSiSYVKitsFqUfS/i+0NOIMaC
AxKrVWBpjWQm2GFHUzluvfzllnVbql++mmSr/G8l/utSOXMh+drcVg7mdLVOBXA57D9NiRu6sVTs
ulAddWB7nXO1tCXkMZgDHX68TDCgeIXetcyIwJFhrbzTkJ+n9Eu8l5mpy1R8Bkzau/l0lL1Pg82c
0tenJYvQ2LPjVRR1M5yLqjq4bYWUuBwMnZN6gJYuhNR1XH4NUXCg8g8wzZJmE9WqnINm89aIAXCW
gZzUJV+AUTMuofTnuP8QMJQQuO1HXTwi1Qg1O+0I3KSyGx6vIXL1e+YKwXmpoObnln+mePgaCJ7o
xw0Dtw7qGqxKibVkzvxsa0XR/gAmwt33uqph2UOxOmgpxKs/ks1Fl9Z4KpHS5Un+p0E1oTOaHVn4
2MtUwNjNcQQRAVGbhQ63DrXJgOPDHNraMcZTlVzUmtKuysVhp/ajZ0RYV53Y5GTCSlqC3xiv/NOe
fOY4ypRudHlWyU/Hk9ac0/nadArlbEPKs8qdWDkygwPfPmvrs484Me1vmNJGowlo0BdSsYBoALyn
Bw3JXg2bi1ao1CNbmGw2BycsQt4Z7XRb9kplaF8xWyd5QzP9zSh9HrmlK2CgRq1kgQlGEVmlVWhv
TLkMZ8483Cn4tDaYZ+LfIZ7/b31DwF8+dCq9l9FUUxnFYVe1MxTdWNmtrFa3Cedzl0n5JEZmd3L3
tG6dskeqMEmd4lz0gzmhIGJwv3axIknU1oP0DL/gCO49VzlGS6PexQN42+p4Wci3kb/AGTbOXt5z
MuvH2ybD3P8LKfeshD2n2Yq+NSj/btqeMkIhaBpXG7t3eRA3joEz+ds4PHrFtuE6Xa6mV+k4QZr0
Ff6fl043Xyj1HpVegkpTIJ1aWa7m6yjz2JbRje11YN6pwNHTbs79zX5OmFHClvx0rnjhi10YcRul
c6VlzJwVQCGgNOOjFyvPkqu7nSAgsgnZCoFz5X6YSWMJdbLc15W8l68dG/Z3s5OudCf4gZhSJ2RD
bLkqh5n+/MYrmKXXmoN5T0EQa5wgpC1RdiVMKNkgj0IY0anuYgCqgri9Uwr50ibRhzRypLS9cfSF
F477LSbIVfp043wSme5CNDOwrkUVFOnZhMvUtaKadnZ7j5JJB0fgkhsp7fq0omFSA7TbHoMRcz2j
AvzXnNNUB/HPxhYWrEK7aAD8Ls/RXooLIzaU9yHY+deiYZwD2o3I2MLi7W1qXmD9PZz6oZo0/jAy
4UwwWnjaNyybtT4T3mrlZKWSNpV3lU07bWiIkaXFEUw1cWT6HkyaN6LSLQ+SbrfP/JE+JLYiPXBo
7tKi912C3lV6E9Ie/hQyfLLaVmqMyfnrrR/mZcZQeBFCsb2dIlTRBDZ3W/lMJPR5XJYgTp6hKW0o
xmk5JDdbyNUh7SpOX2u2vFy29ZeJfCC5Fh4tTKCm6HXcAzQXehREYURZZtQY/Z362oxqNe8MKesT
edgrJ4eGPTB4AsTspXIwBy8dS+oYaUTqS4Z63ubYvY/bM50bZYcqjnMO/Uxr7s9UFUWSYE/i2ayC
7q112p3W4NjDfGKHy/e4jCruBJTAmwA/De/pIjaIbjt7Y5ObckgMheBZKMOzPYwdVpYe/BqRCAqs
uHqABXvxqaS0zmJYxhds3T2Bq7MpFKQHaR+p46Gqy4YmFQcoe0noWuAZR/tVUejhkVZ0QU6qoQz6
YDNxGOOHMpXL8tI6cCll8Iy7G3ytS7d0qf2SXw+7o6lPCL9N+3KnMlzXDfnutcHXtXFRSOYPq+kf
LHXes8omzZjWQj6jnbxr1TpaSqZeuAVrE61eLJzmmPYp2WHC8RXPIiyJ1PxzOG3gvH+tP6ihfTDo
/E7LZfMqEpjguf/fsBn/f8UKvGwpbe6MeUlZa6WV8ZidxJTI1N3sI7rMq2G25H3fE4GrmKAx05dB
wUCdlDRf6SyJVh6Ftf1eoZdq2sxlAm+ipUAM1/e/4M4s2Dv+u2IBElPJ1o+gni14kXUTBQnRkqsD
sJRmAAfl3ZH4EvmbySTbA6GtLGlC62cNfsRgavNv0EMTUQrTnsxkqGo8izXwQ1Uxpcri7aEzCCUD
yoXTqv9qZysxr96KAY/faAn/B59rPZymrCwr92TgxlNVnXJsxITza3Y11shaYvuHFiuR31YdsW/i
Ic1y88FLzOyFXhZwiw7kMmT7CIxDpqlK7xPU667WWbLLMVh0VquWEp6IxF2SnbC53sucJ8g0h/va
YUo6BIk0x2MGjoTz80te1XGlUEpcYMxcgJfsOCFOJbnznRIlWgxikCDfXufDEDwfqzKzYG+6yYAX
5N+jf4nu7aPrK0/8GdycipSEDf2G0miRMfjWMdDjdhfAHY4kKoYNudkobCQ3QoCKwvVqlSQ6191m
ZEBz6fNl8RroW/T07RGQ0EaGUNF0k2bX3lKwpRzLOiV1IDPeY/s8cT8gsDwx0BHEi+gDwRiRScX3
PKHER7JCsCrgPSf/RlR9JIMxUmTPObsHmgCNelmh05JmEXLhvYhK4Q8fptPCtFrRNLPmeTR753fk
rfLkz8DX8PL7GisUagIQreuyXaS/XnYq0Dmh1Ivqn0lI7PJc0c2FKnWPcZaUsD1LbH92/iCYk/Q/
P7oh6JYP96mPd9jAXIr2trWJ5GbAS7tNQgpY7g4E0LSQ6F7cLagDs3kz5MYkDYX59txFOM/ASjCx
plMCKVEzU3lyOD8sIbyOWmIzTeyuzJQUFgSmVwQxLZV/jjlFjHN8Psldbdhj/vRFhsO3wM2yTcEk
Zcu+0Xxjj1QgtDjxzlGrfe0UUqoYDBJube2Pth0RjpmAbEEHdjvaz5mbQrZeMZMth+RRIP622jcb
nyDuigx2WpZOFu0yvLACmT3vDKxqn86HED8+Oka2Ems53Q44iFBKjTl96I/ZacIFjtZ/sjpUzEw1
6kgaM2C0Env+nHty411ATD0+uL5cXNVcLtfkTwD3QJjDOs0JV1eo/rxhOSw5Ef+tGTAM+Tb/bllu
wZ/mO1qTIW8hiMRPMNUUhm7uac9LqFeioK/iWQ9RPsceGRrsbQNQx8HYeU9ld27rm56c9wQu9zQd
uCVg6RINub5uQLmSmtWWzGvHQa6VClgFMybx/lK7Ez0iqsFik6hJ8n2O9bLxFe87IfNXVYyrD/Zu
OotYkfDnHiDOQMmqbhCAk0U/c9uofVoHOYaNf1qca4Rdq8UcarsGNfjwbiIWdvtZ/XwUdV1T6qIm
5DotwjA6khvhu46XRaZ75QnhbCZWFaBnp8kHtorQFtwiZiwPHcWKRMSRz+30t808HeH8WTY1J0au
y6CkqkidCey18zuQnTABVgrhKyqJvolENjktZzrN8NBYDdRYMz9sOrL+zQJD5byxvEFj8igCKh1T
pyUG5pIaKnc0ZnJXSRoue246sVTDZKMET1M71rXV0l0YEkg1NNznamTa5VWVusy9old4FsQTW6su
oJrPBU18thrKlN0mWg9MettC8sPuEot+pO3HZ9Vd1krrPy2i4fiX4U4y1jen4ylodBuyJZ6lOmaN
7UztMjXzXA/tbmCkV/ja3UctfhmUz64ZGJYb+f85TEpAZ9w/Cep9CIjUgURtSeFGxeTn78Puq89E
T17rR+LSHWIkbD3BLs7+DOFumzvkirUyeouD1ht97bTjh+rONewEZcVXVLDTQOt65P/guwwONe7n
foh40FH0po1ArTzqk0ixaNDH3gSccp0L7VPGnEbpMoWCK3NhoEVDPeKe3WOb10gTcKkKPY1SyzeL
fs5BX011qmVecDlxjGw6UXDko4vjlq0km6l/R+PXXJFRV7ZFBk9JN/TiJ5eV/KqbAyYaVWftyfE4
4YJkmydQ5+jjY+rjCfDwIE3TXNDPL7UWbOqqS9nhLNdUgBmliejglLK6i7RkthIARBhfaLDB0+CF
V5arFyttL45X/EiEKIY0aYYzhE9Ilv0B7ZoLNjm1c9+e65HJsFbU5M23mGFPCPLZ5AUFxJ9DgNKJ
TSAl00l5ZdsgQBU2YaOM/3BRe5AonDHTeRY4QFaQ6lPmpOOoR2A5uKqPo1xXUTT8et3VHVmn3gvZ
GInrUKvyYOVRPIRsHjAFuIzUyfimWnXL0x+0+zu2cc1OfIp5Vko+kTCsZ6Za7XrWg+xMs753gMig
0bZ0gWEvvFqx8GES2ya+QYe3PWTUskF4j6tvQie6rBV4wqQKg/HMS+iLJ95yPtrEyGZ/LeuFSVx2
81im6nY89+lg5zl8pUIBl/0BnzlfChuPfloI+yLAEZZFSmP9s3xnBynWgqqC4yOjwyXxkWv0Zn1+
IvQvgzaRFtJLdLiPtynzOcRmrkDGznLlWNqwR6kJdK6x0Te5yeRi8ddP/1luLvrtTKyQdHjkNGf8
NAGeao588CA0z8H/p3Nrzh6iGnQDJUaosUjbTTxHsloVoxVQaLo2eaGo9C2TTnrE6rjwA8CdMABf
y5sWCQwh8Ji/X5R1qaURTXbQ0FqxMZc7wk9upf18njG0jH4MOaHvBYo17ZrXiWeoIzWsn0pTZKSv
OuFa67tuJPUrEhCSqINPfIYgVklrOdKZffghj/XVGdHB81hYb20O3Yw/CSuk5TDUWfYImk0FJYKs
+oQ3achFfM9ImNBsW10CDitW77HmBZfMuFFyon+CxebDQsDopcrAabs9rk8rmeVf85+dWIW3NKvu
Cfh/VpbH6w6fbK+KFstz/U4QC4wjndH5et9zFmy+0dwMcrfTdzdnuQB99QjiL6YhFxpCsKvBLPWr
4qN8wXSUdP8cI2ogtiJfWYursnDEyevxDT9fw00CV8hui2/REoXc5vAJNxZawozF4Z0u0sFARY2R
hQAhEZLwQrnck7gRv6aCGXjrjOu4N2sM49fROOo/utB1n+dPeM20aBzHaXZvpjtYN/Rxy9dXYsSp
FVkPY7AWu7DOhWkG1j3wuaeSiVs0Bdll6z/78GI6jHrk6xfH0UWfx6l1CZniBlqNgQhP4mCqCjMv
eruqRz+DfOfc8AvOyt+spdCctgJzb0eCngCWxST/gJNYGXoUW9oz97L+BSx4Q4bUBcjduXKM1PyJ
tGoqv5rGGZaX65QF/Ud6IhTCPoEqFqkfK3yyjC87oR0kMrSa9HczuX2bpAZd245Lt0aX1yjzFUkW
N88BhVH/RU4Z+fQ+872ENXxzO5U4fYIRVR+4KPoJuvodWJWUm/PrdYfMTEobkqlOWm91VtF1na2l
9niL1F/GQs7u74XM9AKMNkLt6BMDIsXabnkxOrLw2UhhfjXefgpaS3MlX9khHmWlq65EraN4l4hH
WuGkhrDzh7OWuxwT0ONu1wDRmgsiUEjHFUL4wxYyR4rLtCyBFBu6V1Me3jYCENYctkFnopctN+Jf
Pl2BNG7+VtoaXT747v1/xSpK6kLOcrKhgH4iMLu2BBSrpKwNEcpIQe30j1DbexQk0141nla+qul3
TyjnOhjD7SkoH8FWjNX/187PrJl+EYoLMqoDim3OQKxJ88xjHdvZwR9I+y5L/zn7xV6DpZHGNmVP
Tn4MEAhopZv58Y2Yp2ypjrqU/kh24osgfPNKazvqffgzGNl0FBSQoTcochfcGOMDslzx2tfb/OD7
UKURfe/VtT097UTjvHonXh6RtOfyzSlkvhQbKgW8Za9gyU2hgyc1oT+X1o3vtTUyv0YxBCGDyPTB
DKywLwYHpn2CdwhtKbHZ8sDJG9m4gGkXEbvzg+zjE/xHOWiyY5zNsQ3q4cfksoVtSJ7Qqi/Qnqqm
B499/z3XI3O8y4ZNorIjtudj8R5FTMA5EFzwzL+zsdC5OZCfaQ1LJJWPU9DOx1YrypAnnBGrdnG3
9Pc7BVtXqCmfjoZa6flDWRJsk45EQqassCksgUNCd8mJEc0O9XPvx06xFc80zZGvBGO0VEpPaD+F
hYq5UCWko7UDYuQ80L68UOORuUIFMsl00Pi6ipDAqr+LrMFqGFmLX/h8XiDt0WsXU9d2mBhxotig
aWaEGnfw1K8JQLdjqqN3Uf5DTNtDm5ny1Cc1aelkK3wHMMto48IC0pqJGWuffk7vdhTu1c2cxF+x
pxQW2OwlxxaZKKXJJMiFo+BZSY3sKin1I2u7xUcWi29Q+bpSqBOCLFEDe36z7CX5dyU/f8BmUHtK
jXe9foxwchIkG734d/q61CQ6jAsbXDFdENgCiJ7/+MdNBskH8Bvdqb8HBiz8Ulxo8uMsQLKBXBbL
7rPKCIgT1FC+RcsV63Qpe5SCZA8EhLuvPNhl5T1onykrpf+uFwR4n99jVev2Ovv++zuTE8Z0FGvO
H5famBb8yhgR0cj+WGZ0uxdGB/1auGEz0OboOhjxpfPWQluCP12d6taL1Dvndls7fIyfglhd1fDs
FpFP5tpCmt38PrAmthRST1XUgeuCcL5nqddaNI8UfgrNJlVWrCTeHNxvfSV4+77tTFW4J25YzpiW
MimSxpQ8oRMe0rBxL1Nix1lrnRZ7bVS/Y4NnDKq/Q0AshzSX1457kiFCWtKum4lnD0IVGT4cRRxq
4TZ4+fnwhBXv0/Xnmtw4Dkyo1iaaNnqOJJteGZbPONClnnavE/oO7rcfwkxuKUl8x9d8TyugJOV+
xCxcyLB5RgsNd/JqopCM17GhhruTlD4JC5G/xCkMVK3D7emOFxy08/eHuLWj3s+zJKAO4bmyTx9F
GpTq+zP0zp/D31+eg1yooAfNMizaQLu1atv0RjlesMr2BrCK+b/9Bhk4Da7EURMd9qKxrSfE48rL
yrzqF6UQfspEU2dyCbDIx18huSF+Y33Fm2O2Y375uHT6iquKud6kBpIRl+GkIVzzIKQEnimMeNkt
gqn07wIv7ExoaHS8OAHGxf6RFMHPZ7yTE3rK8tspKerj9dkJl8iuB8J3uCfJiwIKEdgoCZhfRCHm
o+qDA6b6Yz2o6bQv7RO9VXTVmHTr0MdoUW0LWk5hLPhK3J0uMYMxWG2F3MSbCf9lJUFNqbx3zXSL
AG4b0FvzWOShANRcL40i18EOUVYioFhJBP1IX02gu48N6a06XWitITpn8H7cbhLjQ8DJt5SjPcbc
Us42xfx6fAuHJkR50Q7lk4NQcZ3ynWRqzQXMuLqf9A439vG16OqWZfZS7AKYA3oNrC32Pa5sY8Fi
vNHI8LhOEfWfyVAk8RQSy98r4Qtjx3ZNZutkhfAwZ19WV2IIz28nUMgoHiYRszjg1W7bC5ZqKUMO
3T8T2Ag1rt2gQhCJE5vIo9rklEdqIJslWuVoQo5RtFEVDDlX7yLZoMVqELtY5+Kv1imeM9KWBPtg
/rgwTuJJdapvVDkNpTsne5EvGCx+NsPQ29OQ+DdimLAwnkwHiIcN69vgahMOX/xUe7RHCQw4XcFd
45F9zR/9zpcbwFoohvGm9JBTisjDsCVcwo+8M6ktauUn1hSroitqTmspi2tXbMlU0CnoOxvjbjHB
1bb2nd+suRfcIjS3K2xOhrqs/8D3xiH/xD95i2byLchP0Zz7QciwJ6hfk2lryKeV9WT5YxKOGaLc
UPOwdq1BMfnj2We6H1yicDB7DAfYUr2Dw6TnlCgkUaylNxBEQrsRTMXSYQZ///G9A70fWrbwd+Ui
6Ep6Dfbfcg3iGukkQGoXZPbmLConpedwyF6N0eaPgoKbMO5yarZEAZpp6RkEAp0bLdZYdlatNOy/
GqODyzRBrngD0Sy68fDk6X2r4SxEH7OfW3hp491VrzM40Kn9RKQHOsvXPN/jI320JsiwLJONrija
HleMPMcXZh5AZW1yyw2dPR2ZBMR0p2eq53cxPwYH//RIUU7McVn9v39lVApJfbROgOVBRPfzFJKm
TRfWcXxL+3x7W99L06b34wkXJKzH4f9Xd0ghyG+Q/FpF0GErTbpo7XRvCS9MZ/jmr8Rv2WH4dCwN
aJtRxO1SFh7sY/Hjt45F/NeSgvWacmRJfhtVUolZCodsxsQC/7k7tsE9EbPCXAbv5Sqg4ESe+gYn
cYxHTHSfNZ403DmQrvXKno0VBHt0Bi9xcH+yoYb/12xiGoWPNMMTE8bL6zkGrMzaz8AF1IYT491T
ax9Q0z+KkKvrvtymoIWtWt3/5XmUp9tfvZQ7DN5a++vd7tTDvaeCLCbhERVa5svLwClFhQ17W1J4
VdW/MQrhc2YqyxP63a/Tz4ExiYrrTqs4cLvKSA04DEyjYsHboIVHe0+SbTYM4n/2LRerOWCJ1U2x
fYx25TiXRSZukbHqpl/7wJsyiqLxLixcMDbmibmH8z+x9bWd1ZlPX/mppUxbBJUlGxlJTT+BvaOd
prDvrwVz88EjXSlIxkhIXIOcTeMZ6w+7x88436rygbquYUTqAnjdXuske5F3ZJkFNrFQDAGyW0Ds
bDnT/adEqpn5jv/Jm87n7JOXT40TQuKIT5jMnHBP+rLRckIe0enY7327YqUbZib4aBAHFj41jFND
yQ+hcY58CC5KoYP2NayLCvn+QlaCxD0Oe85MiGH3/cHz8ofn9gF+g/wIshXPxOH2bDJ233d4ItIW
ZU+KATuZrKwaRcStNDBj/ihH3mXCpIwv/VaFMGWNKaTe9E8ohkjALlNMIV8wlBoVC3n5fCNLL6Pw
q3o8k0UWx9YbVQG1NJI8vkruXnll5xxBaS33euJ6aqwp9/zFOoI0FdrjOgyNg2sGIb/V0xmEWR4/
YI2hdWECeZs2wv6xgodY51EtTF99+rGVonzxbaTRCT62yF554TrYykVYq1NLX15W9kgmuefO0g57
lxEA91/3ASW09ExP4yR5GqDEH8sr/uPV/NB0y5zQK3rBX0jVFwGy0TtcWWGzi5YiYvL/St3mIG+0
Zz7PcKXuh4RnNfIosgZHqEy5NZiEzJPnwtL9PsbdoYRE0qM2pE+ykzv9Q3Vr4TuCnj8dja1SHf1P
dnym8EkOVq/zGA919e5TlVAsQqgPKqm5REGwnbeJD5V9hcXCWtufDZcDt8aDN7BQkU6i0h3hMWzf
7Y8Zpo5arjV3wdmGkD2suS8O5tnRR8ZVvFRpu+Vn/j0XYMX+6awuBIyD2GyFX9Ykbp7MF2Xp6eei
G1l2CHgXdlUxq8/C67tgkH3xkhm+HdPtFgZz95po9EJJzDwK7stlVxAXh0RGn/kEpBn89RTL3UiA
KG02a6eM89KgTGRFJccMTfcbi5jkkCQQj7hQQzKnTzt1YEr8xXwWDnlNZ5JRtGbWQMHsUyQpjOlz
8lKjJ3iKQNhvkfxgkYzJwxZq8f0y8moDHM8DQiCnHKXE+qHmlVxi4cFTjv3+ogDAba+IuUCf1JhN
DazbqNu4BHO4dI+fS/CTGDbCdZcOGvRM5MVmPA3iVqVJPrHf93zbtgLvwHnJv9r/XjRJ4Hl6v4TP
akuMnLpEAD/Yy09prqxqT7jDKsJVSUpwK0dAQgaUDpMM+6q5i+HMg2syFZcuZ3I7S1CB7T+pvFxK
yrcoPKOwQpuPeqOD0SAgX69DUL5aPWdp+4uD3nHw9+zdTZ6gxWUb8Cs+OLoqnPLZfvaQhV7xZtNn
yfOXr/IoTRxdGDpV00pq8KudS/c5FdvFN+/0hgRlMG6Aax6JN3hDS/IFWWPH5Ziwk9QeaSTDVE70
c5muIYPcZylhjUp1OKFonbeHgOldK4EaG5Fa3WLvrVnU7avt5bINU5/KCz7BrNqUjglRinvgeT4N
HXDsq3LJxMGXp6xvA5SG1TTDGSO/SSSKhgSy/ET0MngsgS7G1hsljKwWFGCGQEgpq1cMF3F9Ng9S
vMp/hBQVRLEIa+IHeSX4IMGX9bs6fWgl4Hze4Fo/dOQmXGET9SfPn2IgQh8JdiN9/f+OAs3+1htl
dU3JBfOe3h5MBclsDpc9yZPc7noUJbJ+mZKluEq4+zJjZpMI+MxvB4EzKXApSjNBDhfnd+a24XH5
Rt0c2CC1QhF5+tChfRBC2GiQqwJHY8goS3uRe2TBvsAUNxPzGcX0CagPLL2Q2i5wAERNtEE/6Xwa
D5qf4JOtMSA7aMgbttd3hEV+y3NGeLP4r3gwgkrN8qvwptJFuUH7ik7j/mQcSrnT36NSXWbBTY72
aaGiL12798T28KWLecf4oDC2BftT3IW+NOWiM67PB/QaJTyPzBwGyFLMlM+L82LmsDnT21KAq87a
s1z9kL3Eyoth/Za4NfKu7kNgJw8IkQRt0URajqXUnhRY5HmZVEEbQk1EoYPMfOejYEEm6An5IFbq
/l2YEdqg8G+DbNkfByUxYSZnSCXrsVXcwFyntmiaq9kEMRFPZddWZOOli6LmO9a3DMxplie1+Wsh
r9DSJ0Jzri/Yuz3BvSF73/AN8ln1Y2kYyvvibnVCPBgBn2oR/puiwNKNd585g1fGhcbpjAe7qfFs
eJ8G43asDd7PT2cuCLcvL9LCHqRc8Jas3kkm1dXQLCdvCes1mdnplPCTCLOCwEVQX+cDikfX8W0d
zoXNBwZdpmR+qdlqEuSXPu3C3zCfodBSNf3VMOMwzDICwaX7WtpV+DAX0zVvpJXGR+wxlkApFRus
b69LiZEKEIIwAWDQhSFp/i2cpqLNaDgbJuf8idzHieD24yA+ETrW1GJp92LY+1k76OOnl8QNA3oW
P9LGI3EO9cCjBi2ex+MyGFOxa5hjU/PUH7kKJU+9JM9ny/e4fqbloxfDB0HnswwMV3yZaZwIIPuJ
EGXuSEQjbMYN/UKQ0a9qkaw6qJRV4UDYkf01VHK1PkYH1H8cn9MuibPyd/gw3XARYIF2W1d3erJ9
KmLAfVPxMIGncu8Y7iHZOzDnY4MjQPip7iOpBiF05G+gLulH/HTKCYxzXJVfzn6ZoozbwrXTUJwh
OBejgCQKitTdX9ARyHnqX+KqnrVyEEonhCLhsKTFDXRdrnnCkN7CfLtF53e30YJxb+p9sKweWqkg
BDNNpVq50Vho994K+GDQumLC+9Lj8bqMyaNWLhUPGM1jrglP5weXf87K82Yv+RlOY/qbZ2OXb8uO
rCdPsCXu4IxbHigyM/IEqu0WLze9GuPmLsNpxYl58jGnfvTiHh5qozVv42mbbgheIEXr7c4oSHc0
wvyxvkRwfhIufb/Tglkin/EFyhaQIe9vKZtYhto9aDezjRBw52S21iox7WP8OnClzfvgrdJchXUg
Xtjkwo+V3/RNBI/CWGRA0D9QQO8kXqXYCnTxWfqC8YB+dS8SKt9OXHmhPhtraCSmk5aIihikaT9g
cUck3/5mpL+syg/fVsd2hO/dk32pP3I4vlFcTZuR14tq/2lvZNu78p3g5tQlG2o6IU0d1xX2qF3q
wUSRb/h0SiQ1eJ4Qtw1jqivY9k9tecKkG/6Flbn8yI/NWShkoNrjf6oG6mvoqVblDlRoKpCUWq1+
Hka4JYeQMzdu8ag2/0Vj5ENdEgLtDtK/14omNULlYnSzlSccG8zQ6AqRASRnDtW1tAVqp2W5Es/4
Ib43JZ0PJ2CnbOJ+dgDmt5tm1oUX9XMxrMb9i4QT2if111AINZZ8nBXcj8GgiiSqfEgPo2xu+NTR
AT1GobcUSSrSRvWIUJIXS7fdN6dqvjKOqdujwsrx0r1o2Tzb9FFSbzjyc569or9GfSfCw/OqBhzA
F5bVkjAbDasHlyweGvut501Nuyt2ueP7/UgYwrcCQwqVNfiL7B1H0o8L7v97fM2alQq0w1roSjmE
VV+wLTlo7k1JlaUQUaQWqH92s9G9N8S4xVObBZyXV86mXYEutyGYqYXgkZux0RmurVm3/iL0JrXF
G5LGbscAmIsRiTbzmu9aGtaGdxOFmrTC9RdthAfyIviiDpUjoy+JHFiFXx84XbJ+c98L9aV2gS+V
lmAMV2KiDkbXvR1l2ImuGgqn71PO5tM8Ds6qhXOqwHjfPfSTjjWytfV5hvru1BvjDmC8QsRaDkt9
t2Qxy8yWWOJs0UbZIQi0Oh5gMKBFpD/bL8K0opfAdu72AdI074tVxuNN1bdEoH4+RGvJcZo/5Niv
fOdBaC7VfEZ8UbrlCu5WKnHxwc4xOB/V4XPpS+olD5ZSPOTrm1LJShZ37ALrLPTgpDxCzuLv+q4c
UaUAB5jRwxVtsPjxTmX5dLo9RIC9CKQZFFOQrccQzKfd9vpAWzqfs8Wib7ALl01UqNK5wa2SVerF
+YuWQ5qCkH0bmd3dRoZ9uhWA7RYo/PHmfi4DGdE7gBbLCNnF1IDQOGmQWaTOZl6/xkSFeLr6af5O
p1G1LwX/PR7djJopTB2a9pB4EK1ZfC59wG7zU59n7PrYtL6JtWdAWEuMrjZZIX2meLg7VstrM/wj
Qdpc/42MLn4+3piRwDtBosz0q/rPsCrmyWiKCPybTy6ggFp8ZP4ouoHdpQJXUAu1UMQnGJC0T6zj
m4bgPBzcs/HMrOkmzHVycTG9m8/YvH1P9ti/VarVoZWfaXJPJKkeoUKmstiBp/YodnYRQqQbK4Rd
1ez/eXxHPAc/hot7YYhAy+m0323EqK4MjHnMuGDGp5/1ZDCfcrnU1G6XATDxarMJKSW2oFED84oX
6kPH46bcL8oHQNDDt9X9rTb+4ol9u+TSghHSa+LvF0dJckrmNF2Ac45SzW4s+rFeilDno36BMDbk
rYA9f6i3fLuITJTn3FWD6smZ7ThSAINkMifEHEezNTWauThQCyI6p2DsMlcmhNfjyntfJYubXp8Y
fkkJu9y7RGXcY60M5xVhfFzDLVBV5cNehayCJnznK4/d0EIvOZfutnqZui0x+Bzx9X0RKQvPJYOb
c98q3fWg5dyDTh0kS1fNlKKkHDneaEvIMuZIoLJE/x4NRd6mE6cjTcDXOO7KEY/nIB3p38VBdr5M
WVih+/1/13konSUuBSqlT8ifUVnpZOzIAct7ZgbfxuldHO1YMirZJ88gqd+Fs2HK98ArinQk6CAO
P/7t/LF/VxLtM44MeqjhSMHFsUhhXbjkueDToswA4V8mPlPjXSdDwG/zWXtjr5IcVXhoD3wGbfEP
EU38nIezdUnTpEVz/AdxMFjrOxhGjycPvvBxFM+gYMb9I22CP4cmJ0TApclG6GW7GlLJFxPYLk7x
LxinaiN5/Q8VJPtIisOuQHTilpi3TauZQ5vLXEDDqO5VmbxXUdEt8ToUjsfYw08RsmcEQzLkG44r
HN7OEov4OO4Tzgkjtf3Y4L2jt5rtt90PYm1uaNkeCYEncx1M1CjqAC8/nHKZnkEC+Go1ncE9YyXI
4AOEDaKqAt9pI4oRjcIVZgACuKEANgnHsEk0n5aROpADxKLoai0H8zyfBKshxN0gG4NrHQvQRTd9
nEDcPb8xdPNLPLf9Wc94sXC548g1ApY8pZYVEwS+plmJyxjlYMU1DrEyEkwPG/Rplp8If+4ihJBh
1pZ48kLGvBfmHGey9f7VgbGy3Dz65Pd7DWu4xSBZZnazwa9yYIuV074T0OcUSyjAdOlcQ55Is1xG
t9+Tuj1Buk8SFenjnKxnge90AC+5rFA3mATq8MZTKXg52CwvU5HMBLcdZknxzmKOsp2yUy6pY8GG
gnfUIb/HaKm/5JQa1n8T3PZDHvo/aK7nE+WdqRjjqi88E1cLJumjclU6kHo99wZ0IGiN7E19Arn7
WP4yqhBSntAw2dh+Xv+ALVhtjgG1k2YpSlToVNL5YNAYC3GsQkCw9rZB2dKMa+sTBTNnKj4ivVvm
QnQ6iaEMXZFhDYMCleoLWYs+CxsZj5UGsYUpTxPJpQrAhpo5Glzr3IBrGGuRatL2FdcZ4Q2eBfoZ
HP2EGa4HfZyu/3PVonPpvABc26Hc/M204CEOcnNp4vxfVh7uSyb86Aq2ShlaQKIrqQ+VXkRNWWmb
b5NOB8UvvHSXwz/+DlX5PNESf0TuzOolWjGjkLmQL4z4T8cJf7qUmPLyDq+lH+HPv7DI7KDzhQX5
SaoK09NCSn6bVzJmF6FVqTZj6ePc0OK15JemSpsdQ2NvzygkuqcJ10+zsE7JLQKVSBnjccOBvVaN
biYNOMZ7C8UPyldt1L3kPLHCd1q8n9tLQrxnQ8cc+EjrJD6SqL4HxPsvigth/3muqJSbtPn7R2WX
EhhL5JyqE09f0R9mo+MXxCQN9PBtXDzTrNrCfMUHpwl+F+sunK/TJOfSNSi0zJ3eBfdo0rw/X0u7
lXpMzzxBdgYJrbw6dS7kmkzNj72mQIqW8MQHDs70ALSQbaMjDMpE1GBm81jm/DIhzaFB2QKWjp7O
G3e7yk7biL65M/POcnB5cNjY9EAs5CiUuZVOjKh/tFO246qraAYbQlvyeRPWaHqHB6sNIAPzNjiq
LFxlt7/azySkKQToJ7/AE/XUQgoFtBbKEMuUtU/+ufXw07JnvszQVT366HWdq9xU33Wmfx9YcLwQ
UhejY3XPzvrAFQfwtdEByQ0mzh2A0MHq4uZ/8ukv834PP1V5rCCF+vNzSg9udw7S+rhI6yLIsqlU
BpX072vPv67ARop23xwNQFIgDYUsBVdm636F0fbloYrMMlkx9z0Q9S+YsJORfs/vt2G8Zs+tEWSq
39N2k99GDVGfZeDFlV/dPO9kUqnt1PUA9GzfNchSi3nWqwVRzy7y8OKckIcMYaMQw2vkUkj19Mkx
QagqzsEDZay0Vqdt5+Pt0b8pBUQdcddMlddFFIibtKnMcNGBQtzeyjeyP5p6Jooxn0C2hPPdu/8Y
Yef+1l6uzhUVGILKvGu1gelrj/To1dPHKMnrcYBz72Egr/FIQUzxBj+ubhXEg2lz6fARKDpkRm/m
Budk3sTT8D7vZ7c4rzkCaNBOIySj0vshvlu9rAiR8aQFjrCjAiks8Tr4hq94tLj2bRI9CbcBH8/J
ZXPsL0qB8v38aQ/tl2hyweM3gArtme5R/IyZV0fEJVYW1kq77fafnjzy+lR0G9Mb1FjK43KYGJjS
5ck/UAdjsOAcmtDhvVBXptJZK68wnNt5HrsLZTp+O2rE/WIMzScDjZjXhByGBilZNebb2/FLxdPt
+rJx6hCsAwsCp03BY63wWPfWVIQJrDfILOyA3YuSuK2J/tDAqcUtzQ3nHk3U1PGeIKUY8BULommn
uwkLPYqrpIDfrPApVhE2eS8vVNRAvoI31RdWNlxjkz3SXMwSJjU2t0fwV3AnLpvTkZZp1hXeyeOC
lsE+CmeXQ85NGm2nZ8JLSgVS+d7uaHPlB8IQanLEDxa6hTMZhwWPPQLpZMhkqfnKSeSyb25UYxKm
gAOLWGMgqGp29ZR8mxDfcpCtbWttA06pgGkNKZ6TiRWy+IKHYTRxJFsZbNNhFjRzehsuCPLnJYz9
Hyo68XOMmJRmCuXhOGOK3UeH6L+NXiyaWMJ8Mc/akmQP/OYkuGbM8+yCXwoeIo8xl/ML9JvNkhEu
39VfHsNiDn26oehHYz7Yee3O9QJeiMN1/G9G6dQaG/QmsrPq6D3+En9ROOV85i5IFcsSIyTqJ0tX
l0F2f8r7Q9wZLTBnTNLPNmu3C9VrnN7MUOI5RTSt/BENG7mKEfS1wQ+wEfLX9HAGJgxWryJZnhxd
dN316bClH7vofDTGV7cZrQosyKQtyFjfHCid7A6k7xPJh9Ok1bJj5W7kGEDpLP+3UJptDe5NreI/
iwSXyozgrazRVS6T5batGoT509VTHQgzpve4XA1yp5DqmPf9TDxxBn24FxKDtWGOu4LhEa21OPab
vCEuk54QvV8/dMvzMoVL9W63qOwPz6cD3aOzTxJ6t7064Ioh4CybERBlG9IDZ65Y0CbSrx83BeKF
fFxpvRPZ8gxORvMTiTGKq2dZzsVv8bodQ9ioV0uBOFitIwIUH4Xz8I52wD9+hpNh+yK4Zd619Iv9
O8Lti2ZGdiNu1dhNH+0SOzmjm2peO4Ep4onATS6Z8JZcQZB9iXT2bYW/IvMhhufiZ7SbwCCJETuw
XEw9xuCuDRCsZOEu6dFKWJ9svFsBYi/ET7qFBdSjBu3oqZUsM765D6/Mh/3kJkX5B8dpXK11uZi+
PUGj0+54pO3s/cO/33FUWit9cahHWKd4/lUxvfWgWQ97qKNS2cIZh0FVvDjj+DNi6RhOSXcrSGnu
gS+2py9FWZHofgYRbapN4Gw5hoZLQoolnNlM8sEXlB3gEhbdk9xUv28C9IU5Y5LzarY0jWmmBNjc
Cf5RGhxvwOKqOHzl+bR4qtL9zoYreLB3VSgZ19D2a41wh49qyd6xLG4F+Fft0t1pkdJCcoYopQbp
M4Zf3T5YSkIl5qZlcJVnJLWvH/NrEg3Kyg1WPDy7g5Y+0XHjzhJ5KtP0KeaoHEunwGf/HjTyIWNw
/UKwNo4K3bAxPFXxjm6PoV/ja5eqX7gmLoioR/FN2TK2ZeAUNjoV32Y+/YLX25yaiOUfHaZTshYV
WTAr3pf5YbZ5/+2oofHsoTcojSm/PqmMlanC4Jek+JgeM7oOyA9siUeCD0LB7f6TTDURqrlOHffx
NASQtYvR+VL68pIDlCcZJ2WmvcWmuTcHVMyBI3MzhD43WiPOZQbGBsTGZGT7+eoNVhmglBEUgZf1
xVcKReiP5U1GMzzbl97vwd926CGyG/xDeGYeLxANlMjB0xr1QevkvNVvkhBoddtvUD9QfJNFY2nu
yJBhK8bRpeS9BFzrvusmLjHPWzknXoIlWKQHJy1zeUsHa5F3Zpp+JuopMHGWvWH+2dBDPg6xkV+T
CbMO9uBQytsA8A1j7gcxNu8eg1Z/IMgwtpLEMu8PykxTlHAp3uknSkqCxi8RuDv95NVLgxofDeNn
pkXTCSmxCxfPijN9wCX1ggZxcG977m9HZ7QlgVManmkLptM+cyFscIw+O/d+dEs559DSNWvqJqE4
VpAhLDa6hSnCnPdbj0zkGuZJcqkVPQ5UC0NinLcN5iZwG908MNTZp4egZ4jgEKUZzvgf7WkYPNI3
EG0Jybxxyhs8RLx6gVuwiQD9T+cw5lDsccSu7GwRekwKO+TmWz9sUgFRLjMVmNzzV0qos+8bynlv
ICJ4MW4pccQvjjSxBxRmwWKeDOIdlicKTtBgwl3BzHYBMSz7h9catO8r43Ts7ZNVTImlcCwIcG/X
DkuRPk6SMH1Clsi7eRezxl0ZoVZDUr5Io98su7wwLoBGCfFdN2W4lAJ+QRSBJ12J0XVAaCRk0TsE
ECsj+Tq6n/hXI8kcUHsJN+19myBoAaDj9Wmn+Zl1h1FsPJ9IMPl8IpidxHIJY7NUqw9ypmNtNEGc
XypBOuQqUf3v6o5e0fZzL/fgago8+cncuWvMRaxLciioW4hSJDL3Kt/Lm00LrGP5xEP50RX0yZwe
/f9saU40NGa1vTeH21V/4joWMseJPfNADvPWmSA8ri0C8YC11hC7wu82FGimhzIElBsi4uDKWGG8
xL1DGc3ATrrJtobZ+/fdRAEOrChu0p5oIXK7t/TKErEfeSMU+1f6byLb1npdDv2JQQ+fIKDb71x9
15sXdUMuIhFqpIN5X+JyeX95yc5MB3oBU+VQDd75TiD3mDMI5L2MBSL80ngY4G0x7aR74/6xUPGj
d0AFD8+BeGuu6ebg4YEXhM7k9hLrFE8B6K0aOWIG7h1rskwBeFervSQOAmL9yAOnNmrwWWM7j5MZ
P6mIHgBGE7QdikVtYRA0px7/dj0fhQZYkCLFBrV7CHerHh+3vG/GN4Amb5BHdDSsUqESNZFVN0mL
nITZXr16YYpNPGFEeau0nsLUmbj9GAg9+In2sYgB6Yb2WlrF7TL8iumqy5tcq2m+EKTtdrMSf5vm
jWleOCaWx1oOE/V/Yd3WXt+GeeXmhB4Ci7QTi3IZkSEei6VZ5Yb/G8NsPCI7Re7rWBFN8ZD6noXz
2sPRninBs6G/vOypF89djxbr2Qvke3h6dyULI9bqFlOVCNHhanlsxldCWGaFfYKqZsuz7Bhcuc+v
dHdiICZjbo+kZ2s9M/quQ8uIT4MtgaX3ZV/8NTsGkZoVwO9W7jMRDUKRZAMjgQXtSEM9v24tHU65
MvBnXAFJJZ/K0Vsp9jV1nzIgnncjayu5LABOeNKpNI9KddbTzcjjxGOb52QuragFhKmvLWudPPnK
JsBjCUKuB39wkYDGqQJqMYFMqFr2PogHKqjO3OzjhJNTjae8lyx0aQYskUiSOWHSxVAVTnSqGDbh
MvjPQJvDw7dTEQXlXNoX5OLP9myXe+hhnTE55E9ZhLyb0Ra2SB5oThSzoGLQtLb3MB9ChKXRwCus
6OJEz/r6qvsjFytH4GHIK52THt/gRw9uTrcrAyhC2mdQhaHm1ScEE4WFyEY3O//EAdZEY+cVgT13
aR2g6gYYUmWCoY9A/G1PoLZXydfD3EsCi+oBNtbEPkD8sX628irzD4CVVABMyEfHe23b3NzDQ9nZ
UIQSLBNZm53slBKSxNukNUXfqvW9+IBUPRV8B4/yA0x0Za6W9GYI8zztdC+9DtdrNmbut4ZBXhUj
s0unWCuwN7vL5lfpCnU7vJpklxCswb9cts2fEtL4d/tBlx3ele0TO+kRhUOO33aI+ovFACRvXXq4
bRJd1AYyUab0BcglAZoxiOPfAzgWptZl9Eo+Q6aULWRK5ir7pMRyFibqfh9g4q1ry1qO/L8Y/vzl
7O7zxvJx6oiR66eYdsuWXLeNToxLvBWSayJwdbCLvm3HHDDgGHvFDtd+mcipQ3zFqxfKJijVPFtA
BZNpT8FaMT1iZoyzgYSRzDIvyCioDYQp1Z6rJi2K3/C+2DAVUTRhEnPoH2UtttprqYotcuGGMpXj
VQaPAHZW9lYJqsxcqicdK3uBh0pIYf7AWlGfYWEtAYX0eADkvZchZ2kMwok4+CgQyH/jOQWb7/A3
Au/whSrqNJGry/L5rhYeZECB/NL4/yH9QtTe5M3/iygwKFV721VQBaj/N41AOI13boLN4viHI358
hhGXQ33U/LsscnQNAsARkbbsL0Pw43EsCx5zKZZxeeTPIKQBuJ0LXMh2QgSCwtN+0v+gKboyJTJy
OEDlpSmOYJt6JtYlhWjjspgPJdv+4BYhQppIqhqp+z/CBtHiRKe/E4GjRi3h6PoHErzlSMS7qNBF
aA8LBzNrLbcNgZiGDoNBg1V1h1Wpr0AdcY6NmFj7em98vP2JXSzsyBEMQa5cBx7I94+Ck/gYMUoT
uUV4IIzP1F9BwoRflxVK0N2l7rE3WB3CKVRlxOFwbo1KmvPtIkt2vxYxJCXVWZ+487AAuOV1rmcf
fNv0pssrlpwLH3usbaMR9boSwfRtvjt9L05KeQ26cT7ADL6OUkKnhnVDCnhbBpuq2j3BQ8pp+bFo
bHLN6bh1Jo5PEV/jjGKAkWAB/97KxL/tTZvZucPYXSswK6K7goNTzSa1wjiwoYswebdj9VK1ajJd
s/AjL8/nci+scZgnxTir8wgh/7KU+g461vNK0SuSHYfxOPKgPke6Lu51Sa1K9fWUDkNRrYe9cCTq
+KVAP/W743I+13XK7c9+WNcLELCieH+7R1Cec2/Aq3mmvEAlwvyVTjxMHPiBcuoiH4QeG5FGvC2u
CGRG4+ilaPl9O/zcogyaJhM8EvxiZCpEU3AVKrdqvP9fSXSQAHrUMXk/8LPId6hYEFdZfw0LTxrq
cLYjZ4wu+xNAhCJ/UO0Z+fXUrYnbDYnuIzgb1oaai+hGAA68KpFs7sjvBGvfWaIq2LKBMjn/sUeL
2oGpd41Qxd/uk3dH6s6UQqGwyfg7LEFowQ2i4+LAbuVFOqwx9j7wVuWxyGtImleUUPuga5SvQp2s
dM15PB/1L/jlpphjTUvwynK0nf3jfbY8sJqn78XguAi4TgBhYPVfYYyfD0LX9UTFEr/J9ekKR/pY
yvfYn/f/tbWeGghrOfcgFu7UT3E1Oo/N2lQH0eHBg1elUScN7lnoIF86FAJ9WazkMkDW7HJta896
9CXlqvWQrw/M4OwWQO8Cb2wRWreE7SU1GMdiR49dWCWLhE/jGgVq8/IHeLtdwYHWrZ2QfERNIaQ5
r+KuRDJtx8vfNUK3I4KLvUYxEDbjbpQRaQ1aQ2n2/SRpNSTCE22F4RR+CWPLQlC5I3t4a3pwLy/3
3wmXHoDabQ3En/q2YHghpI1YzReiEzFPdA0epCYsVjQCk16meQ7jV+ZjMA06Sz5rfpkyxLerAL/r
W6FBkj5PSLz8iDArjHFdTA5a4v2F1J8T/g9k8RmpNWKWYGCM/Apmb1QYXi+Ks3OMSL+cH7LqJvfR
0cD6CpBF86y+xzekBw/AdsB53+zJHz0k/00X+hpeyYSJVPrv1IqWQCxWZpuBPP6gWWCdxDZQgqZA
UBSMekXivGV+yw59zblxRa9ahCp8ojKJBNQ8CZvoXnF+9/+kIqPfypLXaTRdvru4CmsBfa3ln/V1
M8kcPeNXsfUNCeGMS67IPxLa2rmbXxcWDSVV/uBw0UbE1IjzJ7ZaS4AlJHCs5PcfLEdV9Rdu2TPb
EF2fL/hp/VGzjDytm5YEbRqGe2sAyO/MbaD6k/QS/wmeeRB+ISGw6XeCh4QFKtkK37bWQXWl7eiW
qHaXwx4TOxftAMu3EdagoHqfkW6YvaagnglaJDbWmfRoangH7S4gnK9PFLxwV1ItqbpVxhamrGfw
ezAvZT15YBUUvpzxn7hLd6Q5r4jYKf+8XZV06gjHEjf/BeIRAUo+rWjt4aUGVnHYxwra0iGnn6hg
dZE1PZusqFyhqvxhusAvxtQ8N428bDLCO46Snx5BcOS5mR7ha2CimQl3tCAsIUIed2CSbnzaXzEz
/7JDbxYK+X/CWo4ugpd6olhiivdlXngkx410G1LazpddKkoqxXTOSdRmQ0/lQIVAXSZj3Nkq/QHu
A2pHygecSZG6MmqK9PPrSHhtj59ow516LOsi9MBV2x+dKVsBQtWFAn0ReAm5ylu1bAloVgJuYP6M
pWSk8uG4GEx4PhXWa6mmOMdEPkpYXPDLghf+1Ee1qw3NeMgwI2iSLVHl5/fNxPHb/WJS9/em95AW
7Qy6FVJaPjT6HP9XFAimIjjUf03RsHDZseqSWSBqgu1wr3musFEOcMp9N5UBQcSyJ1phcECEL5Qz
uReqwaxsVhpnk+tUclAe81HNNJ9UUVOA12bZy5DLrTZB4FXFsCGVdSmwG61c1QTovqKAduBaq8FF
m5KHQ30jdb4TRKjYR1hrmmBdYNnz5LY+Tw41kwAU0sjP12N9uOwSfZMRC4+bxc8de286Vu688or0
SWx29hPVn3EL2qOH4AGhLtVeA6AuIEXlyAlxAmJpad+5NZGy7xjlFUQZ4e9RaCvjDRl5T53E7fYs
zO4taMAVDW73Gff2zlyKiYtjNuuEp6otVFrYt3uIRRmwhmP4ISuRnpAvFNB/NIik6nwOtqBow14/
Wv2l1jgd5FJJ2IcbR2Aur2Pm3psohs6IRUvfGJKLmFf7ywG0O3Aki+MKa84DhkvtK526BCnoSANC
43ddCWdzpyPJolsCiFwnQ5oXFMgDukM2Az4PkVsUmpDO7uxQVjFH2yYUdYiclGurjzLEsIKyRN9G
TQAOvVLi7bjPwH8mqZ8gk8s8c2d8LNODQfTpimRSh77sauHoATWzq8DUp8Ou8e0V7ITp3TtHxZSk
VKhsjWb5cKJbOwl6xexCS5wTiZRCixUbAXtHm5NLKTvscED0YEm3tQVyxkw4DI2OSZEP9m2KbXNg
XOzIVJvNLu1DyDIeZD14O+eAMfOYiZjnzG7MhblZWwNZmwl6SZR7aSpUVfB3mrfCWVSCzv4mthVx
o9/brNzGR7LoK2SrhjLMxYLjqfr7k7XTThaA4S3O6YKMfyF2BnRHOcuds0vu6hBqzDTYzWGuu7Nc
LGOBb3rOoXTE6XNxNYPO2BRSEicW7Ccu/ataMi4wiaqzbMFDbhUWWToE677Qk07UQkzsgNourD6o
FbuNHnq5Ng7DDC1WvPwLhjC3l7WS90nG45JWvwxgV7SwWZ/OqOonlCGVyCK/EKRfMdR7fQi3qr54
buAvuUBE/hsoEFOpYikouNY6zoZrku88nqKCBNysaygGvhJNUFLXQEwNJL5lilazEpjoqsSXtlTq
jr6hwA8+qH47NKiMJ6rGO/iUDgNeZM+5JfQcUHe4G+6vPkFMlrC9hVdD7JARWsrTWkAHaZqkhuHN
9DBIFBSkfKF26oN79919pAkuvQYW+5IybiXFT2ahN2tIORd0y569QT1Ma8W0keTcOFpcr1Cw+9yn
tdDASJD6fLiyOsPpdyexZhAORIaUY8cKPBzwxE0oWlPg7tyqpqqC7KScML52SRcsbDc37TTir3eE
oA5sqZYJ4Vgce+VPdo/FG0TB+h1xiKlpPnDMgrCjH43vXvTOmSJCjYOjg4yh/OQ4fhYlbhzdA8Nq
0ILTZefsi7kGRj0r0ZVAcqm/D3VCwtKXIN+4NFI6/Pjpv9ulgC44pjMw/jNP12X6SkDVlh5f5CPs
sQEs4Xvloz9PBlvbTNsIPGiYAcdB+0mIYs3NEZn99biR8FxH10U0IhXwEIMrRC4auLZ7yPUlfZG4
yX0jhiZDoqeZHq6bMD2cNySY5gheQKFUQARC+QYjN3r+G8+HZjG01V47Gw1Do46n4KN9RkIrDAbW
8ExjxygPL3aSpRdJrlndS7hyUnVUn1gOhwf/1E3ejcBjJr7M9C96R1Y+qHHgTi7/V8MfllwF9UgI
IaUBus+fw4JvTOf/7QfwVV3zby6HQLVb0/dtfklfnvrr2+ijhje1JBDJMuyi4ZI0Xy3wh0EQiKVg
LOeTs/uhMTEi8ObInMBsi/Z4nK0gjDbkpyOrN4RFw6nL2NesRq4AxcDCVBoK1xdR7jKat+JvWhHC
ydoy9oFJh9jjTOPIf3i+pOffuYJOLXYz7adq5yMQX7AYaDoNDuZHcDz7kL0IWxIHY48VvLbBhecE
LavdSdovNfjYFJxI+xuhQXp5oAZnqsNgK6pUyBiW17c/M4DM+/CxyvW6STDOiEeM07oxcYVmFiO/
CIGzjuSsJ7H9HboSQ/yyxha2SugqXMl2rlpbeYDuHnQw558DfM+ltuSRsLvim+v4sSOzvAV5rMsv
99XaiCPtz1LM/ZmFAzcBz1j8jbyrp6d59rDbJZT/pmP5CLwwJaJebGLbJq+hvZFvuXtZiuV+SeX9
Q1hpmNRJUrrZe0vaB1XoDiRabjSA5s0FOP4j1uxDoRU62yC3AETo4fDuACjBql6+U8vqwafan0SZ
kutdsx61t7gr8Z8v+DKCdKSsAfhVgrZ365KOJFyfppZ/3e+CCbEOhiQz34ExMGplA8QF0HEKr90T
6R1fv3g/yuawoM1lVjyeEh7UP8ChgFS70hYy5qmOO2ecBBKhnhFJUb8wpmlKqTYrulC3mUAsWD0T
msOXjAVcga9QSKK4Avdyo1q73fZiTNY31OikSevghrGRoH6HZAdzFfRP1EYeNnmMuDemUUPvb+NI
Tk+xQOHCq25RA8LRh+JTeIPSLTmFQZ7zpUZSh6V4oBwoQrZdBQkLddD0tluPH/I2aHcgqw2YvmAb
gxwy1H3qBUvnvQgRK+nFjfKegQu3bAs5weoQl+oJTGL1Q+tiAmvg7gt0nhVCTKqJplQWoCkotSt6
U3abJ9kaMNT7dTrJDYbqOKFPidORuab9qiLPvOvsIvR3JAtifncOtz8Qp7c5YJtwRzNSLZAfuNh+
C7zQpMY5xWP9KqdiGaMdwUJlQgJXdTUtp5cyC5zSeL8fJcyJ4Ik5b9Zv0RaK5L5xWJb2mz3omHz9
gehhFSQDhNWiShjYFYX5MatuXKIuUpIrlE1VJdZ2w3qKIoqOOvUVMeLBQt0ZI3cuOkDjvnfZA9be
HZj0UWBGlLAmE8xr2CWJfo7n9n0pNlwpXfv40CDQ/N1zpcIYD5SYyW4ra6hnBbEA3cu/tTIuM/Bd
uZ3gHVMwb2yPaN/0IO9l6kXiDoph+BxG2b5SrHCl8vLCGYNvAgNXQ8J0h4xjJ9hp3TI+tZK0lbtp
8uP5bfPZyNCMEPjra1FDTagXqhMwhxbjyGeh+N3mr4uqnWadIDgwBhFahWSikQvoAC9g0DBnnsZ9
nrCVda5C1co5b0311RzkVBKVzGn3fq+1Rd/Su+wGpoAATG3rv2WqqwJPqrFkukBPaalW9OzEJaSv
pkvytt0h3tKoi+bztDMsJVu/V44nNvOLGEvKZfMbrgfxRCUiGHkejjjcgsWNhzrE+PrqlyU5KQOf
iy4etTAt+18E0NGAJfg1BYY4GD6tE1vCmBQmUkfk4XB+MyFT6xIp6/ctzZfM0i4Vt/uGjmiewA/g
AGrbwGExBJJe/+wLxD0U1vhHV88ET+5PntOD2f7V8H4IDx4HttJ0Jm+wc4vByrEY3KoHRyG622o8
W6FQJFUe7GZ+UCswy5Il2fYh/JJO7jj69j9jAxUuoYaOtFaKn7Wiu3BIjSRxfvb6mGtrG/i72mAM
EjjxH3u16Pg6qKbpcOPIfij0AqXh0WK4LoGUwgGa1mzDSREV1cIEUEDdvaxcj+H7QImvDt6HCJpX
eDNHjrw+/8ve5dvwXrPfKEp58AZPwtBAQ2bLiC9L0t7SO3Mp1FT11JBeMeK9/tYlW6Y1mO07zw8+
IVr+zdGZgQOAK1fzclaPbFNAP+TxBVG/gW8yCmpUOwL6MaCHHREXXI+Q97pefbTfl0ZB6bIypEpu
wFnCBKQQrJJlD5iahDZmNKnjFSVk3qPn3fO2GT/BJ/XUixJfZBLU6onbgiJ6944F2oquBy9dmX9r
dZqC0Qao9wrW7993h7tRt65yvuTg0JM7GEaR4hZw3Scxdj8r4sXGQvReEHoSiF9HrGt3Wo60YA3D
aoYooeLKbStYeHdzWRYKhMSv15dG2Vk+yGQ3tKPPZBzuo22ufWVm9KYkhQpr/Nx6SSM6IRE8mlwi
XOwxVRNzygGM6HWn0iYDWQpeT0xZXBjoOWf6RW/vqLa802aaggu0pg+ANSfa0BNTmm0b1Ug89czQ
mtuNO6TMsbKPhOPVMT1n7NlAwXaQYuD8mbq3Yvwv3qyGg/T7ILWJnWgFl3BI6Mh/XJ/zY8zf0a6W
2VSgjgUnpt/Kzx6sAjC1I2uBS55m3HtZusKUKVaBUV8urVHfeD7lDIuYjrZFtKn3q7JKzDD7NMGJ
Ob67A8PK68FaM8wJU/nCbN/bvgijAc43VnqlxURmR6A63dyTzC6+i1eEVVxWTT0da9euoPGn/Utv
PEEwPHm3wAZe6xx3czf+hhzjuZpQSFZ7FxBanfWb4lsPdQJi+EMM1f653zwHXldg/E9SwqY3trHd
ALf0J2OtRpeY5B0ku6K2xE5Ba/+onGjumw56ZqNVPltkcYYToh9q/btxsAf5et8Kge7EVqGw10+t
pFNL43bSbcA8kDq5XQzmslEdxy7U7kGfRFLUB2Cn0lgmSdeen/m5yvs6rOQwKkdNSH8zn9dsW6wD
WEbgucX2dwV7+NUFf1veETJXAmodyBRVo7Dn8C7iFvY80JIPDjYUkB56R2hweKk/TAEEOfCQfDwq
oUtCXrfMp1a3Z5OyquRHT9stAqH+ptmFpGfS0kQCykhiOlllHAHyqhkrHDLR0v4ISrqBFu5w+wmA
8O3eOYjQaZns+YqqL7jQOoEgL4pZML3FchU7MNr5nIEBFZGAbi5rVZLXaFJz3sPiNGI0tqDoY/tp
x/0I8s9sUFyZP9jjET3GAdfpBjLwqcgUdDJaAdoYD6seVoLa5mAThWIfBjuCYct+MsqDCDdsOWUj
ZnFKuT1EqgmYfTQ8n8q34wArG5bhdAvluW7kyqXwK2xd1RSJm9bxsnR5x52SjO4WP689ZG+O9OoA
PGeC4bOLz8EWLNw0kHdC+qESAfJ/wO2PZNsgwAcCACa+y/46G6ykEPY3ZtxcWeR2AvLQ1WylS3Ja
EASu/XgaLixsOyfmJPJjPFYwrJRPJV4fNEJt9OrDKBnfsQz/dSTg4nChGZ3n/aQyrwPN1nBQFtbG
F6vscvw2hF5cNz1qAtoY12wl7drZO3FQ7XGCex1NEzlSmJZZF7rkYUCAMNBaYWjSk4Ch38MZhaN7
mfVplbcipdQ89YXRFaxO3sJomSqcuSqlzIoWD7reBNobDP74Lw88cU5bPqfGmrcgRd1qBmUTZyXQ
jAmIWniO+qZkmMheUMSGUlIyH+p7UaNnvAsDivx5oMJX3jDZZ8qooR/Yn1o82aAVomtIFC+15aBZ
HadUEKXPNAdpbk32FJyh0kflfQeQAqA5//si+WoWy9zjIO9UxlOetj/xXzAw767EjiJePJyGlyU/
mREAbBmdnTN4oWMNEv0zJZyXzTdZe3s7luCdeYoRkAh0zUe3cc05UXpOXzsE4aKiMrWGNkeghmEc
xi6Nr5JyggYye0adf8lsUj/GSiDD0xU5UqdVKaymmSi7pdRa5xt+a3NoSvrXuKZCh3rOK/vSz6o4
dulBfyNu96f75nl9IvTvWnmRvFtc3mCDJkrUR6sP7IYn3HwfgR3YGJw/oSqsJJjqzJn/hJiUYgNh
rfkpH5udrMaYS/9As3ozgc/CmgwaELD/QfWIRBPee5WPoVjYgdBIlC7w1mPNeLuJjVF9fSU7VYg0
uSdNLZgB0ZsODQt3r+bYUAOup7TvFGg9AawymqYESw/GdZnCBheSLPKNQll6KJTl4Q72AjE0DCBC
WgPoai73UbApRarBAFzOc8fhxRoQjWZCRka7vMO5FEn2wJtnL8/hN8s/7xlBIrlURKE6wPikjuIR
wJRXiljGPdREJqhQw65fu1PQdGq749gs3Whzu/lhNZ7qh+WC+urV1ZcTUuEMAjV+wUOcwljXIXv6
8+Y/omP7s9uw3kcHgNslc1+WpFy2oVIczQzLWv95oRHcMe38C26rRC4o/FEDhOPVvA/kJv4hIz3b
0AZewpgftFWGeoIm6otXJkM/T6kiINyBdZaW1A9WChR8ivH1Im3E6qsMQtn8of0o2mgTaTYDz5q9
zrW2ubTxgRB++Jl6RAxBr8hQFICAETrqPYvMRh5nBG5iOOSZVstyjhvsZ4N1s5g38idn9Y9Q46aS
2QCffEHFeX+/vtugWSQtcnhyiueuwix5rlVJDckD0CO9KRiRzQEvvFP4+c+ZbhVNXK2Oxxl/sFUN
m9uXak1H33Co5GAZ9dNUszc0s9Ra5QXPGR73yBsJ3/3Lsf0ub0Dg5/93W2yMMGbnGDf3imkBxswc
6LjsfyhL3gQ8d7S6mpLqKlm09Ocr7YJyCbJyb6z5n2/ZxA6aIyKwGH4QV4J34+IdjUuFufUNL72/
6bu+j8IrQnGgE8215S4qqIqnIS3Njh42iWjbDG1IzKSZiJqpIpPXXy6U6fbgrE22GVqXGSokz0nV
Agj1yxvczcnyK7Vi2EBG3TjZemFv55VxB6e75XD8tR2BTGwVNrEIZmY3GjirOGStdCLYQvUy6352
3j1+JgsocFW4vu5WrG9hpBE4uCSa35SfRmvD4dV8O3MtY65Sf6MJycXZlYhAAn2DpX0HKka2HRql
ABTxApVlPdV00OoCrWSOK3bKQhhjMOwn63jyW9K/DFlJSbYtM45MayV9xQ1a640SPr/wa0Xe4ARr
RnQWsQ3nhtYsXPTyo5yIeEY39xd389Y/gmO6YSpIDfYbDJFvZs5lFpX7x3bnnz8blnNZtoeQqTK7
Xef7uMUB0ggO5XNgbOUXOVR/vlNvLBhOAq8Fz2WGkIGHM/mJTNwZaezQ7S11UL5PjCZJdsJEt4yc
dFxp8Xi2wJNzXfN+/gIAriTAC4BTy51+V9DZ6YaIFDig3/fJk5xMfmzIHh4KuSiV++7EjicG/YVU
4yZpZEuNMTmYzSoBeAU6i5dIbngqXvuQR5UhUQ+7wbLAYXGnFaMwA9qUmNLeQndDbUW+4ftRqyi8
VecIF7Q9VnuJBbINsEgpPG0T620lIHnrmcsYxohe6hhaQd6rRPN10PrdlIQ9MHAjxvqC6o3d9QJF
MDZRXmE/+XPAhRQA2zRiWIQv5CwAOhlOlc6Mkv0/UKNO1/PY7kQwITBPHDervkqBvEb4yI+TJ/1t
YCFilNxueVc8u0wT/K8Thas/fVTcN3EU+hWvvkghuR5RVKYA61CaXBGrFQfGluGTsYoK1idc4WXL
g2mFzMl1t3STbId7L7vgTun/9B45hRlgItGh5ZQbkQkeGl2S/aY1XNFt9CkFodyAW4gnyKA9LOB6
cPWXdZwjso9srQ0/MzY7KQti4Y3SbctNrxmH9pYAhE3YiEoVlxZDm6lYEXuqOPnCuGmFgTvKbAv2
xtAt2YEFq5GijvH1GhuXKfHesEI7G6KK3yIPnxU7/6pXwX+XvzV/s8gZHoA5WSTE1+p/kqfpjPVe
D6zbOJzfT8WHS3v8aFmszrZJsv0fPcXnJry6B4zeCrPrnMyrcCc5l2SiH0ugviMFq3daDcHTBTpZ
7wa0zHjKuqz/EBehO304+pgE6fO7Z/k0NUw6ikgl01PPNYrNreo88n13UozWwNCXDXY5G1WnwUF3
sbXttU7VZJ5gLidkyVKNo1bFlHmJpLdBV/Ycer+131UgUAjLrgCUeRnknLSQt1owmm4xc7bqcEJQ
TuuR3eRLfdLv+7QjeDFqZoAjkH9e7ifhN5rJwBixgUqFlU2XbjkBq+cLDtc1iXESZm+ey98kh3VM
s/1jro1GD9xGDASBYPzyAWE3mwzsDtmG79xl8mCgGtX+vjdN+8YpqBLYRgd/8ANGquidQM8RPApA
7ryYQzxURCzMdzk0Zf5aivNY9Sv/1lmDjy25IgihT8DdSiC0tJLZjIww6qd1tIhzvwJ4PfNDmjib
8Zv+Kf4qIjduqynBN9KXUaGQtRfpgLPS6YicFn9EzHBmdqwqbA0eYMpek/Auw+AbNMailOOewpYU
DRutnapv53YLidmDYiQxI5bDW8Y/1XF4DHuG5ZZ19vM7e7C3zDmsgTfr8bGwP/pqmZVzre5ZkYVQ
AdvCsC3YoR2UU60RNQTQXBjibuGjFzuQf+JrV2C3L75TTolaJtEEeCPCGPfRyWpf0v0juFRyx/JO
aCa2V5LCYVdAtr8bpFsDKCq6snE5puzaWYMFBKRf13kNQRUC47+Kpmt6bQ4diTh1TEY70k35O8Jp
a9G52vMWuopqAyyvG1yZ5OsAeUcnhBgQS3BHYFKvdExuQe6p0saR9Emxd5XXfHEHMTdtuCJH0f5+
hbm8dHFDlbQdypCbgAMniSIzf3TdRE07kRiZ6SH2B03X5j9sBWxUkmiJKjXWqYFv6fXD1IHGPfBA
yCTyqhWwka8M0Iqf382GuaeriV6gVeJf5nTl1nyCyULXek3xV/yhKCLOEli/9l44aTL6d0NN0pWP
uxXW32NooolDhxIIOnMagqyzPE4yIryjb5zG7mfX6ZZztO6SROFJ2K5+RpDTaRc+vAwfMzMCQXdG
12vnHrxBQgT2Uo+576wQ4ZVAbFfM5ZYMOHmnbNfiKm5EznhW5cFmQ75VaOrPsNICvWArRvgvd8h0
7dCjgKEKSQUjgKKLhJr6SZbX0AQFq8H23DSj2HeTM94THkNLlyQq83u1eG8p0wHCtdswN+IoykMz
ll/gpmg10KciiyLTjdyT4u5vMHcyWO4SWR5HpUykn6RY4PtzNozK7Ztmmd+WPg9nVO5rTRMAFPV6
r2Bb19OVuoSw/2B/j/D5baIGsm0xrB8S+tCd4ajHER3kvdUDfoL33VbI5teRz5Q0RtvMSSV+0WqB
EdAk1vBtrhXBq6csolC5E5qmNusAHbWThTKcwst7WR6xvHIvkjO9CZAs4hFfEgAuR/vFbE/wLNvx
l3I0Dfb3MAmngSIY5tR9DCqAOOSA1IuaVS4kYXIfhRMjmJapM7vupG/IUWtOMVh2cjtVye6s3lbv
4XlWQDWsIBgdeb+fMCMtPEGtLjZHeqOj1nZBOquTcXd5rIrlFXmaC7ctuz+8KxWG6XI9Y6VF0Vhl
GADf9TDrBJ/gtd2agM7I+tzqZbnNAJF8qubinJUoRWFnEcBN++oef68GYdbCOyeF0hSemyQHdEL9
clMvSq9OP1TC3EqtRRg5DYAs6jOx2xknddDgtuh0G+W8wx3wZNKo/CaCzvEJhP1WjHxHEYrZoJfO
XRfTAZvMAeZfPOqKCNGZy0Zsdm2M5/yoXesstgcYEKU+DAvEETDCiEn1n4uf9Fzq3zJtjI+ih37q
7dYeB6/lwuWwM+/yuFSJOfVzPG3XzAwlr+aaop23AuWCQTU0fSuOOKgxu2QeamuqZ7opQxlGlkNW
+hRiKXjzYZV9GOqZXxjluNO4CIcNes4qmCTPK/VaJhG59zpXaQqRR8riJlznrj5SUbI8TzbVgvM+
p1bpx2XVZBZNTj6BgSG0WL27JxUVfqD2yw5ItQmne0Sdlqiz9vZd1T64q7TXv4nrQWULOi9EfAuX
UG68/bd4dVSCAfh9LdUVOssm+iyr24wfwZ9zgEYAysnBKVwXkLu9sbQbM8dDdoGZFaXyjl8dsXgu
tkFwy4pMz7WI/4k1o+zOODpnyrdds83Uh1kb8A7emB3OfiwClSV3o7VlBuqVIdTurNd3k3AKc7rQ
Izb9oYTesIs3BwawpvQqJh7DbtHFGQYvup+KxyeBzy+deuyna7VK32kRlWJV4HDAWpdeq37kC6eE
MOemIGPhkdzRetVXnBertBdv6IEeN4X9xwqkoKUbzH1TcIDk4I2P9wuPy7C96Fuw5C8+NgOcoLI0
nNJ0wly74dh28UISLXTIbJ31TTteDcaQP5zpvjWhPXM6zpqwdBH/WRK/dV0mzBeYM6fD3Oj/MPG0
d+dLlIYvBKlVOuMJ67MBX+F4HJexi47ECb5/fucCzkCEiOR6rrD15igDCt37kBS+IIaHehr3QBu9
UzBHRvusL87ZGxHyNZYlZ4BQK8e3ceVeZ4sxC83m6JzHdcGfVQnRhPXgVzoJ2EHwyTYlqrHiWy9Q
7Yl/IEq/TP40ynMEukO8+A9bdaGXw43KRVtscQGhPzQvt7KJ5n02mFTRYKjLNlRs/lJWKc/J6KOy
uelay5lGBWKpCjSTykaM0Rs2cnBVpdySG6MGQWXwAp05soYC6UxBp7rxSPlUVBu6aM+gf1t50+x+
vTKdHHoZj6iWjC8Cslv2YlGWznuY8jCwYtoA5ZYRiaTnVyb7r6YerzEDH1yguAeBmrOSJ2tkRKKF
h+LN1jfCCRPJOvLMqQmXgrpHQvJSl8/LgyRwPqPo5IKi9MIQ4BrrCNnhKDHBSCif8uRM2ieFBcKB
SFSzca7j7uvLEEcQx+mVrFkDIaZ849FzA5+q6rOYcb1l3yyc3/tzgOyK9H6w1ioRdIoo/8FHp+/t
+tDPuEDgmQVQr+cunQMKkK/wN6W6H+tKKptBKKUHMhHkT7TBMnuQM6lSuH8BTTFqx39MVnFN7BrN
Vxn6Z7vF0aWoobYOd27q3EFc7x46sgBj/YFvHYOiw+jYUkhoxP2ZqrWvTZkQMEN0+5J1M0Tu5lRb
HOKkPBgqxXQYqBoAZNsHVm9xDniDJPbjxdwQWuECxuC+pb9Qk+9ZLBiEhsQUkqgE+w9LvcenuZf1
Jt1N9P0Agpqrb8rO6fzUKpTMzdFZW0RifcqqNH6WEmXiy/ALs/GRlSJil+CSPEMEl0950agnK2t0
6pygIu4ls2gX7uIgEGoNOOM19zVRTph9feyif3Pi44gb3rW0nuHuK46ZA5cTOEnglMwaicbEyRcD
pSL6NDseGWGxZbtsnQWKeKhUJ13+Bkv0v7rzfWIWMIRxVoqLUnQ9Sb5gPrQcC/O14WbVpq1DS9Fw
rQCvrH1qkAYj3jmNr4KrZnDt7eJ0Yh6w4jiLIvgib7e6gUPouZJCvmxPl5CCzXiu7xiyc7k9sz80
sS7k6hArqtsOauVFRdqDRSBMN1NiGet3psyOwKcyJSLMtE4IR/IXZJbXTrUzLCUhiNue+Td21YgH
iTMgvazSr/F0QSZZ+TQcBEP0ivzCqNLvTvMSqXWYePQPmCkypQCnefpW4l5FP1292WRBwHNNHXc8
nkiIEgoRb93/9x4K4xAXfp8h3K/jKbzJQpUpzwwre8OeVOtQ/lktKMaw+tdKhqDhXL6NZj6laQ3L
9MypOWfIKxcYDOFzYfRlZyxKj/K/qkFZBPWiveaWv1A6KIhW3KROXkOwJRq2UOttf82FzmYHqVEs
py6w0C5TL4rV2s8ZMUvJAF9Rn/bjqoaFr6u52tza2uJH+1zM5Jy+1ZaClMYmBKjjDnRixhw9nx4a
4G+jEwlfPIj7fOMKX4SJ0ANSqkDtmQX+JFqRqQRZ/jCgXpIc7A5zLp9aBfowhOtAolkXg2oKlFC8
4T4QOC0d5jdiVvwcTxgyWewLPJEifyDrTQUoYutaAu0jvQ4GIFvsLmnGNcwseSPzkCLb/eflxcn7
rm5yO6bSD83OLbNz6k1gA8E9EA1v7mjbCWXCRhzujLzQG9LR7dwJJgzWpDhh2Orz07GZDtnNdoGM
acMuJXhxRhRj+b3AY+oN/XyEzVycQMW2sYUtt/EgNpRwZkznlGiOul0ujOo6HR7U4Vc90Xi7hmlI
925hqY0UAbIy93D+jRttdGE9FTqobxmoDPkZ7uX1F02NQKPhO7kl/dUGqsiY+G3m+XmJspYfR80b
anGClPh5qSVkITOOZI4bYtfWFAf/m0/rz9cQDnCLsUQnkUYj8psmsHX/CDFCxKq1FqPev5wb1aHv
R2RBVHk+q+gzH6zczYYhJ4ifoMCqSASmwpAoyNYXe8ZWCbY5c0NlwUezG9nH8OwzDhitTYYq4Vqt
dv+Cr0JTcmerbjyl9DnUGxOa1uYc4ZInkAQ7GQz9jBGQM/13eqLFcUrivGCECabAs05fIUfXQcYA
xIms5y3ezP2+P6e7d8hEODp1y5ytD2xN8xZC8Zzr8B+Gdqhh5xoVWWt6d5ytU2LT4Ba7QDEk+kkl
ZXDdw7AZyfabBtN8d2lqXnwmDnw6TupX+THYYx0LiS0rCtDSCSZjXj/eddYfmG+CEuNLLOmPhFr5
y4MjzcK55c2q+Jvjnv3mQmlJMnE4mlyRCmAEiXSZn40eOYIXwD+8xbEQCZhrls0mYnt1dGWjzq4a
qkaQZ0af+3c33zZFMcKpCkmQddtTp7eNjWZABfJE/WvY5NsCbHfKnxeDjLr6Lv0c8eqf7L5jRr00
eA6wmSp+WPG6cTORVhk/EAELFG3yn6bD1kDmYd+bykXiuK4v1S+Xz/1g3Qv0ROEwpziyL4F0kSFU
mmYcDeqM4Nb3esXNf7tuOwJIiXXf6/SUzD0cuT5KTEnpnkGIcAPKJaiW7Hv5mO5SZVP/CHvoWeCC
8HI1AQx11ry1Lx2S9Yog38euZN5xoEAIz4f0zJ8aBeNXUtBNPo5C+3xgkVDPDGJayCE+oTheDD2q
Zp55JWRHd9iqG3X4/NPNwDz4uk8SPbTa4PB+lATu3oSceWxZVzBZ5/o8QUQ1e+msyICPVK3CP1Jt
XiTQ8u2+R1FgAOUQuOEstXJqGXpf5TrmTO2GSVggAtQPL08tD3R4weuvi5eMl5bBZTTZ7EE22t00
YsokfGdQPP4R3swbD9g/k/dC+erCyI/aRia2OQ9k63/F4vF9xhl5ItobVtbmR7ZEJsDVzwTkFyDS
6aNBvqGViB8iB4l8dm9cjMw2KaFr2eymqenFOABB2AQ9r1eE7spyYeZPgg0R35xSf/u4KRUcCem3
wbPnSNP70wkQn288LQNeanygfO62Q/RQbmoQGhx/rNtbjhelU5/qq7ziP5sYX5rDhhL26hg/DkBY
MS0L7O0JfSEMP/VsIdOcca9/knHDtrWP09Zu0eW2uxvtPxHc00euzZCvbnZ4gTo3lkCQk+c5bQ+6
7DPfPy6SaPnDIKd5MzYzOk1hW9KhbHguY/YeYviqfmsLJm/9MHSVJGdwZLFVIad3I1MrPfQXUwDH
f42TjKXMufUxOf2Sqvu136cZ48a+OwOI1gWTckTqm6aosjT6IqPU6Y8foXMTQdSfOb1c2FDSCczg
1++Sf75DYjBX8vgeRpC1yPG7/bn/4t49LrSzXjPFZoZG1vae2B9pet0vWEiRsXPJ/mGrEGaGJHAy
gevjaniOO1iq0938Ai+ls0ebQrv0hhQ2bsQfInza3A3kI8zO5AkFzihnEXaqdfqlF/koQc9H3MJH
Eohn/+2AYbzOcsMXnfvG/0UyNmrSiIH0y6ee9OgSwQSxYGWyaYJKCkz2hzB4LGb1hx9B23/GSSa5
Knv1rjIej1QBMyRAbYl3+ivl+NHKvP4kXjsa5c2SAg9hOSyFnuMxPzjw7BFUOcxzEnbHMJnjizGv
JD8S9txsi0ZiJY722xxURyuEbBsWJ127eIrFjz0zFRdgAYRE3+5Mgx3ga1nJKPKTEc9AxuKa+d5/
C5wWySHPoTYllu5LiBN9sx8WUwz0GuV5/yvnzei8kaQ24j6Z1Da07cgOCHlvyCGIkJRrzhrFJD1Y
xt9sjqdTTecqtA8XzPoxc/Y4mJSJRi7KCZHYJB+vXud1GzK97EpCV7rUN1INuIiqrOmIcDGUnTke
NhQImd3DPMpSWBQj7FSgru/5LpTGIdmJYKwBRJur2PYs0JO6sluWMWhVn+EEKdOz0KpylCPcD0Ka
gxXbnIgkqLFeGS+0sQt5rKVWuaRZxv126bUH12Be4NmklbM2o9gQZ+bUAaBE5sVTg0IGpwc0U/Q9
dTAyw3vvuiQgSpHCPcPZPVziyokHq0nBjCHrMA4u8g28xGFsaF+FXV4qAyhwMCcbOCypJTtAPoYD
5ckgjpy5ReXRL2UuvTNZHjQLGVbRDGptMD4u02g7XFfe5KSNwggOK6H7MTaSpw6DIdJiT2Uz7WUA
BJcOKAuMYfDz73ur722CJBVuOe/36yEA5ZKTfPye+94cBeAZCauPpWXGoNR3imnSFXv2nOu9ylAb
Mk6tO6HVHZg7WXHH62EAFq2Hc3siquJeWZkHGllIVqIY5C5Iz4u7PuGhzXFQcpbLIEzs4WXd65Cx
YhoHeRbb5sB1RTZmy0lmd37JI0IiS966/Z0eTC3NSSL8OHmaKgF5FsAu0jaxjmm8F3PwjzJE01Td
7uoSCYmiiJ9ncwyKGJw76BitpmlkNqPqHJ7Wm5BbQTwDCdoBOhWwJjOZ/f6sr2jWPXAYw1Nx/PcV
56PVzZmPf2q55W0c7otRM/gIpTgrObEP1+YE6ubM2jYPRPmirxh+MVgdP20j0qbVV8QxcXtxH6dr
Q+SU+Za6C5EhQ+WBKh1oJh7+GQAPERKWkYj7Pw+tbIItqzy8634EijdXTGPOdH6747wm7D3+N+cr
Kv0L39lFg0++nQ9/dTFjVzYPLi6Zow/zFq7JwhDjqmGI0Utf8/MZ8+97IssbBKiUynEOgCV34RQj
nKtLYRaciOe1crzNgQgZ0z69MhBDeaK9Zh5pjppWYRr0/kyjJpwFC+CkSApeHF3x4CaawoVQVGpD
AbIN+y7cOvSV8GHSeowqaWAUTQBrqM1lwkCGsWb+c6T3xuRl0o1qy8I5qWOmJcq0nvUC1GbtmbyK
T3owRy5/gQConh+mIVnMf3tLWFL/PU8dVT4iT3c8e7xbpEj9IeQNQmOh27+Y4nNJ37PwFjwG7KHm
hFQqkWCjkySlLFDqN6KhQBTnTqJwk646uOEOmlfd1fwX6NSJKgHh+rr8fmZDuFs+ZzWvQZzwqzjz
8eiyIfO/7v+hFX/8Bi8eVRAm0gYThhGtKL2/2idi3oB86XnOXvALKmwIAZumKqnkO5SXfxpTRwyQ
sLnX+DFlTmv2IvUfDps5us2lchgWZg2LF4oa/qjx1yS2gQenhFNwtQ+tSAMQ0lBwWKcpTXiFijNi
qUqI9DfjlHXmaMAPHIPHu3ITd+B3dueAH2XRoobS9CpnrPvLufGKs6mEi+FPKS80j2Tf65boLfeq
c7voZSAj9hCgcHMLq/KvCulEi1aaMy573bXAX2QhJOd2lKtydyAmp8xPeB2+41byK/LCQg93e8uL
69R2fZ7CFPgLceasibpFiKtZPp63TRAr6bNV6/fAIcabQlfxPOjPFKIITDCqjD+WPfg/7YXjlVZx
dVgQlEFZA1g3VaD+XmdUD8tGgWlt3ERaI+5MYBpavW5wGZE1t87dpS1eo08oY96xDdOq3BXYSiFR
y1lvi0Gxze4beKFlQOZ5q6HFeTyblKTYKwQojcvZk9n0xOvMWpU5602JNkupVLayw6BjpitZkGsL
zVpr/nH60sT4bt/gdzNFr6NRMBE/thT/8NdQE3A2MHnGxVGGgSfawEFkWWqZvNYCZPx4OEWYLveQ
iAxd7JHWmQAYwbw57B5mcFyNWQ98aK0voqMg3Ny+y9L/6GWZehKdy3MeRJ9cwiehpCvX4nGgHblC
x3ZV0nSBP4U9yyVCJE0MnkUreB5zWBdvTUGVvjzaAKrhytOKXJ6no+MOsrKtwWmD6VbtUxuELdZw
8WWBZ9ZOlnIhflwQBNvMdwRrmF5ym5MUNFIlnHvq/xL1+okmr4jyWyA1bF2vb3T/Qbugrb7qX4gA
M+a7Fin+UCLTDLUiTPIBqVd/f9Mmef8J4N717Xp8U6ERh15hQ0/zRZORGlZ0gAzGgRHsBnEMTKq3
hLtnEWGRdgASnspVTesdMgrvsmndSbi43dOa/0CKPlwjZsxMblOcLKV6ScnOouDmCjD8i5wiuXYK
kN2K0hGlnLINtfoVlFoQ9lKY+8zrpWWzyCnxgZGnYEDD9X3KG4OQ/cwwfpmjtmqm07fujOSXSRNH
AROa5e24kch0LNyYveZEpEpThoqWWL5L7+yptXJj395FF9rSZokxOVzHrmtW5wGcryS3ZInm7nHm
ed6OuMNAWu02ayxBGdfLr+VcnUTOZHopOdTo43TG4HZ/HUbG6NKoiwVMd2SbaJS5Bu5CzQdfF2GL
LrF3SCLvYSADAd5VsoJtVmyduzDWFplQIzDpRqVMPoZAKOWjb85+2AC3tBEqqLl3uAb2o2Id+rXS
K5XQn5fjrQEGfhiEKdvewPU6yOXX1AK04J+lYBKkBRjZZ72AlEWwvwSEfHWT7GafRu49SFs2boAL
Qvi0U+weI5R+32+dgVO5y+G2UJZWcaszJqv6WFu8X1sm9ND/vkM72ORFyWUmv1LQYOoq+IgqzIja
Oh5LVYpNhBncKczv4I8HuK3v+qoYBHYPVjp0UATacUhxHiAVMvXGGVp0ZWtvGXVMz9mVvHJzmcXn
mbaqj9p1MaOnVO9D/Fv10Dr0OolJx+Tmuam+6CJAcHDL5zNUyut1Lo6jxGdFEmohkX8DylgLmLNp
G9kErMXAm4v6MENayhZTAAK+SWi6MM1VkRWnTn9oBJmAT6iE20K2YMhd20Ft9lrn5lMieROju80h
4c/wJs+SbfPZjBsK6fIusuBApJsAc9ZACDqW3TsGbgqkehm/A7/ebXeK8P8XmXyRT6bGqA9EzgWo
p2G+Hb/lvZkcF6PxtXZBlen5bhg+mDcMdeTLKZvTSxVQZuRJQQ30g0CzTezBSdCqS4c95c2mo3hT
lJHK842cFnY4eIBMMCmTS6M4TA7nwsPxw29wSrHEpw8G/lPjitX2maGM4K45hRxMwpowDccd5L+1
A5FKYQOsUWrlSQsSfMeq5f67bZrMryfZVPgOjai/+JcIqeu+T6q07kh/9iuml8PxVqAY02Up0MDE
clCsWJ9GhjSI+YaVr1RgGylA3fSGeGZo8GlpLmR7CttnwxpTOUHrdNJWG0FkF9KHw+uJrimWxYxQ
IUIu0js4K6RR/YTA/VqYoq1oWkv16Tsn+AQwR4OXPuvLaw3XeA/jLBxR/h9tw0A2NPI2B1izuga2
DAvZKayDWgohtSDaNn4SMUfiGSLKfw00b0eTlgG/l5WFDfu8HfkiSZ9BzeUVyKPmOHCmNQQGbUlC
r6JMf2LoZiMZx8xMYkY+YwXluSQdSN8G9rTl5aHi7WZV7y/fZvavGyoDsVI44XV2FdfxYBuv3r2+
vwVGThkYG58MECSifrB4VdFRDz8ny16JUDrr6XPAEtN4A07XgEQgM3s4xaM9jb3dQa35WAty7MRQ
7Q3tMGmeovw8krCDCcD7NgEskFnRTNkAQ8X+IV6RRB2b7+N/Cc7oXPF4yurM5a/gbU7TYjBCc/9F
ucRok+GCWnXXsYOC3IM0nGPCm0Mw4MRa2o+OJApgLcB+PiY7TRMaEfJyrb4AobEwHPUb2sRLX0ob
/9g6yudmXCCelMt4vncHpI2PYJGGtIq6iflNt1ee31byfVTTz5bg9ARaGqo1Ky6zIOMCnUVfbLgq
ONmER2LMgD3JMtVqpacgicWHrHYh3luwIZI5ETon0busM0zHCqQIhyG4W21lHwKnFHa+S3zIkKv2
X5FPIEx+Ts2P71c2WSE3aI5hG6qpej0fM3gEq02LtvQhJ8pDGbHpmM8hsEAxRySxa6h8HPdEJ+mh
LfehOt7snr4JZZTgyPTHBC3bp2tVTsc0htGgWQWsxJl0eGpApYCx4o4I8Kmh+LW7LKiFkOaNmAa0
tGSt0rikmYweLetxb0ytcR2GYS9NBquf7ExYLnED2I4GeLvQuiY0hC9u8qft5Wta3aUhkzca0QyY
OPiekiz0OS58KrRpAlOSWZRYqrHGknMzFAcah0OZoJbyK18dzLS56d+NlTB+d5VP1RYy6ijkJBRB
iEk77j+kuMD9vGYcVlLG4+938BOJ2cG4B2D9ELmJ/lB2Oocj+fE5GcetVzn/Dg8NsvWBBRI0Z19Q
KQF0JYRQYz20Y3peLb4ePP5cyDVKrqMHul1Ing9XfwE8Ajqd819Gj9J5X2FgV1xV6LhogEclWRZF
hfRPvNfBYrbWZRNTMD+8ENkcGtHaSb5/AqrN6SDXFdKkmS8sK6rjQdRkw0SNQChVI6oYso1oXydR
xS6glf0Idyx/xcoz9WMby43umVK28/Fa3O6tl2A2MPYLXSrB49tyFiTXP6jWhLOu7OrRxUvKVUx2
uyUk5GZkDOs+w8LYqV/IX/a41IOOQFpAXiImJXd0DHp8UpHGh/kSs33+SeFsnOJGVcyjPPWsHss4
jEZ/JKH8wAeP/gWHHpfdku4OD3Q3HsTeCA9JYvhm7hYQqQTU83YE1VdO0MM9rLUHiq+VphR0OHvh
2fLwcb+CELkrSP+YMYQiUJ6hzleQTxodNVCHfZiJtvqp5rWN7G2mDneJKVp1EsF37AgJ20+CxEdF
0sW6soGpQTfnmQNLP4SbVEkWCrZpon5ikNDvMR4cqxcd/PwOmcwi8Q4M8OIqG/cUufhVgrfngMGx
9zx+Ho/oVVROz6i41sCGNSYBOIvCCIRoWHH26H0RdlcVHA4X5Ue6OKWFvl4J6TFMZ47fkNUMzihg
/drHT5lBd1oC7GOzN2zDhnv9uH/P2sAUwa28LpbpLgQHFCyCIJ9k2zZfIf9XmmgD2XydJ94FOqcD
qaTxLA2GEU6WYon/SHNtcxhpYzmrbFSudUTfxsbJmaEHjwdndcf3Svjnju2XD5BLkzsxqJkRpUw1
pxGy6btpvuQOaAiDnG2nhVy9GYwdJhdyCJM+R04/Vn/w7K4xIt+4aog1hzK3yeV1cLzDaKBGPQsu
XWg8/pu79DiSmddQ9cbleHoBYq0ARyQnPuwXa4wJqGtHTbG+3aY3U+e3qzva1Feg1SeDbu6gQTq1
B7ix9jgqoHPHKiMGdLY2VuIgfvWFbll19Y3a/kSLmfqZ+X8wZprlPR0nSbgB2bwpgIoippzShlqB
q1qeNQ1JkbxR0VtFQ3kTshKc1hlUmI82vQIahYAHFX9VaOePqPD7n3FeQPZBxMu7rEuMpsvqEMu5
yiS5HhJkGEum+5dlEgVfU5OMQEskLEK4qtddYX2/Ma6Y5AalK0SCwKgyGhMyRGvyNVDhRPYedzxb
XNkl+PhXPyYlwpSQ2cr7BvsHbRj1OcxXt6oKuryMuTaApg708jL1aMxbsL0+nHReZf0c2PvM1GVp
0do95hqH69mZhh/ohwPL79gBrChild+3a73ZBlTQtDxm4TQdHI+p8rPjGJx8xEQhLInKDjXWOzRE
Z6t+ius4wKBBu09EvljQytZ5hnqLjCvJ3vpVPgDHiSMmzT/+c9HE79cD356HI1LaKn+ddvCodDs2
8x9HLHB/svFwLAISuRfjU2jxDj3mAaz+UOVjFSZP09qDjt1rgJtgLJl6oBWFODgTgnP062e4Qpo9
0j4DJw/o9JbjdB8WdobgGF0BeedFRw0Oas3uhCl6Ls0gkAyX8K2ew0WuUYqOv0O6NxZ3E6wpSO4O
EJaXSHED7TrWwT7UhJaw9xLQJhV32TD64YYb4e2B6jYdTs9ukNKtJLPhe/v80noTPZR4npjJZ+o1
YtEBOHs41Bv7BOX2DduidAzuy10PL4gq9jTeXTmCLQvxBZ+J3r6iz+N9pIpFoG2vEi3TaMxF4VQI
LAJQzetwnEj2uiKv9JnmRR000v2BlFXc3rgs/lwEP5yukEYurM7JPfHPggDHPJ0PRbER6+2sVDt9
QLBjXctXFUGkrkQ7fAJ+UpsVn5Cv0zhu2IIFvZww6Cqs2hfABVikavYhDnBRzaEaDano9wDBTUm7
IjPKE2H4slXZRf8BDL/sL0HVWaO3qwhNPSo86cBfSftlJS8UszgA5FgT78eXQnghEAk3CaG4q1ry
bKyYCZfnsT3fEyXWaEuv1i3p3EmUZoENI7ERmH4x1BS4msYxwDvBVx7HZfk2lN9lSuOej/PbTxre
dspQIHmuXUjSB/wBy7xDbyUUMAHoFgfZZbcqF08IAKZPfMh+nhQ2eqX9jOKlMxhA9cITK+Jao+6b
6EU8yw2/vOV6y1c5Tg/bIPuef3OQ1kTMi4S3PK8OAb+jj0ObMN+zAgkQO0JyGftVDkrHiRz3fub3
lbL/taYPtmSqKOQdu0zB6dL24RALRWS2hU1s//4tfBAFjbPpgfQOjFMJlsiWfq4Kdc473UmhjWAa
2s7Y+YaPt+C+JOZApeL2d4PgFZLh2YG+EuL2rt1l8NTWnrrVcSO5hXw0oM6SZVtiAlScdBd5JMWo
aV+/ETt2oZhx0LyYlBEKYmsTOZiTWflN/bRLmEnRAuMQScsoes/3ZyLFX+bsMWSDHNsj8Zsu2qTX
5TOdFn+9F2EAfmH1+YhL5+1Bvh9hva/8py2ZxT+uiq/vqwlXyf3zXbCvigrmQM5X+xqfbFsG+YL6
WCZAtdlMPRLH4E2KOoVKeX6mxHPmwQsFtz3Civrh3qNw6ilX0N+XP9GYstvpj+PIYiqAQ6JGVkjm
+6HHJzTS85ktq0bCZI+Fo5ilRipivj3SOFFejWfv/05LyPLHTQi+xisauWT2CSYAKz/MwRBz1BKQ
T7zC6MM2CR9H0fqitvuXDCO4IF4Gx7IO60nZKzhIoSR737+B/aB0FFY3N6W5LkvVmLLZXDM7nouZ
bRMc16tD/16xF3JA1vOngT4k4QfaPR9X2BPhXkXN40RSrP+fLwfguNlt7+dUzx/E64oQURAb/+MK
ljPzszaCLO7PoX1KqCrQERw1SsOkr1cKtbvZM2s+rrxt5iQAJ+gZ/8ncbCf7iennfD2uv/GN2dNl
JJcO9B7p+27uFM1uy32hLfonvLwMlRABk4qgsx1hu7hRKCNYfzelgusK428Hf52vB5H593CquU4P
lfl/sEdZpQ/nHUBGFbslEZe22rBaSMcUHJpRa49RJVImqcbDNpUz1J7zshVclwi0/2r3NvAajMcQ
pIDY1LhdAxWnCof57793qrh26dESQKcLDhWUy91i4jq/DV56qkQeTPGXlkOXSbVuwY9zTC+62XLE
0+zJxhTel3m5gERtPiHZ/u7ly3Cy3hYV7FY9YDW7pZKf185L/oKdKdxqsSEGjGaExW1aQmUHPjUe
Lv3W1NXAE0xeGA+K/XuVzHsHv4AJHbWg6HFNTjbwey59hmgtwp85TtE1dWDUD2D23Q6jUQQkbazm
+brhDyW17p0LL7+5A8MT5SDNzEWikvssXpI2giDvVMk+OygJ6JDPmW6d9iVueeO6U1raKLutncCt
Lx9TApz6hGja6YGkLNbd6MzfMXasRzSLMYg2SU6T/A5pq2/4qRzZ8RMpWfC2jKUeMija2+6DOfQo
Ga+jFqfDHjYgP09njFp7Me7Pf2ybxUB6G9Jx4Qim74z5NmaObwVRXJbIYgd+9KBq0srRqkkEhxyd
Y2OU3NbwQPCcGf2MvY+8o5dXkq8Bmf98QQrat5Fi+ao9orvO4u2O6iL6yB73YyEOtxNu0NahiTpc
IjV18H/eklMa/Z5WzgytNtfGovAuOXQrJuK4GMVXeGeHBp9wXuH3wIa+fpHmRq0/TxIkOXqs5+8G
MnhYkMaSTTczPQGizvz3oHc+XfqXDlS52ToJZVGyjQdpxSJOao0q7/q2GrS5jj64kd0/9XvxcJZv
BCsSrj4ZFp5KfH7ISHg7m0uejNNz3/e75PJ8RH2i9GvopfPD3O1A+ESN2ZyOMd4WkLdp94iJ0Rs8
Wg2vUZeqSEzRAqlLscWAQXXVBwhpIEf8Nfnm6Zuoo4UgzGj4fKyUxwsVooMRc/7oaUAkUx8LrIRh
AY858F3B2cf/y2WRNSMn4U3iXGUJ86wSx6qw0C+aRqcXiEgqnGNitutJ7S1lPkhNYVZwxA3310ve
zgyHwwtH0nwY3INa9mo0SJwUhSN4yUjO/o0t+hF+nflwxbzHj/pIJktfohjFAeyo54iOmv7n2qlX
RxgArnfecLyLDgC5Bjlup1Ju6pM/jX1FBosfwONVOgiTlOuY0LiTzrey0PVYSJFagSUhawjnhfr0
TwsJHSm3Um7BSCtcyEOvLTyVcpAZdTlZO28RYX/ebuo7JedRWbakZ1fHETfmFadGKgTfv3qYUted
o1TYtp3sFyeFfQcNDlLAXEFrtZrT6xXoWvFklVkpQCM+dn80kijvJihdJ/SuSxlREp5svCymYcYb
oQWEBQDMIcDBUI18LBE0GhjjuMI6Pgs+qXkX5MEDsrCogCjEukMEKgZv9woDjfWRZcz0jjESkZQl
TLfglD2182IxDlcZgYU+XX0SFy6dgfgxghZssnkK1+sXbECRdCf+MpQ30YyjDcGOgf87jUJm+iRr
hjtGrjlV+2f2yf4KR6IxjXIJ+fpdGZFB5bmlRBRBlpE3rhETySaKDI4U+8BdBgD3j4/zTzdFnlye
D3WcgeiK/uPGlmSnPlN62HqkuRYfQYTOvDYsIMvySZhrfy8Qpf48LrxdI979OhtD3oxretkOw4rt
XA8xHG9fQL2xjGCpF4TSEziMUReBvzAh36yQlF5mn8fjghxP55dAYvoon4D0NjSvv6JtAkKuPgtE
/m8XiHPrqwTR7/zoq3N/HuiXhk3zgj3854IX8sfrSHij29hJGVqxV0g9z6O+E7LYDN79yomAJWjz
NpAwsPkYN7bAcK/RHZSj6NebbocqwsLrB0Tfrs5hrnmGCt0k0GPg2wSqHRRg5oNcsJ5qb5vFOVOd
IXYypYwr+/9erBmJyF9H0DLiI29nFguxfd/q3uPfu5BzuvxujlsodVzFgRv9GCyKYkXYa5zCB13U
JG9FH1MLy9oGvRRg6YjUJdh6bgGpYE8QlDt8MtFW/ikCcysf5PykAN3QsQSfkbjAi+BaX0tYJf8C
7KpV0tAvs2FVpmjb7Xm+KprhtH5gt5MO2sUd9OC1LM3v9awMD9cEkzM3JHPXA5cjEpe8B3vj2kdI
RsdoZCntsnNVY024bjF3xDyTCeDzknM7TnODx/ZPdRJCh0drZiMv+omKmw1WjXKZgGnWqw/p0M0o
nFp7y9G76hAICtWQSf6Qmzv8B4o2OkzORr+16QZouj60GAQemolwrgXicm7VBGwkeDxaJIKX28tB
o44FhNjRJY/os0K/tZw5iifta8w5WqXezyXf+7jUdScIlXHT72uijK/KBjlpxfx2JfKJLXVu5jnE
tXsd/IzIi5dBwoprqOEZVpGDGMJG34s2oyppK08aHKk7xM8ewtWdDKC9usfBNIFQYKkuJm5Z7OA+
stfMhU098Sv4tcaCHFnQ+YidJ2sKL0y4kiQSabf5UP0US2oecvDQT8C39zohmhkq8PkTv+HOTbYI
4kq5uGbnYc5BMtomBxgnBcMFI73aqPoNZ9yA4NHIWzGbbHKo3IM05x+oQwvl0UMLTR0IuT/9wd6l
+sF36j7g7KU5kxa0OhYb1d74zdtbSH07RnryPdYJ3uWxlEYS3uqNzhhyYZ1IZ6Z3arRLB4JWTJCM
AvtdfgA+Gjzgwv7xqXyq0KaMkZEi59d+yqvrEgoZKjHX10SJBk0F+6zsIZmefGPQeKRfIOjPsTnA
kXavJCTophBiNMuNCEGWVRKaa9qcTp098JqoI3YcpK0dpmekUcWumTTSrgoGS+BF76+c7d1ZkgJI
reu1Y7ISuuMJwbwkxpjDA8VbAqkQ/RFRPxh6G22q3EvDe3kEXakV7qUGsQo/3TYnpES/ElOcVQ6c
9SRxKP9HLihjOPIzkAWmYBzjer62tiw3U3WS/hgR/MFMkoGfcaZRLmeOOXGPSZAC85rW7AWEYhVW
Qywhsw+38GYMoJ9gaYMmUHPsFdgsCPAm8omQ799HMlUaMjCtmhgxy4BJcFYV72CBgBSByh17wYT6
so588BSv+fuRWRDpvYbE+wvZl+LhmJoQ1wJ+tFCSbFLDV4xL+ERK/TVF7ycEeW0eXyP3FL2q19XN
96ce2yojyoeLw4lNQFAoUQJU7qCVpXWnibiFjUukkaXmo5QRBr4u7iswY+5Fwp61HvNrOBPSQziR
agSWQ811ACo0xbu+h1f/cYK+FDonM2FgNv8QajbTln4+KiTD5wwsj77NkEoKMe1d0waE1divdwdz
fGBHYPhW4RYiSqXgJkW7AtkGD9SkY1+Z9ZHyMTzPVdZbRVIm2i85w3yEwFs0hI3gpc4PhpnNGXxW
Li7Rm5lGpxg5Vhy+PC8nTR3r3qvK77XLv9vNokBzxcGAVSAE6XVxw26XOTM8lRZQs2FSnzPOr3DW
omz+pT8UcfJICOzQRECLjduZj/9k4/m+bQoQLPjD/nDgRA6IsSURZQ4WOrMKBVH4c6JZxE8KbWCR
eBFnyqzjK79PnN5x9xCAlVU9dveoO9aiwaU0tx85bTeGnBdyKtdL7Mmsh0CvYKZ+UUH5SaH3sXbd
45ubsSVhB6VW48YSNxVfWdKbsijKFTCfdfRlKddm6k4TVvwl4NJWUPp6UsIP1vWtiLcoVCNUnUr/
4imWKLWnQOyG8IyiEIlkKRPFv/lmhoqcSbfPkxUwJnwEPpe4q+xRXoBWThaecRFnIuwz9YZG2M15
NlZZVlrzcLtaz0EwcOj1duMNdYiawWTMylFnJ2+hmbvmOtfdrTHLLuDLUHAmvovmio9NXmfASxPr
FllvmraDrxYhcfInJaPXXq1wA6SK5gv99Hr1Z4D9a2EEykGsj+8wweGzguwiZqqpqHl6ES8YjupI
w6K4TclN2hKpvCCcnNIv0QRCdsTrw8UFaXmEcLx2zS8OA21lWo+DjLHVSaM4LSeCHS9udrc0Je4C
w5Eirqp3TrS2GFv5InNRGUR0k+h2Z0T/Nx4J11pZPeWihUjNqjtdwPwEOxnT/56HPLj/jnqe+7Ro
sSHdIAKQnvJSUD8WGjku8smhIsOYZCTbV3jU6/jZVihijpE/apaybdRxMb6fdHULUq1pvjrlWIq1
SZLmXtPeWJC1QMi0clOwXFKE3p0+O7DHrIrz2GaH8vsKuO0E2x/KDnlzEcp+Yb0yO34sEqzz1rjI
sZM+qkHolsjGtZ1ohHFJrqiY86Rt17Ic4Fy3agM+pQSvH9siyg2j5z6/X6vus5/O5f8EoLi/y3rY
Bxq5UCw6L100BJkcgA3z66nUMI7uXgJuWHu0pVB4a1/VQnGK6c2MOzsItYs1klC3sq8D3Vs9Oyt1
AyXdeWWYEj95t6QCidiMvF+tImgcNWO7VKCu/zr64pGCb0BlpWwOUV4bw7/aLnnrrv5F9+vvkvqM
h43Jh54UVI+Vb6+fryT2m2gk9h6CXsGMKgNoy6CX3eUWXf6aEAV6xEA6MAzAa9+3glg/mj/4dCx2
mjbH+WbM/eQa1Sy1F2OQ10Q7fyXEBIij1QgbdusM1/XN+WJGByHh2ZsM36prr/UldREcblgsSv6K
bxJ3aiEU+EXW45nC4Xy3husgt69PzDnzs0vDkk89bJ5iwBOqUjg1x9oGY6WDcM6eegfE0ulLumpX
4bG2lWVMpmCLFozy8aFoTRXmIwEmNIdYTlUM/uEofPKlPfkE7dBCkZJ9/PO8fY4QbdFcGB8AH66Q
gxDjISliZAU7I4bMorAAm2MPXV4Do4kwn9hnGNW7SZIxnxYnPOWY6Yk6hUk/GWtVUP9aiSvfktfR
f3n0jbj6Tmu2yH9+zNYLQrSx3BL6B6P5gdF1feD+x58yEo4t0fqnPN/vV/SWkUgbAeOz/kjuH9jt
WgQSBkZYv4p5jkfZUIzzDQgEy/KRnbeHhEHdMQcsxj7AIU7rSNssRIaRelKlcO9xR1P1jQYOVZ45
FWC6+T1ODmCmD7a5S/iWBOHHP+rQA4b+KjIjvrKbt2SL9BeKoeB1FK3VP/GWcdvxFvImvRyvanWf
NeDDMT5aqWW4wD0JlvULxNe/sojK5BNRd9ojBBCkLpEydryZ+0LPjYyi2mn3tnmYwidNGM+LGd33
KtVUqHHKZWzka/1ps+0Q/1z60c44Bt27qbX2ssFTU8M3j61pDpeqzz0B2Guq7W2Ty8AE+Ao+XYP0
1T/BVS/pvtZDUa9YikVXdj6kR+3akl7qS686r32ng8Ajl330Z8UwFU4UCtaZ26oTOyQO5xCpPNHX
UmfJls4DKY3FyTe2wH/EoRPU4YgY0Cvj3RFBkesBG9xdMpDgwarDNQUBPdLn0JNsbc9b7tmgoSyT
BRh5L184KYj5pqvD55QniyrIHah43M6fLpTptcz+ZE4i1+8RSncUCf9H8OpDlamT7QjoDhwWeb8V
gvXN1gQrqa1ilKs0dhBJJLuxQL/4daKqSWhhrDwSxzWhoPDTQp0QGqryK3I/ZLBNR08K2bMtZvxj
q2+HliSoGISiAUQDt/MqvLn0iq5JWvIknpA23VBhuOxLe+TzH2LO+V7HRzHt2RJuvY4FsXbhfn9B
29VdkPVrE+xv6E0hDLE9p76xe4J8XJl0YxYgpS3yml+7Tm++0kokJTyUy5QHsBVKU73dDY4GOfaR
cdRHzi0hJIbPIRDI2AV6RUMJMa+DDb9wCJPtBUTJLdlkfkglFL4zF0+OGZqx5HHCCT+CrT2aVGgP
C/+6Fq6PkZJ44+8BuLiy+Dfbb0OYFzFng8/Nvlo61zZM2eQD3264YO2jUekFeNVWXm4Z9eIywxl/
JQATfgkaAg8trHYDOjOQxpEnDxr8J6OLXflnQd345Nvql6LuvgfMj1Pe9y4zAuYVHgGpvPJmu/8F
LGa0H501CWt2hAAOF9Mg8jR60PaY8Rb/H+1vJD7G6TJt3x1Jqgdb8lWPutWHHRjIGKoMKlXcYbV2
vsqeR5wsqOv3aE7YndAzSXg1S961LwXCcQGptT+4QRzw9EPBLv+RIH5FamL78a6Llg6uj6QFwD3I
RPpm7AZ5Zl6X33VKib/uenT9ZzzBeEu3X3y5daa/0Z5ncD3811k5Ko26yXAjeXhJDRrjT9dt5Pz3
Qz87MwCE8FOzHaYev8gNkJiQWMoqQa98pw39Y9Zb9RKX2yoqdhxgMUrFQeN5vTgzqvqJJChkvxra
r0C/Tkkl4CLyQbMhiDePpDlc3p1zCMJ3sPOovFWwyjY64AMch3bCsnG8kuBKRGQV+XPf9zoYzV7Q
jhsMLXuedIW4brkkAX7gYpOGsQqu6fCpwWryiyx6YQi2Y1GhHtNddIpTty06yoOR1Vhr/85x06oP
hnDvzC8VXXHt1q130wpWmPU5GrRXN4ZOabKTcCZ3XMgDyrv9MKY3OlvNszBdZn5U9z6nbadwVvFT
XM7WDNiKuiDk/eZgbfFW8uIkLYq//vb6RSLCx7/1UScNsFGMNw7ImkJea6OAEPHKbYXxDFRHZ+9H
mdcUu8wGJkcoRCnrFsG86C3/dzH6YvNi7/LKDqq3bjTKfH0rZ30PL5YxdDomxP8vSnlE1e8VfgC/
jpifir3+/IgVykHM10AJlhHU4vgy8j4qF/cl+30lAitQjbdrKs1nIa6Nlqwt5qpX7a8LD97PNrfj
dN1tegMAC5cCGbtHFZD4rvk41q3QHcR5tZZhi/QIp5LF8XKBxo36zioZZhOiKwydp5KBJikTLa1E
yI3NHcuXAG5wdg/oyFdnI5rNbNBe8gp3nG5Wz7G6ziLB3HAWkCDxa9oBK81/49xGtQp91Kdz19qJ
l3W/s9wJOtMFezoDNPKHBZhK07DbFTDK/lRfhzTmNqQvWovJvwhST90GR/X+igazsNU5Hv8HXyI8
znlQ16v0l2gbU0nm1u4j5M1bY1D1CkHJ7bn3QimsxnZ/xC3OBE6CndCxW4PczHMT4iKmlPkM6JQU
LPu2VfG5cWAgGoDULbjQSwWhoBa3YOwiwLKJsN5rWQYZHjgI3btbdwS9Xy8ZSmlsO+y/1KWC/vVO
Cvi9kgT38q5q4ix1dJXlCMUb5jndEB2cjW6kvN47GBtjAv9OrcG0NLI+0mFvb/JnMDZqPpMEOcX6
6PrcvnvqnjFTUFJnCRMHTqKt+DJrp7kRMF4RPiWO/sBG/J6PJuKaG/62GJAgI9X+gCwjApgNUXd1
EiTTL/yIETrT2DuZeFaShiCKFdrloZuwOpLpZm0y7CbOAMIeHKwQmQDiRjVSWpkgIIpjv5iuFikV
294hufQ+6OtTiA9PrfCQcAVuI7x5Axz6F8JlGhvKkNL2Ma7ABB1m/9kMdEgT6IjCUikyevaUJ5UH
LUxlsI/7K+TX40r4YMyn8E0UF2aVYHPO59Zf+/khhjMbrx36zZEr+x+bJd+KKwXeGe8ZZKeFCqQN
HscQS7rMvtVlXYneNWsZ05DwtpIUBhQK3R622y9zMQHT72EJbeoMXyr2oO/A3bFkipztQsgrTxnD
rBjFouGQEdnHBX7Hb7kbmVTWdW8rIafI6uaTYfMu4kM5/z2SErKP3WQ6LRtXviMYqKJiCEVh0GEh
Xa+RjwdrPXF8OAf4R52Iyg1bg6VuUwhPSlsR5Z1CltKosBqTlx2VxB9ZPrdtg/X1sRgUFQXGeeLw
uhrxSfQItpy7a27p/JBFdMEir2yhOkRNGosaYa0aaoVJ4XCJTtbePqZdfNaah2G/FIW9EAYOewk9
xZQU56uxOV02BQs6lZJgl5dmAAr76Mei4iuZK9d2BJXLTAXeH/h87JmkrL/9NLFoll/KdRug9OlF
zocnCBAgDlqnX96YXeuh4w/pwuGv0+MqVY42I/v7Mhqr2oSUCKwsiQOPVVk1tuC9qJQ54H0jyKX8
4XSWLOanbczPa8Jp9DlxfPK4c2bggbA11NQTY/l6TTOYp6QM49Za+nfFP/7av8yPQo15/JytV6Jb
xyz7tqUSIow/qwVeIHWkSpd++DEll/qI8i0yXXh9GA5AK0lNDUR5YXrYo6JCDPAyIZEEYpIqpm6r
UriagVwftWyHQb/nAyX78HqS0e3nIAiCxTJYQ0M/w2BiiekBP4JgVkb8ucsR/ZiRGkRYAmFrEj+w
edNNlgd75yirRYUUb+1oKfShaQf/q7NNBH8TcXOeBIbYzcRH6XrHM+fZKePME2y3F/tCllD8CAXq
vwGChoFaKVlUkso26vf7hvKGwAaFUAJM2DK6vsbLM52Syo2KDXVYCXGFeBTU3rJ8Pk+09pWB6VC1
ZhYJVeuG8q6R0ASUgAkw7CEwCtOY8z/ihF/TrRC2QRawkwx5GpH6T5TjUIjJM5WdXuXbt0GMpR/Y
AWQjRuuWHnVyvMaZn/2x2Sur9IUR3YuYd3D12Hra3p4gMBRBWxMltNpebvggN+py2cUz3QGKxIl9
tyA0PLgEGCxf7N65PoK7Zh0O5Om/FSDSPGgQ2z4x2GQA11Loc6bttjvyrT1OCD+cyo9DGv2aEK5E
nTmC1YmcF4SP6qMzrrnFysKoWnry8AKj4lXQ2XWKJssO+X9qIzeOPtXzsd+HAsTJxxelCMhGpUPJ
BL5ViToDK8WQNsZY9IU4W90qgnCyG2QHRJYdf5kWa0kZA5B48Y9akhBifXX9sMUVeJ7TcEArpwHU
xUS8hwd75kuHVHoXQbVUnDJjYErZrNYvLpJ7gPcVYtq2a+j6urKfOQ11MDpll//Irnv22ANVj4rU
pgRl/zfkiUbmuaLfjOmV0yDhiaqcvb+o/1yg1LM4IQncNZ8SchGOhcHZeP1eW6lsiLybSHrGsKUx
MW0pmTzJFcSBWfFi1nja6Ck5JLdi95jSuzBITXe2OH6J5Ul7BLKIGMGKDxCCd0j1R03zDcV0ojVD
5j36G7XOHhiTZSyzA2r41GgE+VMWktjHoiU8O+wmeoi3POrxqpFFHGOM0jzWDAWYhaPYIPwyP2J5
9f8d1A6/qQPJuh42QIVHoqg3el8mKCYjqkubEOfN1FZ9dSyK792guOCtZ84S7Qp8jqCcjBdR9R2L
ql4RgskoyqGEGeMhKIrxOcEy5RpNAEB5X4Dcm8cvyynCPp7znHFvwpvM7dgFgluq8QKme35IS0ae
sldx5qEqs8YSvkCq8GTYS/acP/HSo7moGphArzumGyon11ru3z3lLXlrBa74PkTvda0FrIZqvi7V
govzjwDGVVGLCtSeHATzKVn7YDvXLM3nQnhuCb0H4UiZfTlsPl39co/PWXUYX1IwWRfgr8qMCaCc
8Wy5yVQvw7DJ1wS/cHHDuCNOa4TCL+np4D4uD1Ju0AjXeoVvcmNZuOdEy325FqZeXumkuoMLkABX
zcWEaozYckDLZDHKXyWlh5EP37w3sTLVhlCrwJAi2bFN9z2p2NPg+Z0OhI93d2diMQHcra8bPzu+
WSaHZpFu2QTLgQI2lPHZWRsMrFWBs9keAoTYMv0r77rNPJF7JL6zTYomnKI3I08GiJ7QYBpcH4Zu
ogPcQ1a26Fm6Z5mpM5NsOnrtygJcd7IZLiGL6QpZdGwj+GcbYlFF6coUjX7tF9llBsM/+eTudOlo
LbOZBR1a76qSDf5VysXGentAd0+oREUD57foMfts46GuC5Ky/l8CacWeGcHc5tLrkjvCKmZmRb/W
3VS3IGEwOaZr9Fg3OLaBEYls9QdoXezbT4P1A+Ey3W+Bkqbuz/7S1x1nyBTQbb3qFpeHbhHtDONk
jW7fgyfpSawyIUYIMfF+jDz9Qh3CsRe3Muy65heblvByQpWMZ4mDpqXUlDxrHAREDadc9klxz1PV
JZfVN0/AAE/pJDAdlTUZj45rFu2zLY7W31u03MWZ5/CVKohN3FEpjMps0TXnvypPGDGFuM2U4q2R
RaYT5+HqGo7Zp9pSIQkOvsVorptnFsTmYdFZerKuaBjpyQNRG5JXmjR211+s83kvzVx51mPC+4mN
rTXWbrDvnHFjfSJYdvB1xVjQjYd8tmQwzR81N4J6lsdYxB4qerXabWDuswUEHW5AtbJ5ibjsjv4I
Tu78/DUTvmemhlN9NebLk0+VODuzflSrceiRKrw+SdYvZ02df7OyJ7pPqxvsseGniebFZxjXxp2z
Bc0YC3TM5XuHf/N0AT3j4dRrIKoZZDGR2wcJC5ciO5WnXX8sAl14IvElxr4DtM9EzjGfRNo7he/t
4W77zgDXrQw8gId31TsW/WTzX1zV7teXyv4WYNjLa2JFjhdXzCSvGQ2DyEaGnDB/viRTrrifrR1c
9dFxC/CLAx+mtdIm5fD/gb6xTfYvW1PGmVHMnvR1wLeY7/ePS9YiSS6n7diTbEmif00V2TRajwL/
9hZDoA6WUuIn/BiCCgEipuUf886yHxfuT+RbxFhuXp6YgN6ouYUN/c4xVs8xt6CGi4ZN3rbwVMdF
StkAtW1vHVji5mVwmUM6T56AfLv0YJVa70x7I9DSqLOOv8PfhkcNOr8ohZ61LqWlBLv/Co7kLa2n
EYUgeJvNCBSkzMR+luSJe0sxp8v41DuTaRhu9RDdnBAWHwp8Fwlrqr6cmVf4Emue+XPa8CZ8DT6g
8+m9NIaff+cbwpg7CtvyjKK3goF1ZtxgZqAFRaG7plmZt3NopwNSxQN67aynlkwQ3CmhXl1oTGin
OnDut6LgM+GuPv5cIsIxB3DUsRrHTcoUPYPVZBbQeFw64xkD/F2ECNrroUd13/D6J0nWHoTqAo49
vhhli9LENFiWvCs2Cuce9aSr0C1us7xKiv/egzd0+N4okflYNQTOAwLvOPRjxD9ceb+yMsX5KV3Y
QSmyr9h9C+93enWlBUblitF+Ibm7o2xAavLNDWHCyM2E4ajSp37VH8xAlmb3/aJbo9hnb0uUuNPM
0eiWnDHUuByI3BGDbIRKLhYdeLZgzV/Us7NC/hTUc8/TjgCYd5aNWUmixQkRmapILuLonqxBqCxd
POzZdUJJixiW/gfz+f4UHZyilQ9uXtp263lobV+cWHVTiIJJxD2GYWDCVfOUUBH8f48q0Ioz+bx/
Xe+tc/cwlbEv8TM6TASnJuHnsKDFHJois+GYyL5dAq6UcCdE0GyS3gNTkI9jP9FJ0Syl0BlN63Rx
gNsw7gPG3Ox48+/2BG/pMh+z9B2U+a7w7mvYIwIw+0zmXK/NaDxhC1u3YEgzjgjW4Y/K2NOy9b3+
eY3E0kBzCBmk/eerabb0kroWn9sLkqPOGpwwZFoFl3doYOn3jd4rhLk/klfREnsUxps6Fp6lnPtC
2Wm+vwAnZbdgt9yVKvoYKMvirgV6pZgCC7dX4rF6XX1aI2GbKU013iizetoWv4AD92EpyX2Q/Q4O
8KRI+KOoAaI1U77UvFKxDI7l07kjqtHgLAyiN1MiodGkCwfQ5Q3Cjumlqf0gB+FpWq2FdrUSjSeK
Kfwg5teahrJ9tSHiP9gSZRSOu0bU9QRPN8CbThYG8KijjzTJ+94wCaB+2jku2h6+W0QiSxfxF4Zs
oz3Lw8QFhWZRZ/2sglGnHHui/7tysaCPf5wWNEtxW2vgOPjS/QcGHZTVOkbAqlkxKg4bcwxY8b0Y
yDb7qLGRDggBzdQ9J+2keroLFgjshsbqquc6zStgh3JFSOvHUk4EDfKc6SnI/P2yp2/bEjYTlrb5
EfyWPlVAhNvc1sM8bHrwsMP/TJQyE7wOyAAOhMoQ4BiEI6/JB3FdqlpqfUxI/I3HOlcsTPMs7GNz
eJ4FQL1jwgmmOnrh1kq7craAZQfAtIOwHKoeoPOi6skQnqFf0OnPOgHcW7VljOPuXXZHqe53qc1c
JDFofd1NCIWRi6MI4d6rWzVd/iLxgBimdSyKDe00E2yGqvY+uV0AjpbfoCi6YvuJdAJKmkJBf6F1
NJhkiCqDCqqyuqzArCqTDaBoU5dGR2EKx80Y0Qzda7endjOdrOZYgtKB4EY/RgFp1pevjHDeWX4K
nMmSGeJNhNyaumdN7gIugDAFZTvgkjuB/8kGbrxLZhZdWRMdhsmdpRFUpQblIr/+A21V6yBL7Ig3
6SV5M3CYOMe7lAPKub8oRVS6WQ4XcNpfse6sRs+o3YIGjbjEpkAojCdKDIW/47YUp+XzCEnF2oSg
TlNDIi8Bw7IgM54ENNCDI2ZwDdFFpqmNXp9wLywzUbYeenJdTDvzn+FJE46Ignu31j6UmNvdvfgm
flG4pKwQxSwv8nfAuNVT+uPelnEI8LBxyaRFhE8V8ncjHdEZ/Yy1G8D6IpawiiImK2RSmIMNDgsz
SMze9fqfvmtNWnxHI0XYvjJfNEDS3XTu7ySYs/fYmGg/ICwaRwxnYOp1VaaD+2K50bRNbNuRVYAv
cVAdd7/blKOcYN885oaanlQFKsOPvchvj3fvI0P8c/UMDYBw648/kacZVankIcEtB+ekNkTpzdA0
NG5BvMh1jcXD0UG83dqLPpz7eNEYlpy+5O23Vk6UeIFNCM74SZRiuefjDTVLbMNR+pm+PrLwFDs+
gJiEC5lF727nAf3oLVKUE/PlXzwPQj9DjI9b+bxd/JW5XjKKziW7rj6l8qi3tN8/hv0DCrcZiWSM
Qz4UnKI1LoCW0wSG+3u7bBViKQnBVz050t/soIzxqZ1AfS8OfR8UVu0R5BgJGlGbfhXQSBiqxCrs
ZNw/8NkjdZP6HEE8n9O0Da4RrMnSgzBNJnjwKstWyvSt0qoD80hZi5+gIaxFFfHkhOtyajhbTiML
kdO3162SQ7r7pt4Xg2l/zrytKzOYYyOrMHxyTBi1uaD4PBMc7l8ytuYbah7GkG9wkfvTS6ILGCGe
WcdWs56+Z3+vTFCtDJr70wjIWqrUajSVCoMfpVAuBrCDy7jrMJTzjsyExDh82Q4eOz0DYpxV4IC4
Pi3yNtRbJ/OLN5hyOjTQyi0ZztQ/DRsN0hmO6KsrtHvCSxscmAB7odEamFzEPScNW3KaMj7TW+LR
5z5UOFjtEUsnovbHcOG/D6aIpfQwdG34c/u9u3RcjPZjvW98V5wunuV+D55Rfm/zWRCWsu4hPLsl
hCShYaNiOUdEhd1+Zl7MQPo+kADnM/hHaE6APiHv5pt3RdtaQleF+E4UYYwINrFLdthWNmNbyCO6
JrrXPLOqdTIDsD2f4tcitNifP6Gla7PJ4g13IxlRshWUZyuLsr52eddo+YasloA6HWUU6IAEE6ns
zp3CzhmBt7kCu00K+sfpZ3PToPEgaNSKOHqvAo7I0vBtedjsKQ/vq6Fm/jnRg5E6BhL0VJaFI54A
Z59FknEcAik5Mx/Xl/P7lb0MztTBREvP/FzQBUd6TxM/9t+rEuAWtsp/DW8eg6ZxJ77SBKDNoMxT
D6eUYP/QElgWgacxp3Z/DNHZ+f8YN/s5W6H2va7CtTc1kbwZU2nHD0XMPPViJDxhFUzQXEHkzrao
bIQk+wUMfVNfRHKhKCPH+y0JJtWHyFIbmDIuwFQVslBPfinbrgyidVbg5rWX8Z/v9L/Rk7SY78P+
hMg4rTTSew+NZyQP9WLbYsdxwWqk9aZZL/DsQZDED8J2jhXXZAysDsNSJYwlw9C8W40Hg+DGn+3T
bUkWQbV5Quau+JSltYD6+Edhq9GrwsBLti+7ERXCd0enk1pTr007HYdnVMdFoOVS5TVfk/nlyGNf
bpKt9lTDU3+FsOa5j8D1ysVYNJDSVLY+Rj1P7f0uIFYbxYHuSYTS4f+T7wefLaq9oaMI8O6JFNmd
qsbCzZP0Zt50A/l88FhgsEYQrux0q4d7uvywUx1suBdOI+HPmCuB9ptiDlmb1DyXhbchu6aA6BEL
voKJ4J6OmjtGtDO/PZ/7pDCFawrCT/KG/lNqJiaWgN4jSpfB+sxGgdkC6dvSxyp35Qo8l3w5MZn2
SCz+ruAMeGw1zQq/WQRmjMCDtA/VixgvJXvzisw8qYWStqHqJoHS94NfvTqE6dyUOoVjjm5f4Ryo
pANYCzPGCCgnP33WmMJjVAmAe9uzvsoL8q9kQbu6Vn6A/joKwB6XXfW8pP5ZCyk/yk+lZgzepZkh
4dgRzOHToD5p0TSg3yQ2XAYudxfsgdnaFJaUV0Tvf6jlzg3rFDfNfvf4LgBzuniTuc38hiHLNluz
YcsQkISLJIADJSOxNn1dXT9BlCINrnFGc5X5Z6/QAujHjt7KCTOw0pXuXcOU82B4EKNoLCgBLqOt
dpBxf9BKlVK3qqbcL5w1rDqNhZqhm+M0j+1XeAqtYQcz5ozQdA0EENazhoPZgmqBgdbVnGuMDFCa
MUudu/gw4HVUCBDQdwLokUovJ00xZsM6jnaWFo3yh43e/dRVx5Bqi0iz0TQO6TymMESXBPg9abOe
2dcYokDHinBgibHyMy7Wj8/NkfpydAKk/CLHILoEMMUdkwPdAcL/dW12Ul90UOHkbo5mq/QxKpqg
rPqFkcICiFke1BscWD9T/7faz5gzZrDc9Z7HnE5OoiTyzF2t11eSlm8uxF0MVUdbtl5nwPYyTMsQ
KOojmRG0BwkUDSFWiXdrXCr/9PUZZg1U5vfn8HmLLjwfwvKPrYD9NdGjpQe98SPyQUzqkJYF62LJ
vkMJs0fY7tFvcc+NYFHhsvODcmIp3mECbEsoyUpbxyQxDUDN9YReYJlex/uQ1liGH5oh3fsujShI
Lpl565NzyQy70d0cCMdY6nLTEszpazmAUGYktuuv24JfuX6cyLGiP0MRWwMJvxbfTW66RxQQLgio
WwPF+7exlfh5trUvlmzUCwe0Lw+kYfE9YSNp8sH53bQ+Gk5NLIYS38rxOctrEP4k1ncsu53fZb4c
Rv389MrttUbVyvNmLjc2SeQgASJEbvVEa8ATkzm/VGiShBfk7i8DYjFGulbfzp4yBPlD0+z5CDgI
RbVflWjF3VR4JfHrJHwHF8sQVnTm9tGEk/R+b3sIz9NUjvtW3Umkjknu/ACiE/4eWaoO8UQcUGBw
D6XvG0krjRX3NPJ74j68vR1BUy8/i9Xp9Lk/9K9o+PTzYjUFFgicetfnwSvZOgi8U2ch3594IF39
EDN6N4m+d8Z9TFwI5Z0lsZqBddrrMb8skwxbslZGBwCmghTfk7uTu4li0pB+/WKbpuiKPb457eZG
jxybDfjuqCzCnmTw7NRJHtbPbPfmHzNUMHUYXUG+i1DMjJ7N5deu9X3lqJNzseVTqvV4cEE1DppH
z+KavxvFZQ4lgcF+ewC3f1uEFCD8KCNSxKf1tPFEgHzIsReKFdzdzTlFayjfG5qc/Swg3rjJsjgr
H03M4MXc9+CjgvsW4no5U6pRrnUhKqIpb7Xhv8ODTWykvHvk1RunY+cHebA38zugjFIeR4gxVV7j
1RhO/i+E1Ycb+9tu4gXdjiXq/MrumElTnGXZ0h/zXoxDiEVoOa6h1I+CxL2zXFCmHWCeQTqBqT8U
k4D0PdaqXaiPWjS8aWuXwjOnj+B3pyXL8LptRsWNc5tFTjHU+WX4KIhQMgC0xIUNlJE3PddpltjA
DGWNWjUeHuI8UM2acrm7HneWszDJt0w8Jnzz6wzwyOJVzRiY8qvbltoBhXGdR2EIHTVKSzITv/bu
6XWWfCcixM0xif5OWP8X7CqDIfpIbfIQDRtwaKkHV+kaSCbH55OE/M2rAKZ97IxbZM5BbQ0WyIQq
/BKEHdJNsvDAVtHl9ety4cTihQ94n6DK8eJX/6iIpWmFPOGS0tb1SS2lNkMacWDET/Rz/5IPWqYa
a4y5TcGf3Lv2a9/2Yi+JpKKZ8caZIhwALUUTAeAS5If6WLSmuR4qR9H2ov2XbcuLQdDB1yWPfDGt
hgtKrr6Ge8KdlOKP2c6+D729BKQ4d27h3vHUQekiR1ReS+YH+2G/zJEBg1krgL9cvzikNsoIdNLk
1FPaiiZ8WMKgsENHfWYzQ47ATUck5YOZgGTgfL3u9+aZWBIBNo2HsS/BOAFFAb0U1SFM5Ah2EMPY
6FOle3cjnAmGXE8j+o/uqTcnjxhYeGczTYrJGXUYqfUD24qTzqUnQIsB1MMzQqH0lkGn5w9pFJlt
lPhB9v4Aho6Kt3vdgJsz5rVffpEBfnWk8vCXyKVmhAA0xNViZkpluj1cvHCv4CRoSHoP6HUl9VeG
EEw5Zr3PoLPyA0Ku9kOUDJDphW1U2a9IcEAjuDwpAj3dCghB0uEVq3/+TcgSiOIC1qe8dAWU51Om
G3hqkImzGTxyjeFKXnjfHMy3W5NUBgYvNWAU/n03wf6hcNeDBabVRrXTuc+sayTsecbcrSR+oM2S
ak+N9/ufjAdnDHD5+FVgtmTFJFAlZC895Ze7ILDE6mxP4Buvf+c367uiGPNWYIy2Lck7S5VYigHp
fFI7OgyUBS0CAxlI1414K1fwAjqECGhHnl1G54CMV7xOq4dMNVxH2O6LUMiJibylYPEzotqb1fJ0
MadqZ3Om34oh9PyRHAzS60QAVhAW+i32gDMgLmo0opIj34AxtOqIUaF39BT4hTGx4mLr4OYisKPj
SzFsFzWlnF5jWtR8zfxLaKavT41rqqbGlKy0/wKOYA9K3MJBs3KXJQGc1EGu2mfyXuwTYpgd7pLo
2bzuaxSFcO66/PFi4eip35HpE9lAg3N2yqQmUE+mRxWJWJxbebMlle6j35D12fkn7lGSlViqHcYa
DhCAAHvc1T7wfl1LzfJgZPB5QPOQme/vMo06OO1F6IXj/0wbKli4FOSx2eNjIMK5laoOE/9I8ORS
+q1ZimHBFhtj+Eeb2IAjr9QgKtUjqsEivVo5ZW0amARTmMUQfqoImYncGYX3vzRtbgrvKodxPYUt
R5OaAgBYeIzkP1tb3JDKlC2Busx8Mth9XhLltF8OjIg8a7dfYKxr6exYRzAPXl8TueNDUhbGMqGh
f3oBJHHFpjCP5LooWBu7Q/qcF6zNRV8/y9M1pT22xspy/Bvgh7DYHpTq0x1az/RdaXROVOZZHA76
ilyWbXnmgvDNRmkd0JeCVFyVnxDy696xcSTg0MAmBpSw2qWv9UtCcBpK7aW8EwrqW9iIRYXOSfCi
bsL93jOTur11vGlQJyVEb+LHje4TcrUf8mt0/2vo4k72xFXG/bTMbEzSLiOzFB7dGKcTyxno8S3d
Kxust/+uYaEXWp1AHJH0RyQONmQKt7NRyJtgesJuEVtCri50yfBtx34H53d0Y8Dg8mb8iq8XWzHJ
0PI4tTXrB2Rtj36FPc/XxuPU25j7kEJhmimHL/MtyawJ0DcQJ3I7YhIwJvvEvCegE7cEFw+/4gXR
1YmJ/cbV1jKc5txSysFUVdPgtXoIPMYXzVWS0kcRLpKyXpvLtnKaYK+UKEiubmRKfcIMzUnB0V9t
4l31jn9XSYwOOVpUI82bPmnR8kbz1U2jNYnpOcu0HN4cc13sSY3WVnFsN3EGl5/CIAD0nDWpyzZX
9CQbmW5FU3hWtl3AuJohNj9TNPsxgwhm9SGyzuW9QCVvnDQefPv1vquyq0GGcc/uWDmdGR1OZPCz
F0b4Pim16Ji/ie+QonCHit8kpjo5wHpLUM8HC3FbR7v/OUgFpo7O9kXbn53TF5blKTqSH5XniYoA
56ToKwsM77WkPGBwSbfE3ClkfYyfNbm0MuZ2yIWvmYEsFlvYEt2F0dhEmqErv9+nWvF25uF+zzVb
YLKCM1TE4qNhyYN9jLSBc1VMkfjrjnUe5VSHM0rJkdaW0PNYpDh+mBF+WWU+G0V+XklXqx0PBuQf
rMjOiXtWVQniBIGaSKILFCODcUOfyH9t5TnCXtRaGe2kWxhK1uhfj66w/J2/qbWRDuki6WjBvXIA
wYbHsH71kIZuHtqoT6sKzo09swLgpdD/Ej94WaOS97xp5MK4D5k3+bAlKyZzoQ8Cfvt1EJVnDKZ4
qeSUTBSXB2xlJoc8vpRdHlQqvCu4AZtuehc8I2BSLDdJPqw8Pl3iWmhugZhnf6SC1+m/4LsYfzfc
5vox+lWXqoA6fqD7f0RhGpbIpny2W/Q+CQEI7LIQpP4eLPlan+MpHO0nd+HaljqoTNn6MCGmADHf
TttTFCPMsif+VPlThMZGSnTZzAK6lu9UXLArsB+c7KfqMmdg8mds3ZiMJ6a6YWmOEh9nDbcadks0
pH60ZaXgM+EIDzVC1lQpvR4sgbvpqkxMmWlLASodspNA6EY/ufwj1B5F8wVReJPb2aPDqacxxShg
hEJaQCKmFwtD2s7wmvpn6E+zV6ySi/rl7UycsBCj5m7QRgvhkmXZbawtjChEGjpv+Nwl1slh/kM2
3kQsaaRWWPtwQT0UOjq+8eVCWFxo5tXwXeExhMR7vunZRM4xv3rmwA9Lgnjwhb4c3MZpN0kcbgpD
fkO5z9IHFKXyCH92qZm50lX0h8qsg0kwyoFtLdMQX5KNrlFVn2cZpTHhcDuZ98NZ5TkGTN4z1GhS
+wcL8KOfKG7n1nk78GfvWXpc1a8GG7s9j/xu1ud1RtmdhlpVIrExc0OpbeK1ZnGGBJnGLnaK4VkE
t1FvALWRyU+eEksYDcBU+IhGIIzDLYEH2o0Da9QzGRz7imZ2c+PQBqwxYLlw2z1tL/efo7S5b7uH
DtFBjGblAmgol0bzmCB7nuzua00MtISf0q3EI/MV+Qo9Z7LkIzsAkjSlagUKtDc1D04qun8miVLt
HnDdq9vQzXrO9rDtsn9adOfIxiHbqDTgY0QiqYXCnfVuiMQIY8n26N6qoICJdqvUfqqNnwOY8vby
Io8wZDuOPbFb2q3M8joY/UwpHq20Prndr/jmO8WY6YW5tHEFfMt/hVxaiRIjDoPwHkuLhb7IfKbr
xzQfvz/y3fQxHc30K6Z3EGjblU+vfE3dziK/2eFnn86pc1OrHWV2DoWYWs4nxcSUt5/Z6wSeAJsy
HU2iJ/s6r+tiZWRX3Mqei16hz2V51Cc88s5FYliXYXtnuREb+bx/0IxflU1v/IclfdRGD2OhV4GJ
5H6XNngNlFZGZO59jbZS8sfTr87NiavI2qguBioP9jUFAM9Ed7AqeST3kMprwQoWOMSCec4cKLvd
Xz94YF4Lb9MedjlK/FDRuLmctEyJgPIkGrD/u5AgWISfL7ZDyF2IpDoNIbwsRq27eJu2PCI01zJE
DVlPJGUjTH1/daZqa18h9y+FZwF1raugFCsBtHRyP9Oku+0e9r/DbmZNfLoS9MW/X1/pJ3G7pXSs
lGkLJfJqXXP3KL9ixCBI9B41HV1BKb7w1EBFD95bxMuLu9zWjNcw6HiQTBrFMIQOXHW6Dw8joTa2
JMaHE0bQPWEIPdZ/9kB9M5+u1Ocy0pgWfWHrqlB9GiHwPamyB+73hZljxNdAuzYDyalfurX/s0SY
LwrmSK5ORhrOm+q+5y0pN3Ev16r3lnreiyHRR9IKJKaYRUQXixUtRHAifRHAIHhYH8BcbRieIxQA
PYxSzV/lvxzWyTvD/zQUD3yO/mN7Bx22Dgi7XvD1ByJ31cmlxfi0LKwTHzbTcUsTU2UHAni5lsBf
FoGM0i4gJo23+cWpTI5T7uu6IQiiFz8+vuPdu0MiUihzCTtzEKQiCEyoUfDfzaiuFtgYK8G0YZuH
ps6k/W+8FavfpYDwcyPhOQ9aTG/2G5VRrjAFut0NBRyiatt9R51R3wbHZK3fhUB/E6u5O5Y/Odi4
PPdSAW3fW/feItJS8F966OhsNock4TziQy/wsXAXBsDpK7xSZU+kb0iaObgVsIid50FKR6LotGFQ
G3Gbgd0b0Z8aWQSY00Loh8LHQpbkSCtjNEIVeyc6CNDEuLiwnzUFsTaksEmUVNg90D2zT06GRqHs
UfQFW68tloYgCM1pK4Zt+hU0IYiS1XHPivc/GAGzyvQr6FEqTTcrBSV2BjP3yzDPtO9vtRrmUhLK
0dXHIouiOxTDHLdpIAWbf9QDmuHwExqfodkS5ca/LMe9nFLL+pRHs/wgHHVVxwYbDW/b9Cb1DjA0
mAFCQDLKqCbBRF3Fbj0WRiJuAaiH45vreoJGsum7lUPWrck2fq2rzX+pxy6t0r8uxeawdII4FD/a
ZjOLjKNlnOWvtelJy63AKN1r3FGA+l5brCog5HZkngMdwyssy7+r7o6TDg+ijOesUTiylAHrS0ls
mQ1Hz+hemrZ4PLwRJNmjGxNizf5Mq15/Z5J7FLSoWmjZbmTnEXcTWn9X/l5m7FDDH2lhWTcbR3rk
yAEkapec6926/TfWyniBrH94yjNddPiSAcvlc+uzM1Bcs9Km5cOeJZOPPRlFkNx4lFDhhdlpc+Kr
V5iEsFTdZfB27QNbeXgfzhUMZXxej68BNwyiErQmNTLMSVwvlwEYGLRZKFgtMfBELhy68IqsCuvu
lguUTOMGzmNG8LJ0bRPCIVvUMCG2ZhqAH1hngOqA+Prdd0LOkD/Z7QwMoBFmo4htIMyw7PlRHJBi
kihN9dVdk0+M8u6+uDW13iozVFSINykxD6B1gyCl5DeQbTCrxeUlB+9FF5KGYz7zwq7fWi1hU3/t
Yu3cFDMFnjj6cWWeoe5l2Nm8IgBcsnIGUXyNjmpfuH6ts+5GqI2vqvLonXFhLDvYQBkC5UWun4K2
V2D3KFhKH+ufHhmssrloyi1QspAPR05Zcb6XRvWHyRJWVUObXAHKi+Z+kwFV8vfGBA9u87JlW/xh
1JyRAyZSukxaJUr8MqXt5Q2SQZd4lEfZI7VuQJ3/Xli3SaHqIM1llCRyrly6z4tJMQBXwee5Nqx+
m+QSFjGWZYNvFc1qIrIfY7CzE05kk9Y+Fa17dlTr3QSpzPRttzDL+P1T4tATJu0o836jqKh9bkUQ
uyerhzl/i6rMOifmx2C59EBb8DpRzkbpU3EAmaETqANyKJVtneqdeLvHKYZHqW0g5eO1TbX+pxB3
p2281oFaWWBhBsPCkizEsCVVmHVUHMQrANHLfyqTkV+7N/ZAwR8alLNFV8VVSQl44hwL89ES2zlt
UXNlPXTEtNhY4ygRpSUkaOZdGPPjc4Rh9BRShe3qpT4nZA3i+h4eWda3laNRIU6eLtf5Tlqlfarm
cVgmzCdIHE3d2X9ADSYEFPY+q8yPMfwYY8cXvizDQS/YIYX+VlshcA3ZgMxwDaRuePHpMjY2e3FO
EhBfZF8qhX3R4SWNoIts0w8xRlZxSGl4UDbXjwhgy1FfXypK3/ZbrfVfuUeArcJ34+3j2fjxXD5S
VKz7SW/UmIvVohAfQMFwh6d2HD/GCz5P656w/w2MT+h6yMRXpmzdLiOKSuWVXlas0qPecx2RG6x5
RuP2XJHLtK6wuDE+GJN2Z8dRrf0L0UJ2ZHFpTTKvyELsUuHzOTXD3PcoavrkhfuaMOt6bvz2MKCO
YT9iJcA3TmnJB8iNk22jcxR7Ha11zyQDbTYR9WnCqSS6Oar5HJDeeDAPSSeE1RyKCqceP+AktrA4
isbS5q2rZxaMgzXsopxS0i8Xh87ZLwkLd/UfQ8JDnutN0Q/ikVcaTRt4wIwFLKEclW1ybl72nMOP
57aNZbEOrZrX+klVrcsaMvypHpECWWaQqtazv5Dx4QJh4hBPub7Rz5Kzd/y6YKq5E8PdwbkV6p81
wdQ+4mtSXNysvZvlc+elFxmhaCwYQjjKyZ4ka10m1ZTk5JcP8gBpnWUXEUCbU2qvN0ALGQkGrvfE
5jx3skueETglcBtB1EY4b6skMI8wOGJuHZq9aFG8u3Ity/lvCShjOFFFrzz0wB0t5NXX6VfgWLEp
sd5qZwVOPFLULI5b9PX19uG1dTmlLL8WJ1wPNrCf9YoV0tfei0ANtdOg1tTepAtSV+qHIl4nNutA
CQ70FubW8f5Dv1942YBeLyDGh9dRoQs5wOfb5udmUn2zUwpSQeSAigKCpNgBT9fx6EvGDOJ1rtP4
BnXwWn1EOKgBaVOtvtuYgGvwg4wdZL4rFD3ZS+87nq0Xig3Zu7IjVkHgRF4J32FLLVc3Jf4nKb7m
xTmLv5QXqJijGVJunIxyGVjamur4VkqO7DRjZl694rhkQA/zKRLSx2h2qPDDRE+6HM7hbJ59Lz6F
8EN2D+cHgwXG9vJNB2uiKJLEikIFbbAVMpyd3vEey92kWNRrz6hACKwvW5+A0O9d8njOobHHwj36
Wm62WawdmsFT6uy6afx5gurWfovYQZskNYAtOAQiqgvO5uSJWX22ot+wLZWvlRraEoPRw1R4rAmS
orHVrBpUeas7nT9qlmTrQsoTo+LV/vfzoKRMCtypw27lkDV400XgNhtZKsnb+EVpAZAU4KN5/obd
pAreeCh35qugtIP2Kx/6bx1s4mWGiSUViGDpv60o/rWPQV5XEquGWLX32xpqXWUOrJ7YCldYcuTX
wAgHi1g+4x/bWtG97fIzDOvI4FNS5nXduaVg/YVmqUFd0MQJM8R/8ntxOtiqMgtw3Bw82dI/KDdg
b+7aGfN1DE1q5ooPqDTdPiPYQYb07JiyujuF6TXAkct6j89XV0YyfWP+4scMZMFSCsKwtjoik9ri
0GvCTOX4j1082yda4gSodfdEulM1V2aZcMdFt0hKL19+QLtSKctT2xjPbqSDQRlcA+Gto1xo4tAv
r7XRnWr79zMrQBb2iPFvXN0lpSXz/ptFnyYnBK+i4PtRhIPtuN2Fb4QkvHT5b8sLM3ScjcDyhltI
ZrrbrJHTemhQXLpSdp5f7JjI5hARPdTqviIrAi7VPxWMYUx6eZ0FlhlqgtsIaql8OtljMP3VAzdq
kuti6nKa3lMcXVrery7iFWBGteJ/KEaPm0cuHOFCv7PiwMgF7vfT3Reo+2JS+cQ44sE3K8vMeE94
EyGzJ9NDtMwQ2d/Po6wzq7PftWdqGKbfrv+UgKJk0bChRY7BMjbSWH9LxH5DjZotuG2K97EW8oxk
yJFk/H443YVvTyt7nYdC2M4mysfINUu1BWnRUOBkFdZVKuxzHejV+LLNwhdg9ew0DBRd3sAackdf
8B860lr9Db9/j10XNJt0y4xc1Z+y2HUVcPrlljqsCGNx6EUYB2Qf25+6IPhhp3yI12MRJqI5b45Q
a5XKhAGTE61CkMk4EaVmJ8bEAPjhwUFeNO9o6wwLF17zL3WO+ZXWRh0wH37I3khnmg1vd1QQNers
NhqxDSDd8Q/u+hwXo1QlTvlhZa//rsVCgfmQd+/47KGM4/DCL34AMDEF47Gjx/royuoyp+4M3pPR
mTmvz5FivAUsM5VssRFR/fSOthZDV9cnJPrQlMY+nRdn11vl7UcKw3FFJp/niJu08Wtdu0sguKb/
luidrD9yWvA+k5rIzzTlScjbsSYmER3tU8ddUWpOk2ccpxi0Jhbd3KmKPNrw/xOXDVergWdRDtm+
l3j8Eqyi12LobajYd4wxsgaeMKTv7zPTiTNeHX1RFIbuSlR4YIuw/AD2WROvJcBAPquC5iNS+xO/
DAKUi9qqHiygjB14H8obyASx7NV4Z1NVqqnt/ihazIOgPjLitVh5aAxp8DIWTdjmnJ71O550doL/
+pybc6WZEYDgDtlxiORhMFcuyFnNry4BY7Bro6Cdhqndggnzmtg7eampAGtrz43TCM1u0wG8l7Bo
Hxe9yd6MXhv3lidFjXVtEpZjnN0vgw4xXEewE1uUYyrry9ZlSdXAWqWlslDb5NpcHXwpt7ao6GJ1
eDZZUVp5lRLAGeNSDg34XyvG7SLjp+miPrWQCgpGRgTE9bXZSKZOe5Ku8nAMmczP5RgsPsYCuKTT
GQfa3X1may9JzHY5ZBHACE5HnVcK0t/ZQvy+/rYVqQlIvPdX+X8O6jGzAjLM5/rGEpS5Bv6lEILF
D0QODmPVGphj55ZY/cgLcvs90KYBeiDKXuRvkx1lixy0zyCARvSr3k71mKb7EW8ju5lf49PSNPca
utfGf6+3WprpXVwIDhh5m39dU5ur5+JdOXMZsPjyk5adZ5gE9lU9B5V2rponqHUx4tYaLJzS1HAj
Mpf7wVXiXf9sryDxBzJbWUW1oWSeCJB7zL1RujcdQ8ydil+a/s2iT/Puo6AUQq9gYPwhN3KdIydd
pUpTV+N08sHymeSh8DhyKzRWWiNBPN8JvVsU6K1H0Excs86wDDTXt0i6WvzB7aahC7Tjjah+haN0
XEKjHKQEjcELwun0U+UWVX+H+eYxux2dnjbrfVqUCTpL7r1hDMO0RmSQMSiRxhGYROrXdrvsZoLH
7kMjh2eINK7uxoqOFWjmhGGXi+AVekMKJNNNucCbGcdqvgiecNJu9Opt31lmZsnxUJK8f2apAMsK
Biu4SfrcvoKEmJCR1Nh8VG/k3j8zi/sE7o+bkMRU4qzylFmJq1jDeNXFxNK/OTmQcMSs56evUFAC
lJwpHDLiZQT+hFmyRpCJK+YnFXnAHoh2OEE+1eY1De+QMCqM3yG9ZmNi0Kp/wcv5wblN6JfJPCwD
D2WMmUx/KH2JWviMfOCXov+RU8JF6a+Cs2Oonj4zm1pvNanIJNPq5A3R1/4sMqpsWaA3kvqZ8F04
zKisGLW2kC8om7QOS5/tsFVtZ579r1nZCoIUs2Sp2QrRwrmxnsLaJb4KfrxMg5sIfeoN0RC5T9Tv
gN/J9+CtDfUKQKoQegT+Ts3raFIh+noLrrmFpHAAAeSCcZZkQJ9RkMUy/M0++tf55Wmu1NR4rGDX
bIphvu98gDaZi7y6L3J1w/rt6Lw+F+dOR2K1+Ua0rjKH/yVo8gy6Ie31Tp1ndFWa8OW3sZyDxIFR
GgV/Ax3bKZgTvSUw3FqObnTFJwWWvIfr93mOaH7MJm/Q1eSaRjzyAsQHHNgBAxKjAv2iZA0KuqDw
JDLME/qGYh0zygZ6iVvON7ySKakJ77ghuISbvgAe3ivg0OeU1ZimWAZeLB2vIb8HegSmah6ND61e
j+o3R35YMwJeJ6IPBALiL4MNcaiLL6MzZfB/lN4QjMrovaFGrXhBmartdPKDKfR5URQFd6IbBua2
crSli6HFx34GTOj4Clj3ejj/h00jFelXpT6KlYg/hXxQn2Xk0GdbUwBLy8mzfSah8jbdxe98V+tH
7IEF/h9GdHAAUhTyKPZMKt9xW8CukrVLn4PwK/YKhQ0hxCChgdoe1/eMmOALsydJlmuqxW0xrniy
d3NL7ohVJVJMCJPhA61kyHTKPQMu0R2XNyUwuoybh4hNnYhWVEz8zgZEo9045t4tRU8qG8S69o1Y
vHHdrjN8n2Btigdjg92MiJkXe+ExbirrEkfw2A45hxGMuw+P+tRhemyLbMJ48bT90zKL4YoT8MvW
EKf463bmEXlf776cxr2Ny5mx/3BQZt8XC5rv2VB/zGjb+dMMOpnXwH7kq1jpgYXUtJvPI7//efxC
forVJ7bDAsJ7S8XSaBZu+BLPTHIIuW4IW6QY1nSLFccB0bnwPt3/oqIpotHXIYSAY/jepaseJjnq
Zg0GTRMLcYJBstGQ9LJCElQ58vG5xYSmJL2f4nVe0On7oUfDs2YuNfCSihciyKRZxjdINTghMzYV
N/gpCsNpe2vhjjOzE2wlGvVvNfgnbxVtNKmOb3033kMqGwQdJJDlQp3UN55yTs7kpZIJDoay2hPF
84l1fVDwV97TgCyRx8js+fsZLi6S2yEVmW71ot+ZrsL/HvLWqEAHtwTZQ8zGAZzf3kg09XNNYmTA
uxVA92Oy5y4tarLkFu27GucXdMXn1XvZP0HKjHOKAc2Pfa9sjPSUDY+kVSWf0JYO4CA2tEKYmfbI
jBH6kDqJZFWBz/2bfKN49Rf9XCBVLIWYHho+VyeR3z/aMGTaY4sb9TaXy9KkGKMsTrfIWBBSqf6J
1gwOMbA4zeDL7/Kbl2FT8kf84Ne+m17YQs1zYOCzhLTIAailRIrhuoddkr09zzF4fPDJKngtNdn/
ANeII7Je195GoCWpwCa87kB+FVbxoLMjEGSOZmanqGLOF7+U/whzqt4ifkY8IzUbWPn+UwS89ryP
7UVi0UHAMY0U/rEd9hWNYLgSZIBdikWwiA8h1YM3QcOMw6GsZ1TssiU0MLwX03SZnQjA3UOigN44
eoXfzmVRVfkQdqOJgTp8lIzIwx0NA2zjA8w2FlcGEDpjjBVCI/C3H2M+MZu4XmszHFKl9P7qauwS
IDyhlXRGzQIat6Op6gG+R/thoXk6siUf7358jo0tK2cGT5U6DWNR7X/72WmSquOSAnxccppgdtje
ZZ1oM7LIGCDaVXGr2Jpd9/SLr6YWxDjEiG+pD/a8sTRhh2lWX3o/WcFckx/9bpjtVcu97jbCSN20
C0gOmheOuqfrdiK8szfR5OUc/u5b6st54U1hGe3Uw3Ei933mJFSO1G5e30/fJRJezF0tSTBXM3Iu
8xFV0JifR2unkl7YpWDctcyg3TdOUW+26UCrngT400QO+Zoi/563Llj8r4lQoY5I8e3D6PEiUXkO
npo53XPJ0vNhEWuxbEQDfmUbbr//U5M688h+UWGTW9zfQgt4qIfeRVERsUfuwlmUwfiOYdHVGtOf
CQx6OAu+0NXDS79W7wbbErJzzQmNyCJtwdHc6leBD6Z2MPqbbLi/PBm0uPx8OvsaXUX2nt37mxbX
Mv6P7JIQsCdKgPV9tHx5Jmmpzj+u7mjqER6du8QzZiMZOiG3TWBdcueNlZXSYATke+oLDBOiVZ8B
3EFTuiszc+SeSY+d3qfjnEnzzz9fd3Pzsal+oeiJfFTB2IAuqYNiWVp/5v/+x5WSzweoV6n94CBz
mSTuJog6mZcsr3U7YAD3HG594oHFkP6fZIdXyt/EyUJQEjr2sfQsi+FrAmyjh7Eb8uQT5QpZyS2C
6unR+89r8rGeEQkChSz2fP7j47OY3t0ehDGWcHIN5bymezlWiBXl1q3l9szE6tfP6uQ7z7b7cO3R
fgXL5c29VLN6RT/fi5PmMWxY8DlfYF16966Bn6U9aWxV/27p6kB20WAU+ri5kTDhPZRkjxupbeMa
JO0rHCsTJG703Q9jEwaJX2j4CMGc/ZyLdRAY1MJNfj2oIzJE1EVCAuKb5d+xZ4XE5GKHr0X3Noh3
GoghPz82pwbvgN9Ie/MqHSwa40kDI+iohkJ8lg7bWKAyBLeuUJpcN874KBraOTd6ttpybOsu5Lxf
G6uHRDA3sLm4344YomINyWEq98TJzgz7EAEN5TaMaIAijruWqdFospkykDGD5tgXIh6apDQQbYZF
eErVETg3yQGCsnt+d99bLc0CHu0HpJ/hHwZOrILqsxPmetsx+uukBii2d828CupyH9SOqERWurEz
vPQKys0t8D0UcfNXNfO3RFqoHPcRNMVlo6k4m75Ojegp6XyCymBWm8gSCJLltzvgO8RBkA9BNmvG
yGKo06jJpVRe2cqJi1rs+Rd/aAtyD0M6b0p+PdmBqDgNrWTbU2/DiZV4IeWzvldBpERygjKd5i1E
zAzhpF48qOqCS5hrvHPJGXC21B8r7zMU6SJXPfElLOEghWds9qSNDdDbKooWbYJHiqbP+iCdjP5E
FRgTG3AWPr9nrxf9riuCBSZfta3MUfNTfbZnXlhguElXklzKTO0f59B1n2mS5Y9KLc7fV6JJ4gKv
5CmmQv68oyQML5YD+D43sWGoTmcQY/jmvZv0pudpzL111+mieyIF9MkVg75uLmtW37WAC+8CJG9B
ESpgwQzc8+5n5aeOmJ2lfa2EJyv9Y8ByR0IWI3nEajRFfCi77EeCp6UFQ1YvPlQonq1stuCLHnqY
Eaxm67RIl1SdIa0kG8kDz6K20tWZmO8B+2aTddArGNPkn+W+HjKRr1wpIGtrIwbZ3t2CUvkPOeGq
AG2Bry4uZIIAHXL+Ee3AJoHf+dZYcmRMnj/RL/B4g7JM1aWc7DZuVZu9+86o9xWbs4oncKdotMs0
ejpsaXKTKYCIoi1pJMIcMWnXbhm2s79/fK5hDFpVFVAK6z8zU6K2mI01mPQWtWkyiXjKfFQu2yj3
lgYferCPZNGH2XJBWxS0AvbqiL4kCYicbkHvP0MR6hyiEJLo/SfTOkj544ZiVfiDCNMTsRxJHJ7A
6luXHxCz0Bhz2iDrt0oBBmuKFhbf1uo6ubQxFNz+XKGLF+V2nTgqycMHiLQl+6P8wTZC5s8eKGGj
6ffp6eBp3cwNm8tc6CdAZB328rpku/ImcI7pSGFD1Io7djDRVWHmYrThftlUMRbePzicfZCebpKH
J8IiO9wfTKR7T/XihryFd1lAfkKHDDN7gLbgNlxu5aPLjG+/XxCwgG4e4m8m3b3Kphtbi6lYbAJX
C1nI1VhwVPLwo5yLZLtjRsQyPSujc6DoZ132c0HwFQF/BgbyH2SSaRVvpYr2Kr4HMnt4qA1P+geL
nVs4HyqJ046AlRQ1KFr/mPW1QA3IG68VlLgSWu1hUiBJ8qoMxXgkPp3W2L94HH+yT7B0eWsNoZpC
cFO15O2wCBFjpizMScYCtJiY3/caBJx/KkHmOgW7wmovq3ba51/XaGEZLhLOrwoGaudblMTgp1HV
eHm3l+Ke7uohUzUkuk0xNXSdj0zNMnjfleVab5LnTc/gX7QXNFynKu1yST1FQzVeCMUlFqaiSbc2
H355CF+vPrGVa4NsH61LeLfk/2/0y36HfmEX5IAoUNP6XarCxuuO59I08uL/BSRNLLJrYSzPHgTz
AJ8jQvorFTjXHYZ2bLx6Tp7o3AfC5UcSrOpSG5uthRWgatfu8QaXtiysGhCZPu6CSognHna9DETQ
aX1N7v8Wh9qKVZgPty5wdrSCgtO7NJeuShavofwaurcly0hJDFsuz80+64WU45o6gQbAFcp1N+lS
mCFt4MxMu8UleSUyvNy/bMswOR79m7+dR/HDjjCs5pkYpW6drSpqdg4qMO/FnlRdC52KpK1mGy2i
Uy8aZzviO+yz8q712igcNKo4jC4JMCLHsTerrQrTvOdilA2UP1WCRIAZhwx6eDd93U1pT2btvxED
rWwRUionON/d7P2EQvEScYZ5mcMua404Awf1YuiYMkhM7a3KYSJ8m58YUYXVvOAwe8F1JjmOBqUY
e3daF50H+5R7Xf/d+4WuQ+OKtYaN92FNb7UdCqTXfE0FMOt/y9+5PafQdzptfUBK4odOxWKBXPmX
CSaZsVKtuadHkALNJCkLhnj8apr66OT4gdU1rl5bbIu7LgR+hzqFSGvSVV7abvK9sTN5fR7IsVWk
BBqOU4ctxc9NFdsSWDha/Q6UfsTMXYcInzq+OwSGw4vWd1vwSBqjcRqnzBMH99v9veuGesO6J3wz
VZj9+ffABiJ2TJgyeCfaL1HPXF0gtJ+lE/8oL9uTt3Cm9FwF7ZaRUABPBOEBAAUFTTOvvqTr7vQ7
EzqlKuHg0WRG1LBbEf+i/rJf5nIGcHgU9f6VpofkqLRMqvmONn1+ayOORa7aInKDq+TkFp+LFkp2
Q2WwkPC7QHf/dXy5qFAJ1X4BJGDrZZ+sX7XQTAfqfUIwM/QwimKJKKcoSObSFCJOcnP5SmhrkH7o
DggYzOqTP/p1bCOVQt3D7Nrd8WndLl8He+JpRPlt7Gv0F4CVz9/n+ThMfBCx1N5uZz9a10J5Q82O
TkfzlorD3IAyqScHb6bolvbnLML2oC1gbiiVy+W2t8QzsPq8KwZJnhN5bRagwlmTIRKDvcB4xuxR
Y/c0SYthKZ0iB4w60EQBvwcC4hz6T+NSl+nBAvk1yb8iJkPrRiwH+1eY9+GOGgNFnqgt5uADrbOR
nrw+oZjKU9KVFQwxC6U23EIP5M/qgfgUtrb7Q+lzYOkIsK2oTsdSvtiNy5Yvv46tzOSvvfpJlI0Y
htZf7mq/FdF8u1OmMCutRJJo/U9tDx1D7G/baBsP9Qr45bTVJCwEMDlNyeup5yGbzutPKnXG9kuq
Sh5vgU2NbJeDKDiXkS93F/QeWmALsosnu/VRUP9B5WOdrHJylrkvw7YqRzZCLdMp9NYH8MMTHB7a
5QS9IpDmXm7dcth6DGMO8DSJl0J2cPVuyNea8T+zfqVN7eg6qyjIo2LyeBdpayDY2s+EEh3KoJBm
WznI2kQi9dUdyCTC7mXOLkeM6ysTatZDsNMUCeyt14K6Qkb9Pn5z9AKNNTCB2B7FHFmTbxdMRT8T
eLLySHC/CGUyyzH/HyrnFNRCOXHjjthEl0/ryTxXUBtLKdTHn0YOKKA05uYJcjVGksor/0wfFiy4
wS0XjnjIVmbKUO5Ot4ylAx748KNpLPAUb0hIeGEGzesNz1QrPINsCjP0LJ4VfiVqsMI2bdG2EH45
G7G49869RU3s2HZltPlYIp37G5V9vBRRqBJbnuzfDwNhx7+JaUo9yKcvmztqZHD8Edmp/acuUHi8
fs2Rbnejsl+3A1a6KrJSv7uMl17ya9bC4KQA2fJVREcJNRc7fsiS903ad9EyToZ3oq2UUXUGfnSc
XRVxWpWChGKzONmXk6F2hvCsQYK4nhKRm6JgjJizkzAJZKQQweqfVCt01AFtPsGqJ+iHrR/33jCX
HanFSYlk+wJmk2DQgSEFy8dbWGUUJtgryq8AkC1rnxSotre0ExZk6LUDa7+obPSIiD5GAMPWlehc
qCQmBGNTafH30aZDZ4TT45X0Sw5FrT3DQTwNMjmX9pgNWmgQoVdILEPH/3AcK9/dZfAKKaA8Xlsx
1iQDrVedxNo2QLHkDgkqZO09luXMIQWKo++fzvjMSJnDQnG3ef+1rq4IvM89E0+InBCyP9TvfwoI
oj6HyY8indoXlasLH/cgbakdnWVrFZh1LigzZJhWGcP7uwOcYGSW1Ulta0et/nIwwNwXtSyYaW4y
w+mMDE6MKEtZbESFw8VUBspLmQvuSPk9LGM6N1Wee1N+HEznaAntCiF6w1tU7Nb48qzZSPqyI6pA
+ZkwA7naRixu9RiU4qGPXMvc1Z3Jcz3/0FmPvD8VtLCbWdJJq+aX6bF4IHJgnnKtGUjYXBnhR5Ve
YLwWUBn+mHMm6Wf+tE/WeBvDfJehgQoOYlmCP304g3IwgZN91bLa45D0o4YWP9YxAi8dDpKuOGvL
h/2wVQDlqoSmcNB1TVlAyZBsslcYAapDQ4GRo16N4clJoJb20UFJsUBHaubtVFLBryYQBwkCSReI
FKSCzPRZHntHHBB1A+6AfmJbDI/zM1JTaaw+3SFF5ACsEMyJw68rkPpCUMQJ1yEmGRgfNVpmob9z
JMS0Ld8TDNmTlQOYpDNxExeu0fyZYC4thJd4G0zEYdov5gev0nb/DzmnDJt8miVbiU83up0wMBla
8hcp5iN9d+CcYV/ZfPGlp6LMjYwpYePYjrj8Vs9c7/B1H00aCuFsVqdTIiXQ6tHZ7wayJ7GGtVT2
qIrf4U5J280yKSyJFFoyV0+WT4hjVY4kWWLvk36R3PJgWlzGmFxTqulx4WvYYpjTrjTLyRpR3+p6
t+3Ui0/STH2kp1EC/rnMBobjtyVztb5EeQ4uOvBgoaF33iw9G0e4bBgP7B6iN/GesztWx5nlM+zf
JmoI/aBKgnwRvPUCM8mmjHvg/ItkQ2QQDkfSM4QtIDi3Du9I2351ASJtlnwCBPNvUPXtBxqx83nK
EByXCg4CZnqoQbQPrs58TW+wryqjYfApaZl0smhZy122WD22yvLw96+X2sU9oqhvguDDayKGd42d
bD1aSoEAJoxE6TcvvZ5DOJPStDlBFyGjlR4HJTjN5guivjb9//zRjzcjpmCXn7N8IACAuKDJdLFu
hBodduZqSdc1DuLQjWC4e6cJQDAMhNMdA3M+1rcCZ/GhVRQmFY2bSgpDLcNO1iSeIgKNl52DGQh9
CytCEii73wavICFXuGaF/tNbNAn7KR2dUwuyeEj11+gLu1C1pWvFN4YFRc26PJh/rl+40kGQqNEy
FOfwErzmPy6z8iswflcipqk3Syf4rb5yCpKxrVN8Fj+wAPRSJN4xuuGfrmEmFzhjQprMqstOCtdp
+FbhUgCocUz4cDbbb3UHuCCFr0dFx9iIk7fpXvvhZQkXxVbvQ2RIpaqDkKxg1DXC6vImQgc/7prT
Tw6EPyYrOxwKP5i70tjUjVrrxbrzcK/My7CRru6U+CExZBDMjEQTmH2c47I3hr7XOcM5m1d1CdNm
DSehCZGZcbcTMz/7/XeQYWQMBpjgwfSI9nMZ+KzCjSESHR8nXTly6pCwch3UdwzwmVG1hT26Cx+P
avhHg1ibN4rBd1GsA18auYlQoSOvzr4w4nWz4xwL3BcgJAU5mIBsaT6eS1Gxs71En7Sp3sNzpIDr
AJz6uP4CtP7wDQkpUm3BxWn49fs1ruG6m1H48IN/5r5AKNR40UwZEYW4bAJyijVZgot/Tce5bNUf
SlI1WyRlI5pUdpvcoVC3HINBN4Hf0a6Du8xtKJKOk3R0HHebI5EJ0aUYJiW3F0ORNFBqfWFeiWp9
BtUWIiC7LDmRmJ9WwDwfOEp9K3Gld2z4Rh7rWLSsY3oZDNW3tGJ806qurxDebhCYWBQ1gGaOStgA
yPyx2Et5YNT+C+AW4nbgphUA0seaFPmDZHlrU3fevRUHtPjbxPBg/UWgo8GcCjIfpmhh3x3rnRYH
puyKXhS+8Sq6a7Sg91TVqq585bFE4dK2m6hnP/RvTlXMPLqU/pGqlXu3mAoPnjRBkkBHKXzYhADI
6F1jRyhmu/KqyScTJVwfKZEKe504Y0DuZg5L9L6vkCHZDY1nmgCMhveyqmLHv1gspHeCVtxegdbE
8zKV4e/+qiZjyh3VDV2r8jXI5fCps5eXFG/jzX/rlDEpUCX7/zJWcyN5v72Ln5VFYPXw4NXK5u5B
LF6iywqFqByAwBz0r4gwb+336FFwlJFRb0PB38RJk7XDTMi4iKuoO0tWgDNbIoim8smvf6aMHLgm
p9e1H1qzFULKw4UuuMoY+R5hOIUOjyAY+WGzvbix4tACD3AazyZvdYBtNk587hhvlaRV0P/iUz2Y
8rNuOcetREkpIFv8OUxy8J0sgSP8Qi67lE/I5IyPd2ndYMHGfY5UcsJ8g5WA4Yl/qMZP61YlzY8U
/CRVH/AzhknSxCkDPrHA3fodFDZcL9Fnt8pks+JJjiYWzCi6xK9Glv1EVHsz1IiP4B0GMWZvdDwr
DI+F+rj1sCYF/nmjlmW1iWuO9jDzCDjqFRiJlHIfwpUnubXHj3lnEsq+VhjU0as7+nfyHzwn0szh
o9hOH9vNT3NInnGgoqHJpi4T8UtGEJ/UQoP2w5LBwXsNQtEucByt5xgNzuCM3NThE5q60tJMy7Qj
/WefIOTiROR+dbVkAhs2xdXnRneI1oXWvBMP9EmDM9B4e38XZHWDkBp/dRFKnzO/wWZCYTE7IcBT
IAj+oi6nNr+ftuWdDPNWcyeh6t29p8GU54PVzceVhPbi0UCtOiUnZ7dI6ZvRGmrA/bCP9IafTbvA
qz5cxktyGRBpjnpz4Vs/ze2kupY24QZzTo9w44gKv6OQhMHvsnghl/ZT+tdgPORx5fsQd67pyQJw
qX0IpPVRcuVvJuolxCEBMWxXqJEy4M9kMMAWDQUH28pWSrjP2N9Rjx7JMQeCS33Q8eESS0pwD89O
HDmR0FpoeBQhR4EISV4yT74/NsxGtyJ7T6HYgMy7LQ50x3XWWHgOifnFc9vkFpt0z77WCRZaMCEw
zYGrOAHd03+uuXButoc8Sh3aRjHW1QSDNDjMI7wajPOu/fkETFvlq4X7bnk/UWtAl4acHQp5/EXL
rpFw2iS6xNcSXxG/E3dmD9N2Yrobm6Y8Jr+5GFH2DMU7RPizOPJJgcAeC/M18/7agOyeeVrxSw48
fXSoyszE7jQuRTqYpfJM2EKs6hS3rE0e2iizW1jPL6SIhnySRkxYlUbmLRYHKQSlDMWPS3PdR5Cx
TY2dOTtIOH6AtTAlgoII/v+86qrSFFZBlIThF1HtZEI6EVmXqyaLWdxFenKkpYxZnLmEUBXK7p3+
CnB7ezCZ+hPn0CdodVQcquoh9N/HNA8F5iB0EW/MCnK02Xj5NzFUUT5BJn/1Ep6pHooUa8SUxuIB
3IWngfwhqmMLFRjmH+KdxNKOXDdrsNUQ9naufXe4VzzzVyaxxN0p1zrkj6ZtqR4upeiYdiqQCnwB
UfliHFLR4m3VWngMVjIV9HepS+bkjmoTs+IJ00yLb0+fzsMGW7F/HafAwLOYPhZQQWdFYy4K+uqT
0BCRdzAhK50MXxeMY1duCUIH7mJIMgkLIrALy388zewKtforpfLDf46f+tOcu4N9tdGTom9gb9dN
5ovGUlE31fthnQzxJJaLbiy6w6qKS0REx9smYl1ljmO3YPafDlq+qOb7efcM/tIIU3KL3jtHHYnm
wOT+AjrFtXeNKyhL5i8M4hB13cpG7eXue8xbqbw3h3wkbA/Nt/kdEmfnCdErdOyXUzUkzlYYft4+
pb0e05Viv7LL84xyH2L8HP2wT6AEPMSMrhSle8qLj0id4DyCFnFaWgg1fc4+T8Ibv6vg9qcwkfiD
2VyBIOwqpzyjJYOaYRU6rJlHAI8aT6AoD/wTe045EcnZnFFyzTp8kRKnyAUk+L02l7ssrh2tSxQo
+lKy6nmCOynFOvwciDA9hHeMiz3vJAFDBKy0vdd78Ka5cX3/AbFjyHZ/rvJHmp2pfvMxuD0xKDFK
rDuMYZ8YsIcCN0bP8qX8GxD1Yz+Qc5og5ttE+DXSUUAp3pQDFMQ7kicKS3Qsn1g5mqY+8FuQKPL7
jhaBabtTcsuXI0p7827IICib6SGljMn3ayH35eanHQCyM1z5o6ImmRuKXD5dcSJ3WmnbdFyjAjbY
BnMJaQvxLQFu14oqag22IX9Zt3MaCkQacTWjs38T8bI2mY60exakGBmese5wEys6eP0tLF4aZQ2k
MNBRLKUO0WKk+S0YVomhnrTyYf0yEFcAq/KqEJJYupEnNI1ocGgDr0ezlUnsTW1uCwpVLUb1facb
BrhOvVC3npJc30kqUQfACKgSXvdEIrgftTmUO0DM6pP+/w4tyXhR5emgiP4q0neocPYs9yJZiNO+
clhUJKSl5rJJfMOQp7pMllpFoxprGlZa1ZEaKun5sADQuMld/Lfi4vLymQy+j5pSPlauiDwevuxG
PdgqPN3na64NSzy34TfZ9yqpeq3UikEGGHo2ud5rUEh90B0NUnBv/2akjlbLHle8QSEUss7RRrqD
VC6cNt0GboM9TjJ7fUoM0qnyjSccHJPrXhK120Nqj5DRwwfHITLqiLYwX7WDwsKeF1ejNJse6BQW
Tnxn93uBAUxCEpqsrQ52o9WSAN4zS0/8E3xlINv9aXmDaWbAdiQx+7fFE9b5z+xDL+hyXQXWtMCE
JLxFZHAyel35fX/PpW/FvcBe7WlGVEe+a789k5eGa8RVbvfs653gAa+XoEzLHUhUklybZab07oM/
P1AT/KKDBz4OIGg6of6eqYtGZbQTmz7/wj6hcYBg1Yx36elZZsp7V6pU6VMMhQ6//bO/mMMqmDZW
X6u3yGK54/vwgAkMr+jlOufhYCgAWrCQOWEp9UPUNjCsY6VWdP3Lf493DUCl1UzcLVjhMoXotFpi
mMCDzEh3nhoNG9NGP3VNEAM4b1PE3P7YCe0ge3c0Jh1kTgfTRTXBeYOQ3i2C7LX0JUMdSw1qE5pe
DTiIjsVYeSxtROFS1hNTDD14FI0nL9VlDTJCVce6EprB5EtGnAvcnoBJdNf7IzueYn01lZhUNNv+
OD+EibgGQhMUVAAkylLvyGi8efrCbrRIUatNOv608RXKgPIlMDdYexszkiseAUSTyqNiQoti8rMV
NBc5D/2ZDL+n0aBOM/nJh5pALHFHgIa7z8cJe70/zsXoC8PFXKNmEH/5E2vJEkQr+fNWBBeEJkMq
guSLq7j6ERhFra4DBOvEOXxtp06NvNJVm0685kRArn279HZ80jVdRXz/+MJU7PX/twvKcpL7PQVA
7/yZRVD+Sz7GjWBnBKNORvMsriUBjcEX69HVxyLTFzH6TzSinepKN+vhU/BL6sVIqFwrgBPutw7P
zzh5yiyWAIbDBKvCrlrhyOTJg8Z++n6a7RrAJb2mnbWCNv2PEee1qdTBKrilnF7KIOGL/Gs7PS2Y
yY1y3UBFyDsjkjXsggTC3ENArfQCXjXHkyo1QRAcIRbR+WTDlPauuxrHBcl04Se4w/WiLDvB1Sik
/FRCSc166qExp0DE2YFhATIiRnKEsjM5S6Fb7G7Y0nSJc3ksNngDlYqYfrleJZP/fBH93Gaf5BFi
uXWcOPUtVL3FDVHgSjqqfOjKhyiTS6wIGdAxIQQy3/0ZryHburOGg2l4aRXw7Tn/lN7yuJWTpw1Y
lDXuo2E/an/zwzIK6pfHfOCUbFw7UDH3raq3zNmUHuvCr203SbLndBsnKHaQzoa3PyzHZLBCYSda
f6pYaovWyohZV6du47uZl7oPdDdB2wuHKEEFM8GLnhy2TdWEwVcJanF/vf5/33oF6HnFtV3fwJvl
3UDUDZbi+Ja+cNC2G4iKX6Evkkkt32QbOVatwoy9EuuofNNefXP0juqyXz4pJpKz24Bta0UCPczY
T5N3dAQWaYIXqaaZ/g1srTjPnreLGjQBlDpZ1dkxsxSNZUWzdG5OwmnHws7zM4c4gdZvNHHPqEZB
tkvBH6ZYKTjJNjQncnF1zL0313G03ggjHKgPdDUJFz7CEoQ1ofsyO38hp8kOW067KXDJ9KepOt1Z
C1SuFMjIKlm3ZygfbxFACYjJlOGqS08EO59225QuQK1MrowrarQt4j0S3aQAZ5i/vTJQLFFuwxZK
wssuBpkF8zfcJ4jcKby/VfYWl03sg2xl66fBVgoXm0Qc+0zxl4nYeEmlCdZ2Dvz7cfOUvhks0AWz
nbQJFZy3ORkyCiMffUQk1n/DasRb/uWeSe+xVQPj4bAGwoYsIp5blf49kOCR8XIlc1Aig4KYF2dJ
Cl+w1RdKjmhhiHSmB8PG2xnC2ZzuV50RDsHvEaGdKIzQ1RfkOjzZUu6G7j+FAMiK+/MJyHYFe9wT
/zlewpycpfjXrFq3czZEcPXap3PSHL9ZfGxNaTatKldFl2JNF/8QYsA0FIT441jEUrxb0u0WkFUO
F6jLPmKnKeSpOWQgemwjzeYfd5DIsvN535S5drN3fDooMXKDBH4SJb0RCwubAo9wsAUZF8aEdcEw
fEJQwxoPIqFbn5oiHMMwNlv6QNNYnD1DBxthgpRAV3UGKcbK6wacpEWS75SkVkwuVcaEmWJ6ihLo
JbGmdZMmLnvkDoWLpoOvQDeaj0DdyX/YAg/XSen1xqIZK2xA1kExca6s0ZsQXEvDNDM+HfoZQooB
0kEw49INf9qVFAy4m5FPN8nqaZbQVLBo09rm+KdKciVbYPy+Q8/AIcavdbHiRIa+VDuaP/wuMR1F
bjyXK29pfjFzkR6dQTR/7dQK8RoyunXhonKEdlYjj5jtRqjI2AIpkrbObp4CBsFH5ksMPQDN56SV
uAJKhGF2NBbWfAhLIy2aAqTv86Pfaz2q9c/FMHJkh/D0zLAzBIjmyd429IswHHb5RQ0OI5tAA0lS
0a2HrRtHfAJr8lLuUdVhjt192Oe3fyZQsPlRsMf+cUJ68gd5oJWoUX/gNybrFbmTgOV9RRi3orej
gDNNkxl3dzegePB1Alkj4UabHeL5MZFzZZN8S8/JNmXBCOWY9RwKvyUeqiqxNVp18dPyfRoufSvt
i/sx2BVYUpB+9v2Ih6SUEvGE4d2r6QXQbiUFN7UGqE4aacdrgxs9DY4Zw0o3bPHIbtNbnS1St5nn
/RHmZpad9lNIpoFeq0UAAzPZMI9L1qotHChXXt12ZEtwLxI01mq2pu2sk8SBiYlA5pkPp2YMfAsA
7sjQAeCXU5Q1zxh2jd8CEI+pfN1nG3TqT5eQ0GKCSaDswfTwggI0mylCu63UOynVMZ0XC4iD8sQu
0Vym2sUJZiHYXBPCTwC396oEA5S/YUdzvVJHu+3GPVH/euawMZxvbwtTRrHs2J1TsQ2JLz2hwlXI
6gZ9W96jtxogPFY+ENdDdSdgAULptO17MkdNOFHpkXOQJKSHZYiWv+5RQmNj5NXuqIgtI/ULAH5z
PYHzFib+dgvD4/vihTm7U/zJUrvQXqyVYVS39DEm8q7Ya47GrRbmulXpleuaXHbcEoUVzP3KD8iK
ruRLUOboT/fNz8idQFh1Nft1nbUfnQUFsAFe4Na2ODQKuBkwKbX44jkUPhR8cwflC39Se07aMhFc
maFDLozdjn8FInDDp1XkfiCT9hhk5oZvBg0GuXBUVEK/Aj3j8EvBbBcMxNDOBHKRktlJeATXHOvg
TXriEpD3/oIvWtI5u0/1bavXkenenBtpo6yxRRu3x7Re50V6pF4tuwrc0OxtxtgqNsJacUUhRpvO
nwmRNyOcCMP3eRpI/xUiymVroiUap2wbiHrJOV0l2nT+Voa2aczJa1/nxI14kj61Un/GhliBZyoA
PCXijMw0VKcWqGjOa3JccFHqxkoL0nXqDcukP8JpnNDGB6hu/iFowdAZv8LdC2f0D3qTaRoy4d1y
JKDP3rFhOPPRKj7rFryqIO9dKAH4VG6wLnDz75J7Q1LON6W3sj4oaDoDwB5IAju9nxgMraIDfnuJ
9nJs5X0TN5weUEXwuLBTnTcRs/4MQE2SaDbxbFeq6H+cn5Uvb+rifxqfWFFdFKhK3gKyGZ3PwBck
D7zS5vNCEg76IibDWzNPtYuktXbWZScZhP8N7UpjzTdUOr3QSD7qV5aaHZcjnLF9pLCzUBqL5yJi
5luNaxks8rzevekaOsHh+rJ2veDbXPWDzBg4+cQqZ5qEonW5LyBGK7o9hIWb2mr+ZZRqclwOjNvS
4fdmLZ9aWmcyH3sKekdYuulQDE8KEAnb5jNRzLy18liXk4lobMrAGVmLxvD6V94agVPBnCGpuDvO
errcF+yM/0cWklb7J0/LXILjKywQHpIn0c5eRZ0A7Wbsfx5/gkhwtN2oIFPgO4SmxdwxEdztAtWl
lACB9LGT76r1jG4HWLkM9BSL7JezZgPX59GogGLmyPrz+ZVhb3Xp7OxNatbEqyOKG8iXyikd2qER
HBfAzCTRRtDLXeiocxgHyiOJUVU7aI5xOqeGFB/o7WegadmveeuD4+R0d1pvPvLs+N0+wZTmqCcc
ArXtdfegAQtUEuD4LKxL456C5X31uKMRSURSCMuswV535kDah7fPXZPLOkgbPON5NB2baf/Mrsii
tVSRatJEWWeYQJtG7HgOLV7LIjnWgucn3CMjeXJk/2s4D9n3EMwiaPeE0dG6XQ0gPCoMK90Y3utI
ab1yR1DLHtRdK3muCqdIOPIw6QZovzVEffKsMimyBqqqk2SYhpT5BGurhCVQIrFwKK1mAg+RICuW
bnfipYKsEkl3z6sUEYzKzUDBMYlctcBps5BCPORAENbexdi1pRLzxeoyp753qeX3pFx43arMzUJC
fq9DRsSDWePZ9UdjLgC6JNdxX3APdH+2k9M0w/6UI1ZTuejr/kHxVbDp5I7zvqNqgj12sln4+H3/
RFFx3Id9TX+ojw4jVO7EX/IQIvBGJ8Y7bZ51XSBh3I8BPRa9n8beYyEGJMtgmGX5mr55uiGXKF+M
OkMMcSav8Tp8r7sYM1+5w1csVCXzyZTfA9CCHatASdUkTizjGtMdcWUDvIXSf+aAZQwInxWSL3w6
ohL6j54+EP3bICq6vi2PDlMP8LzDVMMmI89i06W44BOE5Aq9ewLsGOrCqCh9njLbwY3/I5HJkRtG
PblvZYIwgiVFts7Xh9EpysTWrT/Zrhc/zPj5iAne0xancPdzwh2OHEdIIPmWicUSz5JbiWOdq4QJ
4NC/LVfFP/xh1e2SyJA4H+9RYGxCSFnUxzcQJmwLXyqBq/MJa2NvkIcwCLBPVZdYLhy0at3BfUru
Pn2XS+pnCP7SvTz2kBBuU9EVLf4sPfUMzfUA2nlkX66N7f+iV0OuowjBC3EE3G4xWfMglf4t8qZT
tXW0sGZJJqujAj0i2aHI3wrYW6HhWdQgh965a0MPMOOstdTmkZ5FAHhLHZPEeto9lt16yPRsC9P+
xpqI+3Hstl07EZPVbEPp9XhX6VlkkjyxXriNOWIoAtQ5qsw1Tc1MgRvXunmncUrTQ1aoC6DNmxVP
GDM0rac5CdSGQgnwDFol8y/l9cQ9baMmRME0quAabTn9B9fPXk8A0mZTYawcF/F08j0g65Iu/weL
zID98z8s6RUE5jcQB8fKOLkejRYQtyDg+2aJ9SM3+raYS+/uLaaTsOlGRgNehMY1UqAoAu92bSy2
oEOu0IpwW5VivoYUPEzVPXkU5pniZRbd2PpPrKJVSNmqvIyUirsXCCcH7hmxleD1XcDPSay89bmN
zWyB7f1boNfDIrj6DMnWKg4xzvl2KoMHeiU451Kv4YkKtHUCfAidfFhY7uk6leXCUtnRuVRD3z2k
a0uM2fBIycGFLP65tDaty3AYDL5hGAW8kKep2bkqjntPH3WycBwnaGTpyzJtUR2J3H08i0PtBLoh
IOTcKhvB2bvUhZop9ZvmdGfJGMKx0+36qYndMFEM5IR66uIPuhKzHeGlxqRrpqTrod6rnSK87wFN
Afb3Azz+Rg35KXxr/qga+h38TultEtOjhKktMnxhDMgX5AItUrf4cP72JzcDSZL3Xnl0bfpqAFiK
rMaWVLp2zDnNgC7UYKPKjxOgf1Z3Ow7Yu4L9sVWsI7RMEyGTZU253x3Q7VuaxqCyFZ7e0ssFFt3W
iaciM/FZcvuSPW+v5AVTXtva7BNcn9vMHBKCoFwwhUIEmrba2u8dWnoKK61q0OWo1KEYH8Dd5V7t
UZmV21iCwB3HKCniMmYEuJXaEYwmBa6hbmbTSjsU6zbb+5TYyUOO/2IJvPm0qY6D1aOnoatnSqbm
AzqNkMQW919TLSbAo+dsRgRLV1hcILIzwkHItbNCbooS7P3LRYo1+Q3UhLHoz0v/0RzZhc7mKCv0
w9EiFBueI2Qk4M1NwXPvUP2Lia1V59WxNKIEjLddU+gpUPpGM6/fG3IoJ1p5TULEsTlZ2fsCXbs9
t5xdM0Bn94MG7FFhBw0k0IRW9LqKCH35g1onBMA/AIRXe+jzAKDPVRKkHc8U4lyF5Wvg5atwEd+g
LzHiJYQo7MyYxLOKJWjb2fcT+ydSazz3VjWjsYR3NgfUwt6ZvHberNrJLUZiodNNO7ilBL8ZSuz3
EYwWflTHETQ7eCAsuYjzOYUxbSKWtXYndtxMfeER/g26JKvd+3jJGJzXTiKfOI0PNZMBMTPQzoxp
JFYt3+Phh5h/Vupiz5uBur/dECQvwaRGQRDwEjAFcf04XKUpKksJkv78xOsgdOiL+aL4G692bBIq
LGlMpmPVpOfWELXs/ChhcUA9mXZGlhwc3bqC9gxKTDNXiCS+jnaXzCcsEldUcehBcgW0zlLLPT0l
oUM7JUYXp03UP/AFnHwuRGDQt+83UdKVBW27C8JnE4hpmBo0RYbdhNCxLbMvhGUgh32HsBCuJBfk
ofbI4dXHooOeskyQrciA7T9PAQ39bm/cQWmWV5RcSDY9k/AaiqUTkcXfUyB2jjk76rcGowhpdA2P
L5s1ohKOUkaalyFwEGAJP8gHl6IPIhYYQyhPqTfKp0kV6484V7zpTmTnxy4O8onV0EfuR/t5F7Ml
XAor79E9KnfW9N1RrQgm7b9DNYvXku3g//OqDsTcjjsYEW+/x+3urmo+M9GyXwjbSApcF2gNmQ7n
uqfzAum0cjo1nCh70PpD7RTvBquf4AeC2nI1VE8oDkyzG0ckS17cOyIkcnwXxLyx3cZ5la9bLRu4
vZSCgtj6hfeIhLoXz9/y2MF+B/CyxTXGYfHS+DTajyAouOWyUgA8l2+PH2WC/lSDzwUChp7lDYWj
mzDF29HDNe+QZXF3ngb/QJqsD5BY7CFqA+qZcSwqur4qnCBFmYgplOIfzEYo0LXZm7GjZfwx6eRS
XBsYFTKiRUdkWJe2jwC+1lUzFuG3vpx0XqLu2yhXwP7t1VzRGzPi0CEYiS19jHsrys6PjxsO96kp
IcuUOzOZ6a9/KkEjXV0Fx4wN0/L6woyKyjclZV58d81GhBULNNRwbCGQrJHO56IsWHv5kJNO2DK7
O4uHv+W7rBY/g9SFmIsGZq1giVFWqOZofAuN9jdZ/dKp7U5wOnSJXHe9ea1dHTNSxezTgKVOZEMC
sD9Z/ryCpvjREjuUbFPWYIjfqlDdxExo7SCiVfzqMPTp0LAeuyeUaRwp09KqZSFwbNJivZq9oyXq
D44A6puxI2sdW8jYwI2oA8aTo68Hvfpu/3uCfexXbWtY9E1iYjL9ohpBO7jsR1MG9Dx4dj+zmAtv
I7YXS/h4IpJhnVu0yrLqeaMuGedaI/OdOlruex8NE/mmwECxulC5e8RSt3KoPq4ZX1ZQbXwJdJ8E
haWAOoJqCgQSL2+GZSz7NJ/T3UzAh1rO6xrPcruiZR+jD0PepZFEHlW9LOOmVeDloMSanBjiuF0f
iLuuFuAZ7BaaTqBQhPEtyAiK1GQR/WXn/p0jcJD9qyQvt7CkESHCUXaKjJduXAWy0TvD1YPbcQVU
ZIHcX3QWs/4FPjiGQFIyZOFGJ0USxMAIbwFuEuHCFYU+b5Rb4TlAJ9CL0l5+VT6F5s+Huiev7w05
aBlmhHXxABSs6iakVhuS/pNtxDFGW+4shME75rpxxiG0Yh/WnVBed8bNP3Vmqch2x9lmKEi54q42
nbYpiG+jCzYyp6J+nQ1iGbWDubKSopE8prvJhut75B42kXiJrdMzxC1B7UEbE21Ms4T3mXBer2S1
CZ96m6Z33prPYCffSdXDLtEqwZUT6JlRtqV21WMTcJOLqtkPU2KmW8gTcgke7GSgN6GUl/6vuEN9
ptfpUHhjJzz+txOzZiLMG3upx4N9dqUVPH4R9MaF6ZSgDBRO047qxLpYkgtZ8RDbg4zQSLZHllaS
oREEwNIdvebglaz0QjYJFmy7IAVRDR50z98+v29A3chTrD9lniejL1ldtxcA472LXxSjLALXDTah
rUwZqyHRxTahMUqO67c7ni4X7AygSyIrtdtgvhOmxkxnIocbMl+OtZhfBZ9j399dKbLdUgLbjTC1
7ltBOVn40gJ1bkfDaSomTpq3zz3uJSvhovHTcGOdTOykyUXlZBN2WICcZjaxw5BvcH8nAL2Wh3wu
Psl1RZeSZ/QqZOcLdg6EfVSRgiy2BZiopizAjgk9f8qHkJ1h5ax1UbDB2K3lGJAxZ6pMlbKOk5fK
LlfHYjCfiPg5t5AbQ6L5e7yBLiLnaQjb4LPZLOD+cKo8WJRCe0GXmEFEpSFJucLJ71RlnJgYoYLx
AwXVU95s1UtQSh3ORGZjshcC5ebJTgHXsE4BYE3eK9G2CLzyHZ8g98kpx35qbUPHzBEm6uAdkevv
gD9WAyqqJjnMoS5tNG2JHjKedhpdOzZJqA6tS4dbpQ6lOR/ivEV6FNE4ZolmzO7p3Idk3JX1Yf2g
z7A1myRswzqPO88N0K9Yh1G/3uPVVWa0epxuPVz40B0ooV5hWyJPoh2kHhG+u4YohBZyz0lJFqFH
uY/q2h4uQLydoaD1eZyJgZ2zwoG8xHGc9YPMqBFOQqFukVnmsxlA3SKHKjdmM0a7VBWHr6Lz8LA9
+PepLp3+hiwdbIDVK3xnPmE1aUWU0n/XuhA62ajQuYTcGjhv4x7ftIorD8JWA9HQ1dR6tEBhA5VH
Dcze3aUo8tHWIzxgOMvymZMLet2E+kmw77/gaM9nHzwjmKIezPvgO1jQwCbcnl10HMNVg84ZGWCf
FdV7T0N58E1dh2BTv3U/TGB8uWbS9m0s6rChbBujOy2u7+tWaDRIMwuAvbvn2u5yh/+jCnCtTkv3
kEKkgYPj1c/8oD462fw+QvSaS86WrMuEq/iKMDuhMVFLBoawSdYO3pEbSGYDmODjyOgfns9Ga3Th
ozxhkpz5aHAahi4GRWdRnsBrMO2U+9TdInn7lrdKyCKnV6pnc7PQABFqcTAeYxEt5xeFKPNqIOPB
ujcZX/Y8F9miiyzFMGtusc1fgZYtaVJ/OCosZynI5e2OwfgJiNhtEezVZZKZzeMkgDDPi1D8x7f4
PZc3WLZz7HoPJGZZG+qHrTFSUA04sJUyespWHi8lDcAURmLFx4ZgUHv+OOtW/Si8UeZBCSjeftjW
jCjy6ugPcqg1G9ssi8n1WTccW7vc3NWzVTkrJZ4C7LQACtgyowJFlacLmtnJUPO8fQoUv4c93zxm
kmQ9Gt6JrB5OovFBw/UxKwMwDVDqzAeX2PeM5K7DHhSEFACFCdj9gToX2h1Nr7oIl5ATmnUG82I1
VRicPRHPWQxa9gSYgEZ9sPV8TdxHwRdWDDd+J9vlHGSrb4WLBaspQuny9u3pW/Vs8pVVDDNHcyIl
v9D9SUMqrj353CGWfzR868Er6Whimq8DDWk+IYyiw/EXYWkJxijSVHF/5oIG3EOwWeYH1IuaxQfm
8RayGIM3E83QxDb8ojWv0SWJsPUeSNe6SItG0iLU+lneryjSgwgeerOgYZHk7McfaenHKFx1jjkN
tt1dozC4uJ2DzHQpDkEk3L1fSHvkBL840kSp65mVkskJcc6dj1yuwYEaCLwzh529KwyVgaSVVFrH
iOcbOmLLJwBn9MecU2s8/YZ6GcUqowiRJyS8sa261SGgMBGeSTIRECOEn0HJsHPEJkBuQcgVLK/5
Ib6KEjHRQbgS0fvPSEwJdIBxwgd9oGhRYe0ZnYd9saXSLKZ1eBtw66lAJopiZXR4QK0ITFgxfUvM
GSZr7WethjxxL2JFGP87pfu1c4PWhi6NTbea4WfYA6LLSWnNeaDfTBQ/MhUHW2yFXAEPUL5LcC5m
tG71uycOaDwZnuiLbyAaHD/6MfT4lcbj0WyQFyH1noQ/fvyFTvENxCJ7TFnxx6G/2CLLbXRem4ns
rXEFH6B7SLBDEdFKWZY2dS1PeSE28DIQFID5ORwNCsi+iyVP2LQyv9tjMkWFuj9tHxAzaJAYgH31
34qvPaEPqwp+UNLcDDCYnMG4/l+3nEyxR7/ira9+HDPKcaGwr/F0FPw2RfL41MOH0kKB0afqr3tp
aRC/rGsLuXa2n01xmZt9tDAhmk9sk84WQlH46iCw5A5cwwIxpDHeLh7lwR4QtTrMs6SLMFK4rXRf
JkPRDjcW7msuwnZ6Ps9E8oRw/2FDMYZLquXAaqKiS/UaFb3tqZ8FvfHmt4QMI6TievN0P/wuyQ1j
kym3qXigudxh4f8bNokd2/kcGipx1Og60M9IIV0/BIZG/5jU4JAhToqIMqbJ2gc74a3/DjIezVlg
JY1f2LKlGN9oNTy0ZyXGAzQpRx1XpCN7YeOQqOyfizUuR+fZprioY0ZDnq3ddIFl0fdVL0xMGkVn
K4+LGIOVGfIza/rIB0ZR/z7lAOaYzPTpDSWNVDGc/0R1dC0YS7pkCF8N3COVPpuxI2Ea4qeJtm2O
AotHbG2SRRQVXDvyr3/QhK06Nj2cGMN08HucANKqujjZu9k+4CGQElOOD4EN1gfa+mO8OGLtfBlK
9Y0Rm+gHUDGbefXZ4bi6s31wwKi7kzaE+QhCo7an00lf6kOMlL7xOGCXZaJZ5N+Zvo4s5+8MICjt
61K/2WAq9n0SaBGPjL31sV38MVkniTQIiHSkMZUe4m3UzQPRt0wQuKqU/NyRAg2II/lECKZ9QnwS
gPSKgXCDzPQBZSiSZ3f3C5Z21zcXED4RwPZ+WIAJcshvW/qDmU3N0HR7B/3lAwTg1KlPEOIDsoED
/GgYX/DDyrkg6k7giDLqa4vRzXe76pIMJ7KB7AL/99hOCfsVFoHsfKjKBJcG+qaHbzp0zj6N+nvV
S1IW1P8IFowW+0RIWigKb8VPFQJ+ZayY6rLSi9hw03mis463biWNGmmyuAUfvTZngUGi8WgceacK
fTql7UqZGVJUhbtxuZTfIhNl0bgJWcXRWAVpDlYPuG5r171p/ghT0tfWcG/bhZdD8gxiolToK3qt
8Aba+Fcd4SswYPwZrJCJaFaLx5wyqTlOpzPik9zRpJKH3QEvqghjJeT49jupHYUBg3y2EyStZXxx
syS5+perdMf0W1eeXGjWBznl/12CnuQXbheqGLsjdSpxvRzqY3bE+0r/oo0ElInKGey3nHrg9fho
uaMkDJrW/7WSj/Wm9HqBv14MbD9xiykxbtbLEnQM6gCnu0Lbv00774aIU0FCXn6AaNYtzeUQJbWf
/BFSfCuG1wpoHLkpd8qO6CLUhumWAnhjP2lWrNBrWl7Sinbe+86jdLw5gEI6dJzc63/rHiyVUMjj
9wAXcIMC0luPBFVoB6CWj6TjPTVEtWBtRFyPzYXP6EAsXNAM4lb9PRlAqjCf1O9LwusDWCVfc8cj
tDuHHNgopN6nHvUuMtHamzpqd5pC2FQHiryZwcEqjlm6aM4m8GcouYNJ1HfS48t3DKCqGLJeH6La
1jQ3IVTvdIURuP2WTmdQOv1H6GU8pzS9HR6BK0gtKE/RPT74m7W7O5oXV6GzPOrOQcMmaMEf4Tix
wIWnZXC7+EIEtqy7MhJLppAS1PDPfCO18xDfnEH6uVbkNLAOHJUCLJ9HYpNi3nJuZnn3yhFi6t6z
M1B9Zrx+ENmbN8cBjc5smY662V3VGPa4pQ3+8PnjTdLwwUV9pO3M7gz7qJGeCe1lrWgVnncTl9tw
f+hxpVnFv5OstnNDfJGm/uvGN4m6AbW0onpNNZ2vI+XCFptZqY4qaDPX6tzEx4eOyDkkzGGA3+7b
1pBgAMBrg5Vab6+K15fGMaei4pKJjAogvOgfLKudTu6jBT6RJ+bt4VoUVO8WbiWldltWuSwG5y1/
/gzYXOmS9Jl8v+iFZsIgKaBfWUtv5HYYad6YYbWe8dEAj1ohtjq/hlFLDnwkuie88b+XGmdBXpDE
jDOLAHAeKbq2iYPS5oAhI9wxnl6xgzv8MdJMJ1181airuJve+GtE20nDjqDh0IgMDnhV8jfxM/w6
nhK52YdUKn0wU4ZZmV32IjeQDRjuo6XdQI07xi8m0/RpAFNBqBGfaRHye4R83iGctDAXbjIhrvic
p13dm2UFr3m5Ap6lD7nm7PVyBF+CjDG+Lovu4GkhdBvp2/s4D1oOsCSOyG+5vdP80Lm3kCNFAFy/
H83BSqDdzmIRq6GL4h9lAZRCwM+S5ahVWxKEEn9HcmkR2cyckda8tZXDA9U7+woLK5JtmanZVlio
k7H505zyRXN6iqYMSEg17VG4NkD8wrkYgTVPx1SM4Pf8ENLxxJJGtZhv4yzfmW/W+aGiv371TiAL
oO7LeEiSo3HBaVkEyBq8LujNykNAMgPEx/cmm9POK+jjod2Cs309ekmLEjVx69wcetH6sm7PnJ/a
vGczC1t3Vs0aQYGHDl4BuUVAusNJ4Do+Mkk/vEKOmXQNpOVKEGjxMVoVNoI07h28mD8H4zX3udKM
hD1A4mIyCj7bab45Am1m0pWnsNKixGqtUWzJupqMNfGgzD1jhcx16PVelG/p5snvipqPgLB3Bz2O
2p1eZG75j+hacpdu6Ol1xVcQCFqaPLDgtE/VmSHV8d/AgOSjc7rB4ySePSL6IFoFFwydhCKCQptT
vyZJOxRCEZ4P0UShcgqiTUcZ+RVeYURBB+kDFwz71XJctBVZTvpxHD9iU6IdiIWUg01zr+Ryoh0Q
wM/MhzSbhENouIAVdsE6qMZHRxKGZDLCcEfLMCw/hRMW8C3RZ4EntcA21FKxKYBNKg1jhIqpwQjS
Y3y+lB86Gv7eY+qgRdJ70hW471NobMZ1OxMB99IXYx4NllcBmaqs7rjtPUgZq/QBIjMb4vTC1u9q
Mfdu5oDJAbK0VJsQnEqZt2NGtlwdMiiGwwbAvkukk9aWevynkKIF7lCE4Opr/YOr3UCVaiT0/oL+
ZFRVLwkNngsHR06y/IlGUZtvFGJ/oW7tnw1YHfYJbj8GQetcufgsyiq4tt5nw3+VnJjYhs3NKU++
FNqEL5WQO1bs9HFv0hVC5ObUP3k2IIOrIyLtUEKi61PDqr2paVKiuLXPPaDQippq6bTRCB7xLu+M
L413Q0I8JmuN7H0BegOrpjLIANUk3NwpQIVX2gjPTKKzZsY3BDtIA4LGkprjRmneFHDy2FEE11d3
fhrQ4gLgzCjob0j8U0TiW6yocyAgNdeAg8MHWSwhKrF5ktxD9sgPQzuCW0ISvG2QAGIDx193/lUO
HmOS2ZpJWWHZzMR90N5N5TR8EX85GLcka0paLjqUYFN/iZUhuGbXUz8F+vfwidsxggn1qWA8tRBV
zEFQ+Ne6F0le18xbleOIpUWP4RbXhFIoIbA31/5T/O9Oia4t2FmSFx/CvKWqpzp9/zZx37KYAMXd
SfbcaC2GmC7I6tapZ4+8iV1ZLI6b2McysFDXn4OvVeWSICajBSEYRgEViFYtxtZ7mG5oQ471fZ6c
p+31Zg2vfsuUQE6eRGYHW53fOD5HJtVVcWTMhc//Kb4PIcoFIak2fqTEXZ7E+hTNARZn/q4JTign
ZdO3/SvgC45R1NlqmTouCMuDC+wgSHue4i+teW8X8fHZ9QRVApzng7yPe1XiGYCJN5FHy38xOfms
Jx9hiMrFeqI/OcC3vnFTzH3d2T8/sGvssvSVHJHiOwaFDpEqwEjkJF5y8EGoePXXnHCzZShPneSw
Fg0PfepVnTO5WSBOWG0JIaolMHjZ5aLKq1O13ZFS6SNtKfzKUYpMYwbh5V1DSvL7sTQbA24qWeT5
1WuZG4dfRyenDLd1tsp8bjKpTtpvOo/kO/jeuQTrhNRe0l5GGJhdbeo3B1pycvzSXoliOvYjOadS
RrnDoKJLNYTQO/KvWROl4uO0HVY+AhVAE4QWRtjrYPWcsheS4eV6ph46mwIQPgMgkMJmF2celdOE
/gZMrtIsI4YghD8Sc2q0aIl8Yid77NuSEI1oNjLgoQZoH5Uh7FJnglK5wAxKX1+T0yNcFgvDYEv/
2yylz3xYY3TlgJoUh9B8fyX5/IICYHTPeVGReWFws+eM6X7of/MpQtPtCQ8Qhq4BiIwIndj5q7QR
4kVG5xLyDl3x8hru2i+FxodccUT4Tte0AZyGEPPAS54rImCRc9gT0mUnkf8/3eQoXSdGFyxLCe+B
miSKELG5ekzp45keycZWo2oGC0kw5g8wRIo4i7/Xe6JIIcR0byej39oDRuwc84d9jEaXNPCHI1S1
/CKC5igQYIHoU1PpCMMHUtiiFE/E9RYhRXoYXucyqsryLTRZHrHodULahRz4jffhs0Djf3TrCnxT
xBRQ/t5pmrtMcQ6u+tGDNGLMeGfoxrzqSSSZL8IAwE2BTNaRts7L/DLagr7lnKyq+vOygu7dekbZ
LMuXPu4GquJRnhL5lpFgAIfjeiApHcEIZ3qmenn125J/2MoghN/lsBUfFZ7yAYa0pvZOaGdEIH9v
t1I+t7mMtQk9b1+j29yS0zXikx42tPq2GP3A6lcHaddvXLEouOIXEhd+lIGyWcorEuEhUtYRbhRV
GPNSSRliSR7ki2MNkTYYELs6iiln4UjygJonBbBTC2YVOuL2vSAz6RI5Ci1lpvHb8/AqN9M+y6Ef
83ySkFXHUok3RJctlJ8R4oMySh3KFIiq+8YjOhxaqPP3xkuw7zr/yYOZWJj+5EcYv3Sw0P7ivheX
seQn4LD0OuIJ0pkO+Xk/ELqMm92yKDsiJ+vUzDSbKx3Pwu3ZUVhionKbkSj0LU5wwJInZEja5ZY1
QOe2VX9tPoDmlKJHkslWZiBfYjpCM9BUPvioj1NABOlWiTTAuUcp20MiIm3T6tsVrOySJf6XJVyY
XhGn6V3x3TvjOuahBwRA2gyJkT5SOoyl3pWcf7mv6H410TrSmumwteaG4XtZUdmrq9yDrYMmWDmA
o0nFq1snXWZUXuPt4Z+fPatb/7P9AY+YNJ39FnJlk99El9/eAa9m+E2h0T3C85IXLpinMnSWSDKL
Z/GiPPfWMkiIPIe/eysQgM0S13aJCTNsYJxV44uEL842eqMJZyV2Mi4FNxLa9fcKe03wSY6uaQdr
6+jjvNXRV8F9Q3aM7krIA/Pux0u8eYaTWY9BLZ/rHiYIPYb9lI2+7XKAcgTvbYbg+JfwJFW47dkm
UcAnJTXHtpEmb51ETVdKkuyeCHL8RiinNmr/IEFJi13Bam0aDwCx0E84vaVZsR1eqNYXg1465cfl
q+juriwtxEw7UKA58W9h7P/MzZ2RZ3vDwn9eELmpKsRs5bZaF5Wg4Vtd6ExnuyaznYuGyUdT4D2G
f4HOy+gLnVRlby1BpvGmN2x8gRTYE7Z58YUc4o7C9SCDxbOkB19ybfUBVQnueSOIDQya9gqf6HLO
2zuzhIj8zFdJ0xukOBYfKLowyaQ7BOIwOtlhZRVxPwldJqRWt1V9VaUvqS1W+gY/Fws577MA8NA0
zjHnSqcT0b1krfTr2c86YsawFa8xnDJkFMQta2+f7oTKtLlBuCWoLFgF4fOkznArKC7Ds1UwXnjA
mYl0qhcUbWJ4+tdzfPFkYDLhMNuke4yVLUEu4LVcUh9y/8xpeY1gLiTmBcmoBeNNTYJ1u3PVwpBq
5VD4cfW/i4CDIYl9YVWEmU71VQvBiD8KesP6EnhlQZo/P/b2PRho1EiGKfOkDHnI5Ll/01Qkmk48
+afLyKtPuH2IY8QKmY8siZsVcdnrzWCW84llCC1o7TwWa353M9alAYswJaSSPnWdrbxGLGNEiC9V
FKoosdNO5YIWl5SZQx3N1ZKc6U2ZR/2SnnbZGeGw9wOb/09tiskVFji7HkY/7cDL6VHgUMolqFAg
2XKZ8ZhyOJ/dHHpYvFZpHzQ0XnzQ2/FyHI2KzNZaZouJDICFAYSwTxRzOQ+mA1MyN7mXpTzsCcLu
adDaAnhFWjURJfKJ0ujSu3ZU+0hwa7MGMBlMeV65F5eRS1L7BYfEmQW6VJKyAtiggCbyrEmOpO3z
4zvACkpZ+VXBMKF07bWRRKn515f1XBCNkWsE24M3ZsEsOE4aW6ZA9wBvMfSSlA8lwGwvnPvn6VWL
1Nul2PKWoEJb8AnJxn7rOXAbqcVOCFTowqVuqWuG9O789ufJl/YB4j4SZxvHcBA2/QKQ9nKRCHR+
hVWEg/zcxAm2XNzaojxn75OE7qByW7f3GgxT8evNGRImtXJQXfSu+IkFCBWVgm5IwDA7KfKSMeDQ
J0Wl7o6nx1X04Oa1laX5mcF7bPw9xkcT7XV3WqQWkN+KsHXOjvL572OPSH6NEyXrxu+nByHGDNj0
vV+qU/wE5kLxwuT5l9Y1kAoKEfS7vbIG+9mlZmeGNvMqVs0XlWKN2j6omRuTIzUS8HXRbGTJb97Y
VynAZjhMm9RD7YkHhwISceaKkcSVTUcm7kGqLqt25qFCrcQDExXddwhBQ7su9oRvgvlxJ2b+6RM4
oc7SZ6Zl/kOY37cpY7qhpFTCVJg0FYy9byvMxt9jHp6GoQ+h3zZXoM00xerrUwHpL5xbRbUs+EUq
1qt9glpdbGPYtPSMygtHlN6+rjHxmyZIKeBf5HsYKOFDYgouX9ARlkj4oJ6LTomVbf0cTQe8u82s
l5j2W8aydPve/9CWrb+VLhnxqz+8BJhTBvvuggZZkoUNUok8EWFgDl9vdxwHuccLRlMYRAtBsRUQ
TG0owSSLWHfrdzvYgfCru4/R6Rga0I1XyBetCZeCsCprDGM6hCrSL74CzEcAjYKrWetALc96+T/T
Xqa4MktWQJwiJzp1sZwRze6L/kp+atb4TBcpgk6AqVhgEs02G4WvF0YsnYG8pKezm7i69R4466Wr
i5ptoyfmC7QTgdjvQ1DHREPtylaKQ+2Gf4xw+07NQZs/sfEBGg6vkT0KbTUHkASDQTlWZwZjYUC5
Nd+cKsdoCrLq/9sZDUai9PFSkNySP8Bo3MJsK+4VYKPPwMgNmXsO2FHmRfaD49jR0iKckxldEMI5
W642uUgEKXAUWYpjD3NsOYNx/6IIzkcrHcz+RityRkNxnfb+ia+J04qmOI2qYRJuLL9lnr1L/IG8
asLGVa4xvSjSNyw/pvQILW4IWKdpBF+KvuwAh4TdqkPXTJkxcIXZ/OZLxoWhghyrSLwP/FHwAMJV
jiHoauhKfIrL+bTz4sgEbIWlfbJXOZDFMCLJGJs/kRHbF24SudY2zuFtf232bRxO1N1SIniItD7w
xZO5W6iB4MwOj1Z0/ozT7macs/vSvTAWeypJS5FjZJDRMLzenK3THP24N+cMhuQcsHS/YfzcCer3
uq4K2Btns6HLzo4XMa+L5tcxOIZSThP4QRxK2mAfSWaKv8ebzkN7zAAmJPSwWJUCtRAssCXZ4VRY
u79PytPD9/NH6NNf/28zktH2Rw4xY/bIknLr3zSJJ/7YlMYnqbaMy7Zbg7dy0ggJVjPzXRq20cej
Rc1VArT83I3PpY0/ncBWpYmpT6VCAkVJBy6scwHnH/oDEHg7NGJqgh/s0wyRSYzVCKNea4IVpak6
kq5alLnuBbfkbcZE0QiQjEiRyzMGf4ZAZucRstrSXmW+TpuTj9gA0b2ULSTsAsDo1xB9qMi7oZi/
GRRRIZ3fhspS7GhFYKKf9pgz5aCMVFVZQPy7XuMOYB0KpVyz+J5etbfJcLziDoY/mpkp6PDjL9Hj
NQPd86PYCgcYZbwy9GRd7bqXGwYKfT4mnXgxj9A8QRjKYYZcngIx7WwPVQ6EhMfpVqPZchPff5Xd
3zivszHMc79EfCjJ0fr3fIzLNDOQn1ntHhG+hBdHLoJKECRLLMl9iVv0jD7a2C3T/6y82jUeC2Df
VpN8UQZ40m0f51yhlkassa/R5HBum2NY/YD8AtnUeiPiytSQKOOYC/iwYFyvm92g1G+kosR2P2BA
eqSUgw9IzGl58bcNi6xnk/2oX4kTswlxzSu/xjYSmAtB67OgiyDNBS0bvQ2kgjW57jCi8ttinW8E
olGTDm2FS5RSMoDeyqBowDXrfy42wv+Oql8PBuAOkvxa6hp/GviY9vd1+uBtVrksjpWlyhQBSORT
Wkbo0AMutW5JnqSzCtwCBKD+axgfmhiwsbB9Wu8+3WEPtIsJdVsdrh1x5fIS/hujeb1K6jjs9f/8
6+CO45/FWzDGKZ6TGNRyRqxThdZuw28oWqW0w6wSadDF95rrUw1h3+8vC/8sUkJ+MRY3wandNeuO
I7vofxvf+lY94VEWPg+Spj8nPCtV5abq10YzKCZjHEvgp3ad5i8e9PFvY+ojPTtgSkfLCSgE4BxM
IM+PvX5u3aGPrJSxJGlPckOI5d8unDfvayB/Zoj3HDbLKVyUL1/BtQbpac7aoIfDXSB1hZGMWsxq
qmjZZG8JcL0oQnVit89sRchfKc+96sJhFrLldWdyO1LAKsznRhregML942Y9WiRO3WsziaFFg+bX
280GonjoqjbZCqKdARdvjPzxkL4hz+IC87l8qi9JHXo/LFEGMm2bK8sxshVjxArAYAz+PTRZPuD+
z12LOr7yVz22Q9meb9/cehXb0amW0t8Nhw8y9ZoQVaChqZH6FblV3tePZX2UyphEDGyPoziNJ/NI
ALOuYnYsEt1HNBIHFHr9DTo6SMTTcTYAChFRx5BeUkACPegeeJVHuL8iv4wsvk6ymx9PwmUC9BCG
YOLiq5TQuRJ4LsX3yCPmA8dBy1RmzPEuz4cludoUV0x0aV23IfitosIoWT3N/wg4BAhYznu+huqA
tnSfRP9d1RmnYdV71n2zjX7KJCR+oAtyS6cXOlJEYG7pa07Ap5cLoe6jrI+mjTLyZ44V1zUfegRf
NJ6fvaxdJ8Opq0ITGT71dYDa6hFLIAMSTCZWSmReUD2giw80dwkQ7agZ0Ge+1kWAMFP/yFxaHJ1g
q719AV9FPbdmv6X7yhIXqDVfN+vamXzmhW7OYS/hGjHloSro1t5DnmS5v7KcR/Btpzuu7hnOwt6x
MEE4f0c67z1kkmVTBEMSYTX2l2v/E3kXcqwDZVj+CePvcYgSlT10hQBTFKDZRmwsliGDl5En/7vu
XBEB/77bXSBjnTDSBwScHi6LvY5yd/aXDXnF4ItkYun6FbypVBdBvJBCDzl74ImBDSLJRc6s4rzB
AYrqDbnEFxHRCwyCVJdmb4IbCHs7CQGQcY0jK6BrcMwGYVKW+36Uh4tXyPJxHXNCsiFZ3B96TG0Y
g2O2x1LfPC3/YkXzs7Gwov83cvrXvP6qN7fbiWMTTUeCgIwTFPSlNKYEr0XrnHPKygOt2LVR4HYi
GgSTJpoFSref5E4vuk4V92iP8s3hIHYV/HSjDtzhYpCAvtni992Ua9yU3pFtlKjYtQYnszSz+5Jn
eMByn24FXVPmG0PLftj0y5lsESJU4+QFzS4whHR9zbyFvWaTselM0Y9RH7D1sYODEnGTB1KHOT0G
ZJMhtNkwnyVtjpVVq7uhcofHafJMX+zg/rUyrvaevyw7amWEsDJfj5pbu3RQqqlp4Vwmnn5AZbMh
pX+OMx871tuuCJbfVDzs8zZ5Nyjl9k6tbqDJ1ZkbVhXJf3hqeT46cSkd78mwSMPCgmGZKiU/E2CS
Qwfc9w5Ec+itW0D9Xq8lEk9ajURgMqqPZNxFeGzn7OjoX9jSibGelxI0M+SV4AHjlt8iXGQZMCMz
lOYjJPAsTXE2UKwWG7nldD6a8uMeuAfv+ZmvHPBkPO6q5A1ha8PCBr1Y1KgysFP4O9s87SQjS/wK
jx3J3WP8k2MbASIMJDEG3Ql2wZytXLNxjbpWse0hdVKmzeoKdyUMjqzg8OLdVmWjIoPPQR4VkFbd
kZ16Gspx1d1nbK1RGkKsag1m8uyZzwEzory8U4r+gB01mg3B/vMA8RN7MhPpTSEQ/y9uGn9CeCfC
LWtdFTSho8mV6JmX4jcHxwj4fbxVl6P0nsjc5WVAAK1vjkPr9MlJWz5TsARJwBLmWvg5gfaf465e
vcIkwaeoOLYnlbYWJONJnMRwkYtHXi8Ool3qeZgSihy7/mcC/0f96JyykynANcv587uWawEdN90S
5j3PCKQ7yw47qt0vhWeAK+34b9zRJvz7EY7p9Iot3v2anj0OksNvw+UOSGWpjAtyTSZei0z4a40R
hI72WLspa1DEU9YlDJsNKbIpm7wk2Atr946XAroMA4DKLPfdjBVD9FpGONxCNJ/FQKxqDnNAPf4p
GAJ7Zy46SY0nkv7vx3qQed94WKr81PuyKYKX9cLJTi0OJ2P01ca8k/azuYwmgTM70oIxLdgqdsy6
dqsNBmk3PjpAKvw6O1oIoRycm4Cb8YTLP8YM5KjdEwVSfhuSzMHs5UHZo93NwdZz6idmwZYDZQBh
5Mk9V9yn72bl+S9X6q9/dddpSRSbBph6Pgd7GgsoOrQFL/o0IRY/vaDFIiR/YOl9izPlZ1JAPQLd
vVG76tnVRhahlYAgQ0q712j3fNpbTFT2QDWq1+ribO87A0lGeqiOQS9zaMYDLD60EJri8f5Cb3ko
G5FcQboOD8io65Pe18TonZMNjrPfWRbKtpx4SYeC9F+zbQFWu8nkIRTdkCwVLb0FcaRBx5WarFKk
iDvz5QtuHm7GtqxOhJFglTD5pUV+Utpm2f9HsV5LhhMWZOelwh7Inkr0B/D06nUw6uxT7w5RDWKX
mNXV4UasPSYEeqCLDvovltAH/TTeqlAV1SLCYeOH5mF+2jP5t5SF28VAcbtIXv+lKHIVXWuRw5IR
5vBja0FMRoxQlO29Il6q0orVBAOzTmUjj6ehy9LTSHwdUeJ+R+chlur019uQ1NOv9ZZhkavRxUiU
GKpLi8kX4K4A8lR0C2+YKAi2mVcCEkfCLU139JZ4D9Lstnpv8ZqRUilWrXr/y6LTdKbD47RYbg1o
vfBYL4CSi/Tt90RcO2/H7LiR967dfzt7EYVxIFDPnB/VUy3riZbpPxmZrus2seBpb4S2ordMi/Dd
qhmrvJ+ZqHTycedt0Z1ADxG6xxm9KEVHoPPXkirCAvx3DsDVVAU1NWVjS4N9Qz4IdAzWr+y11fC4
+koo11LSWAXweXBZG+RMdWQSTzHGCcI+PMpc2HossQD95AlZ9eQ2WHuI+mbD4lxF6hyXTEHeN3zq
PS6PcK194Cru/scoslAheGJy5/tLkxpoz8PTKKKRx5VSy3iWL5SbL60X2/sIQ4dSrbpR1RB9uDxx
bcNYvfi8biAWbpeQYO9njWM2fdBTVnyFlFMctcHXVbZoKMlEYMgOY46Hc22dpne85wQ87UftkYkm
vnWlYGJro0a1tNX+Ll58s02gO2hEywSto3IP+z/AUKwE1CAGsnH8S64fQB3y9sGKXgtR3ypxiL4Y
trFMKL54hH74iXBo/btXYimiPfMS9fOqRY8u3k1YcpPM6/dJTjh62QGHV6nzPBd+YOiM0RNmDb6J
1A0aub1/hrm4DkxpdmS6WUxVZfpeFQknaU/rblSuittkSD4pEC7HaEhVi35ISsN+uewraJO7k8S+
o2vEXSQNLq2RkCx2siLliMAJC1G5g8JhPK+UA993yp24XcZOVG/OtvxR1PO40To6uQpWMOWyX5O/
AX9ssIGQSrE+hcepOuGLJ5ClVfxsOeVZXQIjIk0/YuxUw1C1+dVVN+h8NyIoiQtcZULa00VXfjPC
XBztyd7x5d+UXaCPBecu89X1sqWmERNMElg8Vp19yh5deYaXO8Z2doawx3hJpStQlDjYaUh5FVbQ
iv1EE+YVNi6+PqcjAMr+5POgJLfqeYLXmUH1rIxSbDw4h66sTN9pUeBNHYuFHhcu3TBAv6VCytJE
yhZqjODOsIsVev+SE+iiGParVg0trJLKEXjf88YxhsrjtBW1IfWsrLGIy+5BemM8DaOgdYKyVVe/
k4AdG/HF6NA92MVitaK/AtZOg9Gac4k+slr8boPudoAJ2opSt/mQYEEtVsJvDS9wnsehIHTyVjGA
9lJGwrLlKbYqKUk4CkdvSbI73aeSmpCqWPtNT9vS1Vf0MtQjZv7RZttSHKxb9dZ60Clx1tVoc+4m
hW5pZn17TujfIvPI9YQWAOf3fejAxN6/ACTzB8oMhDtcsEtG2AQjfa7elvq8HmLB2BkLgakzU9aE
sJz8XrrkqDB2AtdyABJ9N029XCchuQZuVbH+mJDfyWQhu5/IKK5QXQUY8OF4NXpUZ43vqD+WkNOg
av+y+JoBu6jcw/AB2FKS2fn/ldhLwnlL522nGR7GHtADKedCF86flnGb5kew0cW5KomEswYelFfu
0CW92p2tIb9rCROcvKdTucGEl4K4vNvtTlqxekHhgHJ3Hk5BvRre2lYTjNj6fIH+T2+KDJ2AEAuj
3aIHxOLOAuKWfhak2AUAdPAkslK++o5CxituBaJTHCeJf4uVrtAQNyytqqrwp1N4A6J23aLbOlAH
FdykNh8Hyg7OXDR6Bqa89XBIdP5UgnD2bZeiMzYGvdW3GaDce+0ZUFbaeTe9qOa7Wp5rUL+vVXgM
eVQCRsQtDKrqeOpyzdRKbgaZZS09EbrufgqhPSb9hH6tmO+iYils9RiGhlxxf7B1xk+O7Nw3/2uc
8kiEc0cDzqxUjbtkQ3xU+sQ2hAiRDPrsREknjyIQLFtyb6S/bR5iPSL/xo/gtNI/+Q5aOOuRQneq
vIOjZiLqsjfm4DzNh6VdCFV2JW9kxe9YSKcjzTkkyIBC4jhyXQ8+iGeDyxltI9MfUE61hf5wSab5
t/XYH1xta2thGsUalh1JYHzRdJT7c0t4MfQPcprgECAT22a/Aob619sl0VySYeFGkLAeOVVpLJzr
/CYi6s6hAKrqoEG5D3B2dmmlkOjKNKjih8knSB4UaY6waKoupTbkkAQJ+lc/CYC1FZP7SO3sb3BT
5wW+VhGURzxuaUxGrb7eC3UGM406VSQq9XTclu7uF2+KsGvnCOLER+oy0dYypYbmbMOUZ/3CX1Q4
rBngO8BqxA1Lk2dDnBxNNyOxyLfzjitYKc6XFL+xzfS+l7kMfRn2CLUv39xTV1m6Cp2Tqa2bxrgw
W5LltHGOvSVaX8jay03hTgpIX41gRkI6KF29v4UAmSIfCSxHABp4to9de5qirSRI+KDC48ykBcV0
dRT7bYlOWXOj7GyQe7QA5b9h5kqWUBv3xOw0Z37JV/lwEft7KTMLPMVkKd0FnGueAkHnRUxklK8D
eZwOI3fZExoY/mAl+SvNV3631L15BxB+w/frv99s5fruoqNc0BzVixknwn2Rbnb5gV+mET7I5gL7
IbAg/Z0ULU/58ZqZzKbi0AuX4vS0yPUujGNQbRlvvpf1okydK83fZtv5yo8s/w7WfsafhGVAouRG
inAd3g4hK8eEZdhqdPBxVxgGxpRJGfkdmgRtqL+ki42Q2DqBX78H/kC/MSp/3Jkf4L8tGpEVlMpg
0m7A6EthGtA5flSlBQgZo4yuipChJwpbNr3g6WZaYkPXrxOqH4mTEK0ojPZdf6CL46OK4vLsjRk8
CHfn1NeVdGSkrIlweTOMzGqHu7AYa6jBi4Wzb0/7ojpmABZaDySNMeHsZBJSB3LJ5BtpxioFj6TR
3fsv99RWfLVpwbp+WJttiwTqi3PP+/oCwhOojiUNaNUnEnQuInGYYthiQ5wKwJg00uNNKNkjzsVY
E9vfaP01WH731ykrirAKCLYfZE42tH3NBRCVXr5D6lUcJU1k0+PcLz3H1Lai9CKy+aJpVTaqUwlv
LYeuKlHeZ5NBSE1L5foDh2RvPITPkK7Hc+7R/C5A9YJLKretSJ/sNVohpWsUwbqpkB4+JfwHJQ8w
ca3l2Zw5E0iA+aabU2Ad9KfQjW4lUYE99QlinekyOjBh8R1SU+kpyhPD6fGYuZz8SOXyZBS0zIY5
f76hGbIrAd5MUCNHPiHiBEqodUyIjdgbE2sd2G32C/rUeI7dCG9BowGoodKNB/RUvsx2lohfTy3E
zT8zc9R227ejjwMQlhUNgLlPK5r+TxicrVjA++RnvMWMDB/mCN3Eyn7leTBd+udPRvQcfPDXdxkI
XKZ7hfv9HQcAIAEqRrui6dB4n4X27uboV9bLYcu4L+7q9oojlO/2yR4VPeYcsBllM4Apbk9fhYiP
tsDSnJ3fXpmIl5LxSig5owkdV3H8Rp0BvT5/WfiDXBHRBWLrbLvNBc7zI8scM3Ujg+i9lvtUYzqQ
LN3oNfD+7Ff3dyCi0MTqGPKYbr0/ZoDPd+HYFss8uO20+mKmI4ofT5z+igzbt6YjYwkSmlXfSVio
Apf41KxGMIm8cPTNrQhf+yfudYdmLJStj95y7dAH5s7zCu387fg4O3pSnhF5str1W3+yyOcdu3Kp
HoXurdS0CHx32B3laFsIjt328UbhEiSfl1VvDpBtq6iik6OAPRGb3aLt6b8YX4cNRd1nNBl8mc9Q
kg2GMQEbQ8v1JOs1PW/fJ8VKc97lDiYrMxQTuR+hGT+MxtZYowqWIzo8g+GUGU3/oq/kY9Dn0pIB
FfeJlduN8MIEeWjYfOfzlenaQ+LosCRlpXPf0gteR7NKYHUdIHSr4olg7c+ZbwnnPLCFjnLlXGcn
UVAwM/JLtW6rVNkEuyu9dI6/tABRv2My7fmJNRxOnqaxSEbV6cPVrxLK3ZbjTuZYVi5tv/t/8dBf
NTqlGeQxw4AXGwJrmeY//O+8yv/efSr2W+sGJXncFgNNt3gDtCz7jkIXkk2pj15A5fzX/bRFYptA
nkbUky/fCnB+xrh3VWxHNNy5GOn9VQ36xzbSXi52S5EmzkyvbIgA7GXcH+mCZomYN4YpGT8Pv3Bv
ZQ1kQPKUbLlN2XDmvCz99F4Mfc1BoTHrnBdc8vwanIzA6mhO9SZ2EUmzBdw2yAf71ofX5AOa1BQR
WMErK9wLsc0cjjnrOeHk03TG0TgDxXcmUzokg/+gQ2QTzNwp5gyLOIuoV+GrviLvqFYUjVLNGyuH
qMgEUY6C1s1ZFQ/MFEtmitb83ItnMkaRCRzgbxf3JHIgP4foI2FkNjlVEw4a2Bfq545sQxHgAwDQ
26GGuZ1qJPgO4RZtbML1wzWOdf9jZ0506lao+ejRxRUNH8dUvLECtiiRkJvGEpaWEV2SLQBw4Nbj
tYQTK+Tb9/L62invZOBKj/SniUDDokWaEl3Aa4igsSBRi5uyPBJnuGtlQnvpOQdHZvJfkvgJqq/G
ap/6StAldT0gghpLL2lRcPXmDo6GE/nc0B6roSUb2OTmra7yB/cpGCCaofgiePpNzJm5kRb7d0bq
WGNaMMbzvq6fEar6/NlqupoZmoZ+ieS9fnpGG1NKmzyFYEHoic5BxeHFEZGEpLX10NTG+ikpTrCo
4IFBBy5/zugbgZBkWrhCmyq+B9te0He8jSLdYHe1JxRqbuVW3ViBQ++gYyZ4Y60yKkJHF5/FBXPb
Ncq3CmSKFLfUhcfzvPxZNPmR/wE4nDuAoa93AAk9pjRwANZjrgLGL1K3G5wBRDi9rVjuvumoVzKE
eI7q5+EjmhJnkYqsSHv3WuVnV6tzsZnRQZIGeA8UyLrSw+OFvhBqP1CdU0PkOLbvwgxucHb5JUk+
r2HbpZsEvzTzrNgSXGoHTHr6g7qgZghMRHJf7vGgHfY6d2AgBFeGwkXezo6/JvnD+m9QTkHsLq4m
PURdM57m2Sx4nW9C7o1WJIEFVVleFb6HfKGy3jKrFnN9tQ2G/G5nBxMnMHhulAmoiLgWrF8Wp0yc
ZVyLcXRSsqkiU5Ic2JNwz0i59WU+bkmDjp7hwlafyqToD2QDeUYscC1/4FcwiOoLI6VcRuWvg8rI
+xct5JASGCxxrt3S0Z+735VRskGHVviq2H4VrMVNbxwlwHukpCtmVA6Ms6ipHXbRGebyVWdReIsp
uE3Sbbi3cuqQxqI/0+tp9X1JG2Pe8JNIkq8JvH5XDut0t3QM+N+Xq6hBE+SWZA3knXG4srt+FwAr
wqexht3a/Oi9mib4yDggOnu0JVCsVyTDI5zF96CBptpJsxPW0sb7fLG/GEC+TrRzHVquEY86xPaP
Ky3w9ERmRBca08MNVxlFg79ih444zAbDC0gXj8bufJM3ZlihtDRF2RmX81CgOswcij4u2QyQKqY4
am9yhiSvJI6lIjT+I+O2ZbzEvDafrfiE7FIoGcV9Se/rlGrqOU+mW0WTXfwOgWjKpG68u6fqoba4
weJv8MapyVUZidPcmKDf+gjEL2vamLzDo8uNFLEZrdWWNlV/DZvmxq+l+uLGU2dya6H9biz9HBRe
4Hee2KBgwWJPxSF0IBbeW6AsRG5LxAQoreSmn4G0kPrOpYITalLRrbRN7lxpW1+YEKo9xp71FPhs
V6UfsgRvU12gGw2aIUuOK1A+q3+7UPz9NRa9hlOcbgKx/mOe1TuKvYzOqXz3WY0ARBUIGBWrC3A9
G9XoNfwVyKYBYOGpQzVn/n8/rUATaKaSsdV8x48CUgxRL3Tg2oeF5KXtld64KFH5uOwcqDj23nD8
ewjmX5z9HuZfGOKVj7mYyT7BfmomKxlciSjRovRNgzLT53AsScbbVC/tG+zNese/98BwJv/UFWSQ
61CCv/RPJHKILgagQBW9WFbZhxsJTmhAKgY4ub+XAuLgPSi/p79rogL9NAgyMr6jLyCw8p0M5DS3
GmgzMPVcExC6nGA9lXctkNSQCLP4y5Ug/h30TwbA/LePFNYGisD/6CjPJe/mz4z6L8+Lx1TYtKHu
QCFkNNWfxOUu1vZMGQvZt/M23JvqJEDphzB0WW08rnLDP9EnVebTGz99bYLCs/5wEStCgPv05pbu
DP8v9GWb+EUqghPa6BUqEDlGX2IlhODe1oE+Jkn+oa7ie2Uwr0vQAtUUZrHkQDq3j2cHGuuy8LD+
x1gL6JXyhXrQxEAuVM7fBKVaSAULYvGHi5UxJYO8E2imBGO4KAJpKf87sIc0hSqBdp+6zOX4Jfm0
9UkB4URoyijXypjSPxTsWwZxlxtvCGjsdY5Z5uYkxB+E3/cASV3609zZk/F+kBeiz9jvZx2yG/Xb
8W6bOEnyfUuBFS2bQJM3jdPVQ8+3EplnP0IELHoBcJ0OyTRaTmOnicCL+ukrtypHB1YBjDRbA/hW
6RfbHJZqWIjjKkEJi9uYXGBQ8c9ftwKBO0SHD6z8752vTuPBi2jWhLP3IJ7ivs5iawQzNn49duVb
YWBUwzRQMzmAfiAsArXR3ybC04/m4I3YYa5YztdNwsjdX8F+zACtgQH2ZSF310o8NkxLmXNXifcQ
dApHbvm0mxg3TvSj8/WdqeOhOWn31aOzn8dXkAvofVTcoGSOHkKH9R2j37EXM4NQn0eBruOCfXKi
7+omt4PDdarHSRQgUS7pWJIZ1i4JtL+hcIRoH+oIsa90rSXNulLkMmSFc1JmHXhEVEMUwQZZpwBC
JlyR/uZmTs7FyAj5d/vCm4osGylg9Jrb78D0YzwsczowmATuDiZI+oWRJxHFCVECXEicgamYCi3f
2ZQnfVdzhpesULrQ7k74cnrVMS84agVWQkhTm5qEzetzHI6TghuSkRF3WKQPRizZdbpr9VUUSkCv
YFxtkWK6QUEk6h+ExYgQxYeQjQTVt8TtUaam2X+hslnJYE0b6iBA4QP7ZWjaMVgv84SSMP8aRReG
d+ca855sOPjXf/wI1OpkYJq/K+Gv0zHTQtcawwiiOC+ads2aNYqBGiIFKz+OUFvWESHfuU5IqxnN
Ypnlp/JeIz5wkPsStS25oWGpi6CiCHoJ+6QGiV7NSAZ7SgyHZ6hhVEUbxi81+cdY6x6WBwPFT1v0
I7b0aebkxqM+4CinWJApM8dHqd9OveD8pFw69ptg33rTgIWmmiNqTIPhtRngefXeguC8cfNCDpFs
i47uM2Rw5ngOde6IjdaIAoBqIBpDbofpmkRG1W1qxfQczB6NW+zj5rHOPYjUFJVZKojHLAdGiI2y
PiLDCc37wPSy7dVmegU1ge1t+Egwa1jrNeUh+fhWgWfG7p9pRLl6NoOjDiO3ZJ9CDmUf93lxpSeY
yeD74Q87bS3bzrG33Np0VhBfkeRQErYeo09i4G61qYj1lWtuEvOrjAyvCA7+ATmm9UPeoVAlOX11
Avh4WQsDMxCtivDsL81mRmTCAOZHXuI3Xpr/GsHtFVJ1+CUBarpkQzST9lzwF42R7dTzOhk86wOG
DC84ALDF99UXS5ejDfFWNdwHZ4wvYYoD5B5JSWZqtQ+CHWpmWrpPNdvgSHTsmN8ZAKhmn+xazBP1
NgrZ6C9hI/3oCzfqZuih7d5DYNo+9q/+IvPFNv51u5Vzco0oeXOUjmbLY+aKMiZf6IsK8TOavdfZ
9C4odqtOss7T0LgGXXarPcVruynE3/IV0FE2yww8YryYg+JXWxJwF1EfzKd+x5SRM9G/48JSpNil
Jpr8oKqcdBSJ5fK0qhaBDhhiPLF/2AgOOMyGhE6jvyPq51WF4+CGpmXUL4UOujAxLLjoR8yI36uk
6OoJIfDfvG+/R8DzFCk0tWCDH+5OTfBUwiyqfQ+/nc7JpQ5NyayF6eJbprvOGNVqZeySgkg1UurV
rmYN0ElalnZHu6Iq7XbjWwXyMYwgMF30ngoo4MWrczSl+hm4bNCLjerMNtnW2dGFC9gyrXINLIU2
x70oA4lXS5yyRwJrPYaohRoFL/yM1sak3qHR3tJT8D+2iNYQ0c34a3/K+JZTz6urO1gQtQnDZs+W
CJOS3PK9JMv7hENpn+sA+5vhBkwpMUzOKff9jEUCKSCuqJak1ROquiU1teTNrDGwlMeoq4JVohuR
JD5YYXJkRynjFs2xVTj3lYN8m0kuu61hk4ZMBCbtcOLgkt8VNBQFekzJN5u6UpT6uRYrczyOwpHo
pbK7t/PrREn0c78ABgctO/86NHKD/hEphEwRp+G7u2Wb9Gwfj4gQXR6Jank2cDyuKh6ynvpN5puR
stZ7YqOxoZNOyPzS4XL/orFoOcKdIq3XHBlBkJeVal2VKWwJg+McaxUVnAP966cpz7reviim6y6h
nUjPdCGNRI2hTbutbO6lxdS8q29229UQ+jfnIBJ8IWv2/XtX4Dl1wfw2XQ/T4ekBYZqc73PChE13
1XtK9QVw2/8TuJOA4Wy7qSrbpk28HjlZF7uTkN1Ek8X7zbT77N/m0AKkRXriLmfpPFMMureGNjhw
ddYtlWwUZBP6M4qAzEv6O81vmVEm/oUfZu0/hHTzS+gdKS4NoHXqhL6iafcnQ7OJsxWbWPkLJYCe
WAkjWyOomrYrSLV4uiHXmCPK2vmgDW/sRqln1a8F1xRqEWBRfaZWbr3F8qLlCjv3ANUNF1Q75MHf
aq6wjAQpXDYwFPfJRd1BFcvsowt4cSqXW07imfcfdTepZFdbGXHeVO3XMPv6pBrK/3yewfqx6cax
GRiLpfAGS2NAll0797nnCTx/t+11DtQoQnAkZPfaRuP9OY6MA7tUWCZ6nPIY51b7fxMlYH3LZKT6
VOgyVCmoBqKWfz7ypw1QX+Y1mP/X+37gyFjDu3kjJpiu4oggq6i7XH9FVWceBJAoe9CP20fIeCIJ
+oNV25yrlJQ5AOZ9sqECYrTP++HLdpQMQSZOY1LGiOEyanxBMkRc77z/oq3k/3LRvDkUCjd0zI+A
xmZqbwrfb2or3PGTJ8mEKPT9VZG2+dyPWtofyIj2dErROlrjlL33VoVjzM2npXrIyle3N7Nko4YQ
yOETJEjvhZNj5LvKUshdK8ujVC4bckjehO7rhfkZrkyZA68nqpS7qpQj90sb+79h6WBtlrgQoQpY
nBUojr/jk98LMaxAJHF2j6RQXgYV1E8O4S7yrAGNzFgf97xEZtMwHWeGcPtTMx5wYXpPCMN3R5JO
9MzZv/UKBz3bWVaPpKd9u4GpcxBE89nVtZ7YO4MA8RHyeVN8JmvGTyPY9iNTaTarzPL3hKIzO5xx
OOIXyC8j3ESZMKOG8BqJNHbFUE6bWuEy5j3Kbtnu9fEzAXLRaWKPsOqO4U7q+xWOZNaJnzkDpF54
HuVqM34IfdMfAXFRSroYZM01aEbH9D+UCBNZ6d8s2+3d8ORyh4bwqFy9Ypw/P+3oMFF40/U3JQmj
B6tMpns6e98gNwJQuvpjFN58hiIHuTUVirJ4C4zVLL/JuZKgiHiNFkgMcVYtJkZlPRwOgOvTbf0Y
ymyhMsoTulIVCO9Km5oBxhC+UsKkoGyGFFEUTh3xb47OBECjIQh8tZYqYSOvYnqmpK9Xqo5IG4CM
J3S4vwhdWPdXUs1JlEAqf87AT0w/dcok9yYwaie7yAH7szW8nVimxov86MXNr5ZGYNMa7bTqcFHN
5FxSjdTg+18ZQz4xfVSHdjJqxNitkjtmphCg+ffrrv8L2Ll+xoqm+Yeu5Qc9A9r/xFtG3LYnAsFi
9dwwIW3oLl9GTAQFMSKgG0ELaNdisUmfH4II+wYRdeW4KNfqG6v5kvbDX//uTXFSfmia/y21ylWA
MeDNEIwxrbIMruE8jpLZxzGh6VzXwfwNfpYALBR2kiYBa/VQrbm3z9YUoisWqgfHVuFqb17Me/CB
p6DF70wI4kO37XC1nN/cHhIlIFYvZfPiedL9YCl694l8jdd5nTU7JBK1uHXIZ1iiY6m0HqhuW4Sd
0vyr635Lj8dhUOzoLnQjWg+bj/tsUWgTFC81NhA1OQjC1inKy1Vfu6skv0n2w5/kp0xMCP0nVvnz
JHk14u2oLqnv9CPuL8DUswyCpa2CfyRxob7xRrEj05LfcPyU7CbMrjtiaoLR4OhyPiPD7BRzH8I1
q1rA7bsxCcUt3stFnswGY0EWqtktJvepXXTlvLNkm0YM1Zz7rJPNMsBVsJ0IZNmDwuOVGfWPXt7r
gi717svHe8g0QLM4sAoFSB1ijGi/MTQU4POPvFCD1aq5GlFLfYhB6etwc/KmZY2bCh+8Q9XMIHbA
5bBMTtOgmNXQ5A2Kgal0fm/we8f89LKsK9PD0euTHWN15LuvQHVKy4P0XGMifV5iw64xKqUnbOGP
H3tzDLj4nraBTPMoxL7ozqY1AgTxTpdF7lsrUMd3nRsrx6kfQz31fAd8wZOK6gmJWwaZg4Bu7YUH
AIwz+mESAOlPSVUhzM+FkSE1VG+oKIIAAT7NOMR5HcWJGeYZwU/ilOmHvNWg7wqHYZ9JUnUU29SE
oD9LMEQfAG/LJPi3qdLtQYyCdyuhrQdW8mslThx8t/SI9IT1hjuIsSgUp9tcBeZ03TzMOD8r7L4a
CZ35NyVnRSsvo8ias4ydKc1KOIVIokKRCHTp23m2TEU7TXALLT2WcBV9IuZIQcdMjNBumsroWfKl
AChPiYgn0vwc2kXvIckvG4ogZbJb+1zdMO/HvjeANP/V31Y0YSSnlz/+qjJkHXQcw19VJAWJ+JrS
98RAIGiYyHLhEVSReYi8qYyw1hgH/MVr3uram1OCP6sCrqvQ3c5ZfF2uKz6rGeyYzuMfb7UX7548
UmxY+Y7ipKiIyUhEWvK9WFCzEcpfID1i7GQbTHIPgFwvifiAD9er3UgDEw27N6eT6WijM9TSGXb/
EuplVVWF+sMOIbkouKXyshURtZ7CNtTk7u7v6PwnyaDuYavVd06XTWuFrrENK9OBV0kjGZrGAT/w
K4/tj7W12XJQF6ixayAVV8B8KyHfH+yiZz6kpyRq3IRFFGlIEiOVeARAURkRO2TI3VgBk7imKV95
4rRnBRZql7m1C5eO7XMwhTCLtEoRfm5q8mrFTm9nU/O7daMgkFm0DHkRBHSuZjHJhBAZtKZWx0wp
guUERu1o8agqXC/e5yrFdlOhBFgqJogWBdmVA1YEuyZbYQAKaP2nOxnpMeqnKi4EUE9J5N0PxaX2
D2EETO40LGHMiEtXGoyWnmM9PRiX6xqQQn8E+om+EwX3W9XrrIA2p32+87bSgajSYAqJcsit0t9T
XXGZYbz7yXc+tnC2yRfF6PoGUEyc5v7Sv+bCPMGYIpffl/S2U2cqe62qopSiPPFieN3SO3K4YySg
09g8YL7FZ1H2PHVL4dLx1zX1McC27Z5JoStp9Xzisv4NaAgW/hqxT8s2Vss/61Tu/ZxWjOUKU6Oi
/rBKjtoHDspcFtEsTm3w6hKSeWVGNT8TSVIJMVtEo99gA0wEy6MwXp6M0NCVCCbdCtMGIZwiSObo
asFbGkQB2j/C5nxOTwESWyArZnOc/pzh+KjAWWThr5vvdq5771XUc8e4Lr1b4BPuG2fSzR8Iu5ue
dZ/6gu+hoekAKzoCRvN7TFfXeCTeAMenbzCubgc1WvBa1g10h6Jitwe2tU3hVySEqghN+WMuMUM6
VWp6X3PvE/dinvoqrhYMZmdrDVgM7BDZyX2pReA4NzOKhFZdt16K7YYlpGTRgva8e+Ey26OZ6Zo9
pNCB/o+NBtC63F3vphpxgo9rRmelYLpEE+XpArWvzhBus73zpoj7oanddxJA8wbCWy3cry7CvIrB
EqG4s3ez4RtLjpyGMVkIhomGjHuzWSRuoPoH3AvPCSZt5bYPhykxv6xPyODFckZiBYClPiQLXXGS
vLM4cikQDdSy0lb4B5W8fzkL7FyCTIMJrgO8THukaUJEU97nZWcjYY9fgjVnusCuAs34eGrdJh6/
2fd6yhiif7kFKHeHDQaMUpQe81kcV1ohBtLfOwJ+ghI0wCNdCu7XjGYy6QHnPWjY6qPC45405kxR
7XGr6Ja9/hQzyTs3t38mLMqlzVH4yRCUqdTrnOvHzMvcD1RcmSxp5z5NOLLwJkTn4MsdCge3v3+N
AzQodxRK9rcMEp7wrmTBRTbJ8Qu5iwQfKdmQT4uKTbALoT+1dHRELOYTnEPwSTC2EjJwZbQo8Baz
XhGrlRuU82J4vF2uD4y73acyZCER3q1Jk3kRxcm0z89Dff3du+v0+wl5v0ZFTLgfN+9NOOqVvWCE
9eSf7FQCMqSJe3Y0QD0JwHdxdHrrVKulWhR4yrRBh+SrubkZVAiByUYLMdhgURsKHFXNghfGaqe8
6J76DiFCMbcT8e01IDONK2MMGMEJP5Z1yUxxgz+FPVaaEQc13E4MfyLq/3t+rdmGJ9WFo7rqj4Wm
RaXJYIIgYbhPKU8nchB+SNSwEkk9040SDJw+mBMlPGAjdiPk7MUtkHBBMN05+7mouNdNIWDfcoYn
ccgKSv09AGsftY116tWE6efR9c6P5StG3xbk1futxY9NgDggFne7i3I/x8TUvvboK2H1ryod5uuf
NjC97F55DaZhhVtxKnlQBJNPjZX9NEBDiyCxhtB4NRNT9AF1/vVlXZmkUTn2IiqcZqIh0LF5NmwU
OHNV8DUN7G7Ntz62GHnDy6TIWxwMCdHfjiS2ULnZRwyZcs/OU7/62DJj14tEqA4oK2uJ0Zmb1+dj
1w4XXTkaelNsS0OHGH998Kk0QQAj5HMWBtP96Cl1SVXiS2HGvOCSJhCqgTv8ZbmWnjcVdS2JAxhj
pxo1AlJbJ3j2ZrZ+Ve+1HeeJ9ttQ6ToJbP6yUW2EwmCYYH/JA/lWq2xGkzvisxDFeNCbfKehwzCA
oQr/YouSBoSW3RgB8u2Ep8JSUUCYfP++SHMW2st1YCXrj1tAhkGxNDZftdRIxRYBuyPtO9wknw6z
O1UWiFErzLXFZT4GUhJzTgnHq1lgNX98s65wl34B52/jyhIbFEFszCBuAqKl+vaHdkuXsBSI0Xle
p58qt3ekxwMhmkMP13/ZYbIDaH38wuzKh1grL5po/WaXt3wwoxEml9l5fbHArr1DjJ0DwHlrHUVV
77HHte4OpoT8Oak0ZOAOC10jOKD6T3yk56Xy2S+Jjn84febaF/CaTFlqjV22OptGNl1eZoql/igH
Jeisjtvd+i71LDI9GrHEIkkneCM92sWog2U3Agpws5tcB8ttK2vY5DKevLi+LDroZrrxi7S7QRgW
fvZQbQlFsO8eUihX0a0ye4qZi+fBhout5sjxqII4rIyW2K6yRaEAde7IuER7o+Y+fnJWI+YpCj7P
fKvUps8scnbKlNOa2HDeVa4WUJEcrAiROGMFpkXZjy169anB+LlXxZVlEmcwzXiQXWQwws8iN/X/
37Eo8v3idfsVH1+VzH+l3m+KhhesRiT/kMg4YDpZNxkg6llsfbNXDSrHoU4EEkO9SZ0aXJJuZte/
81GRz6tRumLFjcYoSJoG5+zOAKXs/cX49UcbhZonBQzUpzDhRrG6G5fyd2llu2Nfp/sPkHJvo3ph
nStKniqjV28O4+PdyHJlHyE4wgM8ZrOQ5p22NC7ho5K3EgYpx6MQUIfhb2tkeXeRaThX0Sl+S3Oo
poLmyUsjQQp+c7cZGym1lZarjp+DqOhibcBrarC0rXaVe1fFkHdt6lo+nWWNwGE5w026jUHFxKmb
XStkk2agD9UyzjyhuHN5Sf/2GyZ9fSHLb0NbgIdvUyIrpPYZ3M4mC5ITSUQdh+gpp52rBtx7zgqG
SiCZ530ViF6fkefjpnxczRhLcpP0+fFf+kB2S8S16QVCkUbSksdQcjOXT65V210gnERuTgRj6LO9
f/t05u5CiK5MGH75IclON5lDBbkam9naa0W/OnW9G3MauTMrsG7N8uqr2jd6oNdsMYUKoXDvoOwt
6/+p/F2ZtuGIaQnDvowA/d7uHPxBXaia0xleTqexad1IHuNgbXXaIVV48+ytF8qAklOrmRhIDwaC
y7y2N7nIFm6V5eYHgoOR7PU3Z99JLOZgcGpFs56Jj6sK9RJ7M0BnHo3DWpz4hm3KJUhiDVJHf870
kSWSASohqqYM7nRlLLe9KKL/0SRxsOjhkXRWqS5923OflQ0KFtyuPj1mSBKbMhR9kptNqy49O8nX
R6+GkIfnbiWCx1oJopnViIXSH3gFPlBDFCjqgdvwHyz/yHJPHViLmV96sCykuKTxGy6INwKMwc81
OFISsjBa2QWS1V+9B4CINU73+K1dLFX3+Aq8150NVkho3f5GJf0sAvcxwJw3zran8/PGt27Fj3vd
aQCFdMxsV9srV2As9SXsgVugmB3gXj8JVjas7Du5/bv2kSxUK11Q6+LJ1bODgXU3fPNgdkZGLxf6
8aIPBzNqtealxCbjEHcFt92wf7+rOk5eHewPehc3QIb//shbql8RNL2bahA5Tj3hsbI2oO/mQ32c
+22Q8aKEkrPax/FVRJMTaQJBd+I4j8tG3Bdq2a/s9HoUC26A/mXhil8r4LggZ0XvfnMF1VOv/IRc
YHpURkqby2N+6IUSBSlRIfOhdzgPfsPSgCG7p3sq6u7uKagk1CquVtgdEbtiJ0/hiN6sjsiCBvNm
VOKtVdPnpj+2YkUeQ7Goza312f8r8HQrIrYHDZwlMtHKA5Be2k+O7nPcsYGK0Ir03yq7UHU46RNe
qAO49KqpJ2Q5lJyiz8L+bvKjqFY1pFPQxAh3IUslToDgPiAi0S44eZH4wIS5MD1UYu/naRZ0fp9z
EHq6iw3K6GxFeMu0ugP8RTfG188MlZ9AZBlsGyE+mwvSkplRHel6bKrAe9i+Ey9QRyt0/zB6kEOF
OITGXo3xtfZGYA5yl4sBt7qBuRGSKEFuQlHXPDLiSdbeZdXuHQR6vIb6muE2M4F3Fj9yYDYZAMD+
RFh2uvLNOc3dQmLeljfAxyG5H0YASG/BRduRImxkPi/gspKhdsMtEXF28APh0RRuSGj0gneZPlju
4fy/+RS5tJ1Ns7rBBeKzLbZi9yFeyfk/jwJSoWDByi/G1m/8RJUEl4/gzu2EHLduON5SMBvnSKFa
d2Msw5Z1wUOtO81+GloCUljYrmzkviG4C/mxdmv7vxG9u/41iGvHMcBE72V9WofRWZcwADzcj0P2
u/9W8nV+4lQOJqBvRAg0pqznWKNUhz4b+4xR0a5m+GslkNaE9n8Q8yXT00ajEfbT12RSrf3hKgoK
FjMal95nP3S4o+/I5naeuTyfngibF+yLuWNUuNMPE8sMdLSSpp+rvPfJ4Z62EtNT8H05xRh/h09U
lUwLKW0z4Nt04xvgKlODnNX+SVI9CVtZNPIITl/1UrCIUhfbXUTJwLrKyXtHJ1JsC4vfnIraJ4cD
a3/MBtELqTndtyGlevoM7Aw07OE9OuVjQ7hRcI00X0M9dEknzoqWXAM7+afyR74uVyCY42IkY9wd
NFwWmLsrYjwiyDEH78GY4bhZnOmqwT1S+rYVknxo98S7+dA/OcsFKMV/eL+O3+Fqt0n2W8JrN4bo
4I6r8dWL6qZWIK9tGsAKe2w/auUYQW5NdrJ6AjeRjE8ZFe160t/E1QfQUU4+HALOU45b8QSHaUoo
DkAuNtyB/8bsxQ90GwklE69qiKyihXQ+GvoxtTDCEZIsP656SlP23pG7DKuBGAX3RED3yoqVKw+D
RdPSGbC8iHXvcxBDp/nZsIlbzqFI8I4jJ0Ylc2i1ZvifTFbc9ZdzWogwUKqU25vhTk4vqDw7VLTp
q9v1P5MQrP+FgIph9YPSEwXwrYflBFiEq24Tc4CZJ+NvmLmXM9/JEaSs9YncDSbxDJ3X+E1BUFsu
u71OjsVbYxZReVTnkW3kS3PQodkem0VdRo/9KY5o19Djne6cihK6oDV6P+1llna3fRjd5wWr8w2T
lIC6JEfVrexfkcS9YSX+vtD5eSQmbFNaFDIlTggKr4NyvepyejdPMJQK0azj9BWr9zSpK+ILJ0IY
b3S+2Jf1etgp/7Jp/u6sR/EpWthdfXP1zHy6wh65IPQte4RxhIUqMNl01TBB7jPVEXi1plde8acN
QPmCkTI1W5sWsUquRrKU9eu2HUZAjSy6Gi298Wk0Ldw++engF2Gg69lXWmZladspK1C9irO+xX/F
f8tWMWvNww3gtv5t3DWGwrzyKHn0ROnKoo6z2sRlDhr2SxmfJsoZySMkJPJ462gl28dkFuRis+Dm
8WibULWryeFvwK67EGK5F4JMjRPi3MwFI5Jo3h9bOZximqoBdPTM4H+LIxjPEDpAwAbRIqwLCy1j
OkqL6s9vdXonbB+1FzsDe3gA7CyN/32fd8piTgFa41ghIOBulqINUsqVjhW5ZaNXvFkSEmtAnW+P
a1LUal0glX/zyR0Vui2lP9OQiDVmd98dkqVYMFT35JKEBWrDoSNCntRJQgJIndyAgoMX7O7hPUvY
mQkG9APbqI4f/EE/CdmFD67BViFck8XAXBJks9g0BgO9cYhcfdYgJ7/7ftoJu3qiyf5ghU0jgqtZ
VI0KhshlF9A71/LW5GUD/D/9chqJHmz0k7svTKQ8h0KrCVN68OJ5rOlA/ovNgKSmef+LpwlsrV2v
FCg3hiB/Ozdm03tsN6QOgLVEuFu1E/Pj9651PAG6ZISgW8E6QGFDTTfAvaEDUjbmMB/iNRBBky8J
1q8d+J9gh56aLeYlPmEGOQhgbicEwWZkYdTiIu86IWSLIATzkdpWBT99eRjpomVQxVy+U2074bzZ
QiuysxQuGP4AQ63sJHiV8HdwtlsnbEPRg7MgD6W3JaS8NnUzunVtdS83vOnoaj7bqw2AcdGnjIjb
3JdKtiDQkbJP4QL6jXBvP8mU2PJJwMYfwnEZv2C1yH2xrmm67cOs6Ie3tE/M1FP5ucneRJ8761tz
KttHW1SV+IndtN1f9REYDJzH3DbZuLu3by9yQLWIbWKnCkfe1D8q5zQzcdRa3gINBlSQckXdB7ma
40iBHLij1JjpOkDWBQLMVki/Rv4sey3DljYqfAtCbEv/FuHu7L/4D7ump2FG8/KM/LcJ8T+n/VVH
5nr93WkCP6ZB/dNbUjbjBwavYJe5JuiNBYioD1Ea0K6dIveG6h4gqxelzXDqf3Qj7DfSsWSi3SjD
EPzOgmmIbWbfh08h/d7XUgpqoWYHrNsciLMfJ9AXCLbGBuG8LGxFzG7isY7/hyyQg7zRwzRL27Rf
FvG4TCkvGzOcUiw5bkbiOVuhX6WNfuHZBCtLjem/2LJpbfLlr6/OY+Uk9e8GdLyhzIvHg3tQMIin
CplmFO+0g9lSuG/0wbW+DxGZGDk4scol4ijxgS/ZIYtmMqpE/GypZNl++i+3sZkr8J1rKZePMu8q
jibuRnA67VAI7A1SCEdQVDFSbfXu3+3xsMyIYBhd37le9GK7+wy7ADOwDaWvD589zoPATQayEK10
esA6ve1LrbumQ6eqosWFVebVV6geh9vRB5+xBETj80egVrO63lNC7Y/L7K58LILT8AYp1XBiVKEY
kSCU9vQwW9Kt0G1CtECR/34okEE/HtwUCcizxpl17oI2RbZapw9EQkJIk79Rl53NON4TlcvA3o6s
M5Za4+NjgccBJ82TPgMRaxLtHZqwF7MLnGyVx39Sy02sBSpAgvg8FslA9sqJncETVa2Pg412fIZA
6dPrpcVP4CfNO531qFWD3oesMKLRu+Q+710peVXdgawrvSd81bC286ghLmhDUQu5E8vmCiiequ55
n3sRugezrBZGY05/PyNQqbw88dlqC0maEK0Pukt+noC9xbx+8XfUBADyzpuF0S8ssKUIjGWubApr
AVSk4igKxyD2qzH8MCI99npad7OUpLjNFejYnB6leWpJYyHuj+1eqOi2/1IOaBmUjcJ2Fkps3pkS
X/D1d4ChDOG5y0oF8Mp2MalB6V0dR4HxX1niRojyHTUfhJI+kBC6hUWMKkIcriU9y+j0/QcGqDPm
Z5d1g3XJAHRMbxgJcPVbIPI3Lm3rKxFU11vW//fJx5Qut+NW75z5bzs3JDxx0RseOGCV63ytN9iy
8tiL0wX4rc8fUr/R/3EBD8qpECFU7BODAf8v21FUUNDvPqCdA+uDWlCH58rvBuTFQRCjh+E/oxTQ
3c5wXqsN5GrzhVXXU8PQ3GlowO6WLFN2/3MrY7BM+X5AWoWbucID3DU7WXY1Bl5nLYItHNkFeui6
rONgpfFGZ4QE3yGA0+2RPXQud6LbB9HVF5LVcRuAgn3FgQ88wpjZm9Hm/Wd4+mQwOe6N507n1t3Y
6qKmFm5CFKng4+WzRPYGPidua5I8P5KQl5Ir9+QFb60iFXSsfD8RB4XKFxPlrTspalRaflvD0vcC
PX03aIYU8HmKv+9afNE53+kUMERYPG6MKxCewXbIhYbeUsA07m/TIH9DeP76sCK/97zmkbHSpilg
mLPyyRTDmOEqtNtz3DOoLrPwn/KrytDttrU7PzFtxme6+S4s6Z15H5QkSD7G/WsFUnESKAh9A+Gc
aVob+IFzh5DJQXba51kO2oibfPRwgizCbEtmEImNJZTHh8t2jgQ0E+hIZho+FWwml8KYzvKFq5vR
fY0RV36wbfXKzdGP55Z9oaRwbKIdj8+Btrw6SLVRa5jiZsNhmcXk5aUhXu7syLypN+KMgHsrsCcC
9IwTNYufV7BI6zXwvysFKxmDuDFjuVEdze7OskUQgdjj2O57EYWnMvgjSBe4VzjTn5238gc9vpW/
7dTqxz8GURD0Qctbi3Fn4XodbLGIsku9QVYlXELyhoBGhok87y0ttfh3zDfT7G6gKkypCRG2HJb/
qAxSIfUIefOXYDb/0oGQlOOYcuyyU9x86m/gz04qBFVvK5U8K5D8J0e3d25K0o6+wKtjt3z0ev+n
mNIZpeyOKbDryh0+LCKUIISOrLWy/mNda6IsbsPpo5N0ljrJCr1E2f6Dg9P8GMur9tDvalJYQGrl
+PauhC0//jCqIUqHCS01EL5vrl4ftsCNDdKxYbmH1xGZ+plgVBHyrwDAaxx51fVrScqgPpdIUOqd
wQv8CTqePK+D3W5QY6xKO8C9UtUyFywEv0FsosDG3jt0U8lxnoIMj+mZpbXx1M5oYuBjru1v9rCx
iOV1m3IXw/6Mpnmk/qTuH+8jpoT7h490gd39f3BsApWtLtXFUMB40+EmEQrBnqTyCcEeykSYqO9z
BOdYm69NP0TzAzJbFZblkGVGedRVaWzlAdFwdllYAF/yhTjzAtHkDQpKw6mgokH/2j69vfdXDWOF
ihXcbKTcRvFrCgR9uqZUii7EfH0Hj354SVgZItHvNiaiXci1Kb/bJ1d5SYM9+X98zZvlzfCZewjG
WxP5L1bMmtBVaa/hdAllpT2yF9ynS55z0q3sig61F2yI13GLKdv6V0lwI30Aj75wI+Lo6CS9ljTL
6pJcKda+QHEXqo33rcAi+vSqXd1QXwOTrp/hi4Zh8EOdJhqiWTyUpGf0txwO0Ouya+2G6Ul4d/Py
VEj45eAOvC7LWzOO6F2SvKgyvu/JFtnrp4Fq5A74ABLMEkr+dmDBDzDWT2fJxOkR6T8bRf9RK4vl
Z6QVgnxdZUXxJtAYRm57LY/IByoIIe754Gtnd7xU1Z3BMYGnzMd4SnTunG+0kL/ZeMpnNLO2r6U5
S0AYIjjI3sbjHVY/qucr35OZOsBC0xKVPoeV9DCsypmykjqMWLAfyAqUVPNuZ+mO0bivXB/91XKT
PePd2A9BxU13M4mBN4ltwZdgLT9kOOOuh7i8FEEQ7TuhB5Zp4UQqRmu6iP0LzA2PxkGLPrr++K9C
Jn24YdmRNbxibzfCGjmWW66UopXSUveOtzpBhEpn9xVl2ZRLL4FgqgqY/r0LHIc6i7oweJWs/XGc
aBoKg+FfVZxpGkzd4NaRMsBxmqoGO23k+heD4by83kKjmPysLJYUSCX+Z/j44iBRFLWwHFwlgsK4
dXEpLC4CNaKuuKNnTssIRvQV4/AImELFsfS4PEAiwt5x7gi0j1D+sfy15JFqKyWZnubZY9EFsDVn
GN01t04plGhkheuwZoE2k3G69PfdUqWG5CxEz2sJNw9iX5RBOKyMzyf9+dUPE7Srt+p6KACaZSJW
wZsi6QfbX0JarKAZD/RmfDzUfwEsz18n9mjsTc4qmEwEdTPvHXh4AfqDYhJ1K9xZRBq5f2il1c0A
QG6YOi1LfdS33BLYHSbnUH+r8M9WoOiajVJhFYfHap9mg8R4vu5/+fkvY3jx603mMm9FPeKzFt/g
vSjjwrReBZXjb9aexiRX9V65XbZPoSXlQCXTo0cnyRS12I6p46GGF5qUe0xxO/LcFAO8OxIgkYi3
1kteBvb9f+t4DQv1ov3jOOqJvgTbg0484mcsIsQ+Yih2sdXFyz/MRY6j4Vroe/n80/CqnptBwgxo
gJv4S//HpdF3zuP7Vr+7zPhbHsHK6mSXAA9hJAMRjZylEg78Cvud977SFLp6jvohramEQMWD7m4R
vV4STCceB3PeGcZe0Nz1GA0+bQC8jNqUL+Q9fP7PkeuU0H3bnk/cmbAJIbe6Lohz4OOhudYkVn4g
Iccb3dIcb6fsmqHhxMi3a+n9WHM3KzO+4kCIK01XNWyfuPKISXFwNWr2jEfVBCpz3Kz+IKzfT+OH
twhNs9rFprht2jwNDS0waEYN+jD6zkONAbcLOtpg0ZgMI1jfDK+V5AI0PGe+//WBviY0WrgQUiAZ
4lvJpqCAmI3h7Yj7jzl6yg2X6RML9q3TFTppNU1r3RQ9deF8ppwlg37AEqz79kabUhmyVPVrydfL
4ByL0HFwpUiWQG5g/5EtXqU2buCxR1eMjvE9Cj1XLC7yTtL7vW4A8Rg5zdozk/pWhSYPccRpM4bT
IWJ7zFV7lkqg4Rv6+aKHTQkJO7nqAeuEiDSdE7cVoO/mcJAKfx7+BWm04HDHPI9P9dLqMreytU6F
lzLZCyHeRzGs7nV8qNXsqm8jxhnu41TzAa7dj+MtIA2Fuv48G7MdEZ8Gr+vQBv4xg6H8dhfOG1VJ
b4FfZj/wHgbb5SRy75UVm47F7IfqDJVmtLkjKWMcDX6VfvEjYHNovPWK5zRYPmjabiSrF7HVrCic
yQ2VjLZZh/UPNwdYIkIH1S9Hrf5JRV+mD9LqBuL7iWO/rtlbpk7rcsMhjW/T+ouBLtsFu+csN1mc
tsFO6TsFYCj/d2dkVg9SUU9S8fHVOtCs/JCkZAdbQ6EQBLMrWv6+nSh+pfdRTP4YevaNzyFYu6/M
46PVCVZ9p5urrchTIkqRZqMirB4QKvPYLzxYHDXeYr9ke+yOuBUT9uTFr/5g9xG5az5urvdbrqly
bqHGcT3JCt8hhTWt5htaZPRAzmhqZ6+28LGI5byF5c4GZDH+pPwUcJUHjYQI8blMjfzGYFe+jSHb
qLDcbTQzYq9091PkqLw7YIqsXAuBCd3YNZM/J87feq4X8+6v1Yem3YnPnQjVQYKNDEZTRzl2XQAG
tUMxcFH4arCUuofUTETZP4iCcGOS5TyLewphmm7fgnIiLtiDDDfY8EE6rDxDtbeJzjIgRAOKzuag
J2pNX+drTTqLC283vAR8uTmc/p4g+BnpoT9ZRVk/wUCg7Mt4MFasxrRairQR824HeHDLlJzz3keY
8MXZ0cayCXKSIM68YZlLkaAiUayGIpsPNje4jJOsZzx7eov/Y45q2GzV5ns9Gho97lmsJhEyaGMG
pSOqSrcDIPvTE5xszcNR/xHfzCoBCu8CXX88aJsL0mvWW1OTeZ8oJyOT1Otp3N7jHQpflmSVvP1o
jPDyvFvfSGhJzsd36E/Gw3NtvnWricRR9SRbEfvEQxa1QqkH9b3LW5+J6u9HLQe0nENx0oujihuK
6UcdMfWt8dGXf2hxlmQf84LN0s0+LUWLIAmHB4raGOAoRgZtyOptC2yszSFV6FmbUMgrK+CqItOQ
HtREGPS9RbkUMbuG8buHCK6FRH3IUdT+WSpGof09TmyQhx+1ZEev5OERlb4lq9MCNzRHRjoaJpwQ
GXfrLixYz1z03fo8s2Oh5lAVu95XSsMCxF69tshror4a1E2YGaRDFcN/YDMBNT9R1O5iFOfBzCMo
/wjC91l2+5JleXsVKUMDSYtmpMsKGyxehmP2WDCffzQvXrohjB1xITjJ10YzTHaU3vNM/eZCgFVN
VBSzp9Np3qNaIdayJHCheCY6zeaz480Iy9VFP8Wk9lv9Q+Zb6W3VYDar+9JlTUT7NGjYBpei/wqv
aEDDI7Ay10RF/PSZ78dxVSz72+RaM7dfj5Gu9waSiYdb9R2tr8hThsVHBpNYCTQ9UNCtm/6+1wbh
qU8CsG9SDjXh0HxckWpK8njnbILfWlsUWsGR+uFoTbpFi1d+ZzXAaiUNsAPyp0Zxf8bFLL8ZolPj
RHApwtoeOQ1iWTD9eEzMzmFLrRfJHkPag4oz1TlyOWzYRahl7rjNXT2jySN6b2KnzNYjYcAYtlqm
swZswyav7nMrrhgTb+3FEUZPBsBAUVrYkSSbf4k/B+3KuAShPAHqjtSO5UTUpIKA4JHzJiimJV/j
uwEbiKwT9mFe1xbxo17kTQtQ8gjziuX2oibmXn3Qw7vv0qiOippoQEQWOEdU0K4AbzBKn2/F3ZxH
qQdDFRqF8kPVeNdQp2I0foM4dSuVSSwA6b2ehikoKvOinbWFY3NGRO8kqvacdHjfBXB6IMHLgGZ5
juwxpJNC5D/FhFqYRLacAXueLxANiFUHFqzH627TN+NvElDGuEEc/UfPcSwKcS/c2eJQ1RG1Yp32
ugRMgmPEu8ZUQKh3wKo/rnV3gU3g8Sl9l19g48AzFrrnEtxWTqIxpeJ2mAyTa8y0sIRmJMi759+h
0VHAp48hzj6BDZbt/sHLJsyEjtqEznu1O7OrczpEZ5x7mf8Pj1PPJYu9V3pF0aKURC8JMWlZlJ1j
6KwS64MX5gyft6jhFdl1rSYa8oabf1vxrUB6V2BSxbvtKor+AZYWCu1rlIy7eg1Et0RkbjNJnIzL
uDRzonU1MD+d5sfQhWu/dXiZXbGB9y6PpcRKJF7AgSg3Lnkw33OGSpfwfbWIsNPluzJMrSKfDhBr
HjzwucoN1viJdkOauVKhKX+USRoh9BTmy+5TULums6e4MslBj9+KBf14foGAiDin1XvixPNBbsPt
QSClIgnS1fh2plCPtih4v/LQ2EhpPtk69x3Pklf7373DNUwmabxYNVQnVskWMJlhwXaMr2d42VtE
qGkyhlQJ0Bx1m6+l8U3p2qaaZniBJmkrhsf6sUBQMDC8K4FuzRJeR+wkQWywrvBqLpfoFty6sb2B
+VXTS9r2Cvw29CiFTTTx0FzVgVEuNic5T1z6bkqH8NkGV1OSc/1rDOwXSVHFDLv5zOg828uuYngq
c94boJ3LxquWxaKGPiD0RCbDMdSmrAwt80hu5HMzDX1is0QeMXdWXAPcR7v/1cEyThqo1ir5T8Jp
Jv7ag2f4INrrw5Pe4KchAIuDNPi51MR45O7B/QSngliOjmMO+7CLS9+VVDaD+oJfEvPen0hf7Zt5
GQaCRRKWY/W1QUbgiuB0ssFnEUZbIy2Dq4fGZaFplGivxTAP2W1HtiAThCcxYwlCs4/bl4UEssG1
1gg1pdIAjstwzG4/OuzgEJraGd7tVoqzGcRMMllLoPyv9bmI4Yyn1Jj8gUvDZu8BGIAIIW1DKHKr
At2kPwsITrSGTQG1dGkU7Y+N15aVIUO6vR6kVcnNxCaRqFore2uScFdIHbOp84UseaAMcHwRpZap
DVH8cTP01rI9OR1ywXVHJiIlcmh1ltFCr8+Q54NT7xHvUf2ydwH3lM/Xeyrmj0eQMCD+H5NTbhi4
KFTe5kzzCx623HsGq2nxnZcqT4WhXXsJmZRpzKy1XL4tr6HDLoPDMyMZtgBcaWWpYr6z+P5gZhcd
iW3FfqEIup5d80WZ+NjO1VmK//i68XTQmDzKy5pjYyyWLxFjx6i2sEUnW29pw8fCcfw/orXVhOge
7X3RzN0L+TbHa4i3P4dyp5KVxxYeF2ItvMkzah0M49FbZoWGeg60v1YMdKqaKgzizBlq7ABZ13Vm
jh5G7bCt3K4H8ksNEeBkkD36tpoOvzWsxW2vtaSSIFo3R0vX5MSszr7EGLhODRcG7CQnOrfSEuZJ
gNCyUP1R9FBKmTrSD667WpDgT3ApeqGnKO1sevLyppesjAcb+JhOUgHkwzsWrLxIYPc7vyFuFadL
m+LRPwDc0wyoxtq1vGuU3YeUwftKKB1xg425bwnRNp2akNM400YJbUzRccKIS46yj1bQo+ITh2is
p4Rv1w3pVZSeQeu2vyxfxVzJSzNAC+Sfu05/uEl5ieNYr+/CQ4YaSt9xbsYy6l0TPJ0PJVIvLh5B
5R9jcrmFoJcGL42HN1eK6SE0outMwOgq/5BmBmdNWJbjF3s6d7yA5FfNc+FB/vTV4psxIecvcFaA
Pk8X1+cS8uBiHNk9HaSqigBqi1tev4hg41ObunApkue3Pq7k2bVc8tnZjfsherf8NkjfmlsHwA4w
Zs9qE0LGlTWQxqvqTzMdZFpDPpuInhcOaQ9zZI5jfiLSNpTicL/cDEttXQu07MHEmFXjE1iHlt8u
WlGq9LnJ1AFIyEq0VIeegf8lXrcBFnehFqvsDBku+O5VuvzxvFIIUlA5HAUMNTsId3aa5qR7m5Nw
lKuytpdhrD7AoFS0BX4TumBm88aQLPT+hYYktcWp3HlBi3147BEFN5Pk8Cb2pQ8+83JN5/86tvfn
AYwLDMPmXzuqpYATXn0ZSfs1Cpj46feEh+SCABRiqjEkdPA8J9A1zPebqTEU/AblfDT9uewjeg+Q
b8BNXj5GyJVW/cMudZCrCVShI+qWOcaB+pJ3pCNWePWTkv0A2L8P4aVyPHZv/Wpivaaf6QhVhgIT
tMsq/ovhmAV0bwjdmXq4Qrnbf59wFSuemTX88uoVryfFSUpijC5gdz0dSkiDzn8NCblOkPjUaPDD
aGlN/zWu4J9jF3Um7B5tkGAAdGXRCjaJfCtHtewkcbDAZMzNIcsIL/leLEiu0DCC43DJtfWTYq6Q
n4L+lE7jaicuHdZfl/04r7QjbcdHJchpzDW5PV1AttG++7vtvheGk3P4mfRFcvy1nsCc4P8qhz73
9G77s5gQY+jHW6wKZDlYvZWLt0Pg0IBqJsbCkcH7iU79x51mSaRdkpxqsa0iZvRupnOqgRIEXIUA
BwCycQyd8OwFPsx6k0oGyYqUx9LngU4crqK2mJ+FlW3eKCME+ym7mh859ylpCpVNPKFPtGV/HoEX
VNW98aIPIM19tXGSUBNEColgOZKi17QkyNLx2LYO6P340dx4H63sqMWzGk2o8qkKeaSLAIDQyCXh
FJqUyYsANt48uSRiuHUe8rMb3U4pwJVczRxDBbfOnUaVV4NqZjN+T71wZkegi8r62tJrCyoZsr04
5LWAmSWPufGJp3hjlri/GFmZ1OKvkpXF+ysgyKe4SDqJtbA7iwx3jGDIepaL11Fykti27p/wz6E4
KKFToCFuCbElkPiAddG4/LZ/JqCFxUgV8i9T0ZYeEz5KZMNoTkNszLLnt4Ditz/lnJ79OIi3KdVO
cPbf551AlEo7u9WBhA8xbK1cYyt14iZ+idhBzlNOsIsKvzu5qVo5qGPtyvPQXXBC5M+nDNYM0to/
tozQ7xRMEEIk4dwo2AjsSDeKPgZq/cmsGKJIBtFTYGSSt23LvVWB8htxcIwcN/wRq1p9Jh3mb09C
0CJRjsdpTVdchpY4ASlxZYxoeD9si/V13QkoK3vEsVZMSKgv+vdVzOjnD1MbWhOMe4RGTx3ZfbcP
/TXLkpZixoDNCa+ANvbrB3+gcLAEYq2nNNUAtNm6CThkZrjdfdF6rk9kg1xwOg3xQnYAq4Y0qfI8
bvBVlu+hNRtx+Wes/5hdIe7vjeZ14nD0cayLYAjOXHUliE369iFulnH+HmJYgN2zmgtqMKrg6Pjv
pIVg6DGdiafZZd70RWMCiDavzTAmWtpmK+hKr3sxKPFpS0cgjMilo1d1HkfS3of+kbzZJneYSLHn
8ubUFN4U4AEwqJlJcKsN2aqsaE83gFU1P+RZe0ziM+c0BOtRAsCHKp+fSzXF8AGWkKN70bCYmTcr
SzZzgI6YkZd6pkFYOwVLJ+SBi+nbpJa2leBseu5Dh4hGvlehlxGXX1fP7MJj/y9EHkz47d1VE7QJ
Vq+9RSocB6eKFCH9fWra2Or/6DFsnAw88H5fvCXI2PqzbAqG1GpnmCfXcXzMielFvg83Coap+PLl
6K+JrLnzXBXk5Tre/ZGWFbRoy4/KZakr/2J5OEyNmLbBwwdaUtZH4QtJYUALmHxtQExSwqZ3EjS/
b3yrXhELy8MC8Bnybd8A+PyBzG6L8Tz/HreTxnyGH1GMk/Sguw3ZdTJN9WrnM8dh1hAuJFvRjZQF
UG3f6qwQmd0H8chwopfESK/LkmIxnS7ezhE3bSqyPTwBHzuFAa6Rq7KRvAW/795xcpAUuX5Nhmrx
zNcZT30iTM7aWIZzuhf0GrtNtmXjEXsGayNJ5ReOL7e9/k74Cy8ZmFJL+dFWa17Mj75p+uHdtfVj
x6XhJHhrZKkvBl61KVyEzpBXeAn1fr2M8xY/4gCHKC1hzinWMxPqByoVfy8O8yAVQl1xiFLOpMz+
Dl8qDdtkyYdFegEFZMlqRqQrd8j01Cg4ilNNdKt8E4veweStWaWOZoXnyssGeqtpou7yT0GNKYgc
jubO7UhuIXr8kjgVH/29bIxR/130AUuAlJM3yjIYHrRiRYaCFmzcGKBuV5HOn6DxDIDUh/KRnmy2
XwbJIJ0kQxQ69C5FZt66pnrzLeXO6EYb15l2L2HnUgeyyEAX4VAgC73d8DJn//KF9fTIE37uRW6b
VovyW6x3jHOwqWzCcARvsT79IKKizzvQy0wICmAhjNgW7zJwTixtJlET1+U5eimgWOUo+K7t6Y0Z
0zS8ifP7caRsufHla8x/65HJjBSh70zc47jrvFDDlJe/cPJNovygoiYWnkB9J/cxIiJZAMj57qwT
WTQfhKC70yiKORYI9ECk8GPkHiuj/QNYNFRAKfLgrCUubo+79wpQTJMaqKEtMWmhiNMf4aXeW4kN
FsHtmcBdbg6gYFpCb0VHxFtXpKBHCUDaXbpY/ouq/fFAS3tmD5GtN+yMD6VT2Mz+mwuLasCxlI5g
1X3LtOobKQVg7UTonmr4qTsTn0HCr945oNRBhKgVTr7lvSp5Cafqvg8+XEPMPKWnN3pwiBb8YbmO
1ngub9M7tQUAI9PMgkCmjTnM789qCHkmT8VGMGI5uPV4CWEpnAzMC5phySywlsv+qTf4j1F58ygS
Wc7u8OjNiOL3QJIqAJIexZBI1AboP3CNNIHV7IBxD1U5K/uAAcUjPe7+DTJ2AqtvCiJY4EYovvGP
rGpiSJb17CURBmsBQRu93o94TTHS1lEM+h7IpE4tPlN5jOIfYOSZo+JEOqGDmUhkqIPPjTJLiLkf
OwC2RULhocjZmYADutFBM+NjgmjEwEit6uDu1ARd9WeQeqcbPRKPUfcdzw1L6DSXJNU3uTop8LEs
4FISGZYIbgA1yAy6tZ+93nfEjqZVMO/pFlDO/Ocbp9mZBo3eIi0dwV1zrHNtOCRrIuJgzvTW+cAV
tFlN3MWJSLyeHFkZbiarrzgmhVDXiW6+6oAtti103pOnsHBzJwlkP7ssPrbdw6ALn2byI/3NIVUK
H0CIhnP4m0v6tXR1LQLOxlWvC+EkKuOjoD5HYtM2kqQ6lTWuvpeWu1ExOr+U8dbPLJ4Od4g/7LX+
zMyKzfT8TF8enSKwprb6uiKpIKoixjBdFcL7wx3h72SmsIFtivit+gw5fuv3r4ZJ3HyEuLFkIkbM
FEtmkKbAvy220+/rghxmeinsx0yfBlv+a+t/HPYAaVd1JxooVCbGKNZzlp4BUmyu7sgmkZTSgRJe
BEQYiXHMF2sfgIbWH59VK5USPtZFwy7uIUA0G7WsqDCKOXPGVbp0SzOx2R1Kw5LP9dD3bd1NsN8R
S56M7PVsAYaxqhQKIMx4iFUgPdsBtIICNq2yNZHpZTRqhjl079TfBzjSagBzMRMAxoqkhgZdtZx4
dUOgYkFk2HRFc5L7eqFtssnROU8lxeBueu/C3iJtUPZTjpz+QT5BbqYZ7riCP/FHUSL8yKqXHUNH
wejrCD0OvR9HeAhR+oBlj49fMPqFADT64qkFReAiHMAY2erAfePjfnRmxf3Te07X68EC9x7wyeQJ
eImyhV5eTKgXq8M7JyMgHhl6NDVUc+j6Nwft83XlA1DPN7nMTYvNUxR42+GLIvV4sLsSKdMMqS3X
+ivfpa+D38D4z4a1U7R9thZaU/yD09l8rrHbFU1olJbsiO1Y4nccEiPQeF5/QFNdlfZBQyHthlP6
eb7PWXvMuyhhZQkDDyg1IKYkMG2zIw6Jk0l3924GcEcIi9Lo2Wj1foHUhtZz3KL9l4OC/bMx4o0o
xt2xlJgyd4sYM9y6PhoYROkLCdHfPONMo7zZmBH0shMNeXtdT3eQ9rt9Uj6pNdPpMPo9eHeBoCf/
4IZeTK5a0Iiq/Sp9FsZkf+zYlt1gUoBXTPTusguKOQ6VGw2sJMYihZX0p/1Y3nHQm4h1xkQ6Rxbh
NxxV+NvU8yu4Xwqy2oo7zBlG3IZv7zB6xm78XMMICkQfndCjkDCsHefPqniKjAFcfpFXgsmRU4Ph
ZvSW2kYx+ZFqieWZiX6GaYAs7h/Cd1ahYXdl+18f96FYAUQkZnEHVptuT+U7/JpjL0GBPNprraDQ
+h+GJVs+dVaCAOxMnQQy8cVI/p8DuoxDlRDCpGhUfYLvUqASd2OisRPjFI5PuYgd0XNYJPqnpeRQ
neAe3iV/44JoTYM36L9aA1HqoIsL4HnVPLaPQ65genpJriH6XQ6C77p3HH13X2AJbW7IhqVHAo1F
Q7wo8OI0gNz+y7a9vLBSZgUf8lBwukER4dZdSj/LUBzYr7EewoPZsu4f2BYAMxesIaTT1ca6zgI9
v3ZOKhG1hueiMQ65eS17qunpPs+0Vk+Y9k4DB4slCxID+R9DGVLsaBvvJ8QS435zS/9U0IKguSlw
yfbSr1ArELUjb9ITJz7WCl33kI88cUNGR0wZ5cqG876mhTQlrCCkexuXjSwvRxs4PfDX5V5rOV64
rUOBy6YKBB4w5hLx4vL23JtwPKX/z7AivH/lY+mhdjF0lefl8Yq+Vc43SAGS/qiJFHQzGgbjMuOf
qxPqe4UiV5U8Sp+4z/PvVvwebjqqare9u7xV5uJjFZP1JoQZuJl/ifzC0rXmMdaCZKxwwj3XRKP3
gOA86trSX7h6rPeWXCFgrB1oNGUNWt3DV7hT883fQc9i/q+2TR8hg1r17VRAgrXr03fQfIi1iqC/
IMyeWDpSoEVS9/kFdH7+5BU07ifhwXTMGUrwakTaXDErJxc+iKkP+qE5XS+yo1z9d/e4grXhV8UD
yVFO90RHBQ6mQGBKZj/V4DGPq2PUJg6Hp7uVDXvh/Jn2liaAFgnQEbMrPtRyveqtQKbbeRm/UAFf
o90D3V6oL6f2U8yb866/0CkDYy9GOGLuQIKMojADFawGOdqOnxK/G4/njaLxWtaZeOUJnNomiKmI
BCgi61ZYTDjec2cyyrsJFmGPNWFvRV3tct9k6gWP07f626IQEzYG9rnjOZoAdRV4E6h3e1wCs5Z4
xCJzhPNF6i4GQ4nYf3vmBcZONYrZvAL7yHZNPT+MZ10cJJFkuheGnoWbh8rVVGrvhGi4Kcylu9yu
yqqas1iZhlYSvlllh1hlCSwsj/esFviaxMfchTH+5aYrFqqRdUe+t3svb+j9MU2GGL2Spi21Olp9
jP3cUAgYylB+fHJyJH6xA3+WwkKm+l2pG1VKXGtXsUuSW8l3nUfl7faxNR7kKMg5kd55ahHYzbb4
eDwNJOZQV55p9fLc7LnVf0qCj6+CfM5Vzl+e19Hia0e0kYGPsRwh7banhPkZls7BDGNuc2r8T1tf
zreLy+edtjoKTtQ5i793d39z2Lv6c+m2i7xJo9Ssd9zx28Ui/ogGiaP0ClF6ELyqisyaUrDq7goV
6p/new2XI05NMuNOdZs3+2LCckaxw5ZfOCose1xWFnhIP7jVpjRnN5rIjl8IsvnRKJvdMlIy0PdK
TtWm6uX15l2Dsk5rMAg2ZslJpQo2iECU0i59Y1qq1mlursvLZGsAePWTs0cWcGdNoQ25+Pqz26Uj
CeIK2V8AkCBFK2+d8zfuwpkJM6q0PiwgBFwS7dxYBQowbpF0H1zVfX4HkCA4AWV9ok6GhESesCMZ
u7TCJZFyQPh+Wo9d4wlePOZ0GKzaOslFdgTRrIskhYqEu4ch3cBupVt6blbCvgr2ZlpHVSkyht/H
a9xy059obNaoAoj+P2zaUTbMiDH/fclrjm1mtuxf0tKZ79LsgoL44YbR4rzMYhzLc0q9yaYHi40y
G/2FAf7jlT72VqLZFg2C58HKBkxjdajBFeLdAc1ObBRzsG166X529JiF2echbDEeEfvjKezYEdkf
Tj9B8822hIeIjY0jogavm+m20VZdKweAigaa9PoOA+rfQkCC3bwGzszk3EE8m879k1bhyFC/Ks/S
l0TdEto4uI6mU+7LTlIa5VNVvN6+VRemr5gPOWJTiR5tpSiUsFbptkA4buVJA6sZWB1FMNdl62Eq
OsIA1F151suBo3aJsxYHkDSX/swTG2d8uax6TF8vrJgnwSWizqZywyOjik4e3NVNYhI88x2VvuuT
FkCKMkP4X1JauuBELo1uxPiWKDBCotiGFCqRW5ERc9H4XMjuyKW7ilnAvsDjMZmpqPhs33nuo0n5
gEyFCaFG/3ho5DHAi7mpBd6YSBtR6XeuEa3VKs1V2WwUCFetGO5vtTd9xT01agbAoIcXzJo2TGIa
hTcCjlkFInLcLwkds6gzWvknIuCTlXTIRjNGWW47m/lLpEV7sOD9vA1ueZJ2kTScDPm8MUeEFXb6
6ixF9T6wQVjG8zyRgM4EKQ27pHYbb63yBbYW3M5fSHCiMdgwtw9mMqigdLRAtsJY3WUCFnvdB7cF
UIXTmTQyGghtN99G9WDbIxt6xp7VhJfAIfcigO959LQwkwZ94HX07vvMMv6tpq11KzPyVIhD34or
iflDgebsF15gSN1wgiOCfHXNpkiORi9I2rVBEM13Rw7IzND+faJzrSBRrlBMvg3uS8jDiYVUW4DT
Ws/vSStVL8JsG10lq/IQL0l3Vp0m/VmUlrRxC0WyhK8ObPvPYZDcNkwZSmMJ9Zb4TTtFVp0HrC1Z
2lu9Z/vcbow7LibWdGtRxQWGKtMCWentEK3EPGT7q4H9gngppx81+5AZct7bKQsRhJYZfKBDJpSI
UnEejaag2Nd/ZmjQ7kQfcG+ZjvH8KssjFSUNfBN7/xeIr1EqTGPGfPy22ap1E8O8I+i3/9nGLuBC
DIaEtZzA3EVV1g6kStXEVcoebb7WxTf9CpI1tEK65FppwkNgtGxcJ6VNa8luPd8GaLzz6NO2Th8/
veeSgKB93qmiZpVIzBJBL6zE16HnKMJIZ5poS79CPhm8r5wrBvOh3jGI+20tRGIDLhBMMZjXUre4
KREm8dVPGwy5ZIdRnipZQNPSA48XoCdo+hjnhlezaGjhY5X0XRdo9mruqiVbp6ZXJ30s0yVxCjA9
LliLsX006/Uc/5z3yikEgeyObPtxVBIp/v6wQnvRR2VYXrO+0ivoTkEsgwTof77sKL2bWc9e+pdL
66Dz9S340es72jpoDNb/qfY7F6DljRnJwKGJgC10cEyErQdvrtfu4iLb9kcpxLrD6WkSnL/TaJDJ
Afww8Fmywut/b10Sh/IPbhjDCZcN3Sgam7eK1dBxNI61UnPOtJUpEv0AFXmxREK9O9/RtyKckfkT
SfQwQEhGoTgTKI7aQDZeZysTWoA+7rclbF/4fE4CyPQrjxgMBb7xghpGj0IWmZVM1lqXIXri9Mec
dHXzcm8b03vqfgxiG0xcxLELd/RLV+TL6dQAvgwzAeunU9dNPozarZfQJPOL2Ph/qWhBL9ZTRqzt
1fpDRTV2wMAHvx2mhO4vBNTALdjfPYSYuB9x6FK6TObmKsU0nL84Xsgk6H9pHW65tyJtBPdSyklD
rnB1T9iHKTnYU1NiLucmdH1KUuZOORVfbO1b03zjTsoefVNVISXDQOl4cKr1DZQtfUXrDA5aVr3p
tDlcQfvEf0BF92h0QlQ0TPEFpPRp+MwtDFVvyrBqv+KnCK3xr+M9jLtVx8w1IL1mCrKhSVlvBQPY
Vj4eLBggz+pLpnrJLg9FfwphAwtYgAKpiJ901fjusNp40hJobEHzyzTKUgFz17dD1shZg0iREE2G
dS9vkESiRx9wYBpFkJR/JXDr53ufUgOWUhNoB5W4MdB88c0KchM23cnNwFo85Awv1IOurak77FLv
HLkmv7vozA9zDXetL4zmPG9Y0c5wbclVIJKcQigto09+7iMvNuOEyeayVzGb/8EHcRhtnxzVxci/
ekJNH84pwCT7IsVMrimCSk2mfdz7vGqYMpm7wkVLkdP55hnPbPo2TnNv0XWsekUmTMao/vlvXMmz
zURJgQMPepLj8h/+c1/okKhnkTrwWdCfA3KwFMbq34lHvLFfwSM02oYWtygz0MRMT1N1I+F3YOPL
bZI7Sx4e9VduHb7fzzGEQDNl84Ykgvj3KHmVzXGI0mwxXK33n64CFBuXuMvORRpY43RrZ0TnAmDk
PjiyxYDzNEYiJkHzr5DqRH+kc0AUr0Xly7TSp9xKRg+wTM/Crn47yjPeoG1ii52xl+nS8nXP71uY
CTVsZUD3kts9JC1f7Kq2YlMDVycLHz3Mvov3TQuVJCSb0iuFI19zGPjUoTKUzFGoyT8vD8B6wcoZ
FXSsP0a/7K/dfhsYfvAs7ljWbcbVucOSW2bD9v8XHOglLF3yt8I3MXkqvsscrrYVB2GOHFx1jdcw
x86jjkCooRj0q3MJOzoKdEl87MUlJSVYAxqQ41KnkzOnP5KYijo1PWspDqCvYuB+1P19Pk5TpzNV
lVOk3aeJKuQiPQu5eT8LZaRYoQWyw8xZq3MvHiHx+POpphylbkbmiV3hRIPcu9pueLLVygyolgwG
NTDvSn7NH6WghBihgLQaVOBKqE9/L5Is81RrcO0w5PpbD4+LAcE9ASOifnyRCB1oXjR+4kxcCMmJ
lMXBkjYswcVmWpjEPM5Yq55pKSRE+K9aYLUBC0EXugwKVH2JatovluA56uwt+bPR8/4bGRQTQ+3+
x2zrkeitC57BRFbEtqZ0TzXavQdh03WszzlDq+N4P1oDzHkyjawdCqTn+zIRBKMWn5tTdt5TK5pm
RBQRKOhCehiXK7MRtoEh+rfGEhWu1evfR2mx3MqYqmz0R+7n4kiFv59DtyGOF4J/Ck04TPMhqIe6
honWdkcfgKZ46/Lo+x+fFNF09zUP2ZNcL7QM2J+0TEu0a/ptpYubkbu2hKYUHa5SzaSO91wAoyzU
D2bUEGcKhwVmVxGsD61MeStz5tspg31knflBq+TJ80xHuemlch377esgBSAtHhQoQ4iLa2OIHwBW
+MyozAQP33IkxMpP5i8BpWlmV3xL8Q2+b50iP2fT5p0Oqs5sqTztKWV4jh1u9r+88GHx+o0joS8Q
XwcVYgBEZKhNk4zQlmYy1ufX3MXilk0pUmz/Tv+xUEi/gDS+lvhAjOXQrqnr27mvFAwcMxcPodbv
jF3HvYFmm97gjkWhXZ2u7cAxYzTGKaF1KUQIP+4ZK42fQ8U8lN1IR/9qNeUyICrciPmucvG3OzRm
TzV/XGPLOwH+RZM+NouVXXIqc7XAhaUac6o7ZLvGHGjC3Vb639mGH/SbPGYFD6Cbvju5hU24RBoe
zVDa/QZekzblFFnOn1ZYIfEv8lYpKr8WzHvoGQ1w6zzrRBfU4RMx3L6SMJ+MgIsat9YFduRnVAW+
VU5MFcWVFedjtGZsRry8x5MuNMdJhT4BvtNC2hNDfjOjAxMY8jSxM9KxVWdAj0kQAKpy7w8+iXT1
ilxC/9kuCuRHXA5PkVxUoOiA80hlZDY9y5Xirc/CDG+t8qq0ShI6oTvFbUCg0JjR2lX7zPurkuLY
kUXFl9/1zhVBD9yhuodpy7M7YGYl9SeeWfPNbnkCoPb169Jo4a9ULJ6NKnXAnxD6/WpRI7ud4hQd
ymyMmz7bkLqbT1Upn4LRgs9C0bQMK0pmzkwQMp1pDnRfJkwKb7HTz0jeYufcE9NUIwyDkHYOKMOn
0x14AGjweNbVcOAMeYDD4MlC9l5IGRUl7xGl6X/97xecUXNpHEqGVNpk2Lj9LpclM78ofAAjkeue
MYirMvmFnRlZbdw0cEA6APx8ds+AwQhEL+oIa/DL6CDontedoqSSf9J9OmiJX3oubbStOeovqHoL
j1043Gxm1YZ7/2OYoxJqDhcATAe+CG/v5vb3VNSR9uNPzpqZeipUrpS4E4ekF0iegIvsvvLo4bFu
DWSJnzdUl4cDFk4e82n57PWyZn7BJ9mfEDCPG9Qypla85PeOs8I0/Tz9/sAzhrIPadEHbpFLNNyj
TfCrEHTPcLPNoeJ6HYzSRPVgfxZVUSnhJrITAVM8I/KJii0Hp+TrlPj6Pyy4d702yJg6ASy6MTGV
fByAoYLGQn+SX0h499hDjpaNBxP5FlFSnMg9yqzTEpsJOQ3gnsASz/GfxsolxAVEB8fcr7gti0eg
3CfOgA7Fcu3uyxVQbPFqul7Pk2eWO4iI8Zl2irSMRr4F6+4vJ//MQkD5VHA7IDQJMD+KvcLgq6cA
r1SVJv/gjNhp1d/lFFJEA9a/SfxMCIUFYXM21mSGY1s3tnLnLRHh9sVmBjxLxBlZBetuCgJrtLJb
GIpkSPkX7psv1ELRmQz1LmO4I0JTfmTfSq3lltBtF3Hdiv5uIv2663VTW8BCBWC5IHGqP0aGzwbD
jDSUXiw1fLQQpGc0dYDeeQpc0a/KQMQRs+lylWyt5KB/fAle20jqJDC11dGC23mlMIZT0oD6aLhd
yNQdaaRhIUHl2ox1qx1/otBT4L6HsStTwbP5F2mCaXcjYUNz18IkGfkj9iJjei0fim8Hpf3jKQN1
F9rWDLw86Hk1vnb3vFA40FHCcyBjRfJV5kWOD6m3shHuz2l4ptulQ9/Fza50g+hQJmvkq/hsMmDN
5N9biqhbwuha2BDz45oleoO60U9djNQdIojrrjK6ma/b4MpaaGgGICkYW6P9CjuKd4iC3vr0X1AQ
ZC/zzDAIhqJ8NVWCXp84kB/s9o0Key+sBDP8PboklouDDjRhfa8BUbiIDY9KtZ4qehmoV066+sH7
idqk6KeOKk/M9aDfc6Skp5Q1I+7y4y7eybkWRxzLhsLfOf39iwjVH4LEjls98U/DiewqMjqzdy7S
qi7CeqJzK+i094FIhgroq2jzC3kvzfpA+bzqD4QA4+RXUmM8vjpGaL//aU+IccD6QSg0vNPHusl2
WO54N6dUzrz1U3nj+cg0ekO5ZmDdurB4ttLipqXrZfzNCQYZGR8Vwtp31jl7qBu8iBVbPqvevrxr
W00QfraQAyPZBDA+LjvEyxCGRpHNPL2qygZmifGlse7G1DHujydN1yIxlHgicaStc8OCoXjSinYz
kmWB5Qh6svNLpVcGpMvpLkY52WWnKafBCNfrXF0h7aqN2JjvJb9+yu6toVFpKOqjZyOyBGPPoX0D
y4bJipKyxlR9FLBY8tciXvNFDA84h5+0ubDv/P91zfwGJOHjjOeXZNgCXkjSzcbuSU+ixmzzXJjh
xbX1m3DZfiNeB3P54KaUxfQWwMQL2v42Ubp77h9SIXU3G8y4e5OqRPAKsY7VF8VtzCsNUuwVxwVZ
Dp9eP3lby1HeDNSjJZlcIRJSwdfOsyCqUsUfRgMd2IQa1MGHzMPqN3EwbSNcSFShird7Ku53ZT+I
KRPQ9FbUY+eqgVqd2Cyumpw8uJYr9VmtIYjdfkH8bScqHje6bNAjzNrvduuGOn3fCeG+4j+b4PXK
jJGqgZmEO48sjVV6Xzppyw2LsR8mG6vfcYHlpKD8Vf75GY5EVTKRJKDfRWmP5/bPxDTyVqUMrxPt
tRNuNhJY8AXu349OeqPyr5tKg1hpS4dx84f4P+zXeSlhBOx7NMWT01v/tzCTO1TCjrK0TAft8O4N
tmEc6XsuOOmlKUijiQC7InLG7P7Y0PFkaU7O927y0g2gTTrEJ90vUS5+rT485D5rNoNDev7Rg3Uk
7Hd+Z/BgSOlL+8Vc7l2miuXeVboLt/CGxsqabE4IAS6EqVN6g33V4efqcWRgn07Nafo6h8epw1VL
gKsM1crCGn0I7DhWg23piPMySi1V8bM5/Is1+3lChhO40NMElglMgZwuouCcictji4i4JO1kt4XP
VuDFPUHBYPPede7ahJOUdO6q/HtMo2Gzlb56DhFHXVErr+5YfXeDjTcEqVGWxMH/+BCp1+6nInMz
lXVfzUyBOv/1+nQAAkHi5p3KnlaHO+cn2+56vzUNSrcLfPbtMeKdl/bWqXzqoLSuwcAKha2cXX+Z
I35d9V2dHSDAvaMYpBuWxbCDM6lV70ZF9FDkM012g7BtzzlYJuEuasKfH/ATrzIQAS7wxqvS/3++
gNyITDmwcsDCnU1oSefUDh0p/cpTrpPGXyK8x6yZxKe33AEObE2+mgyAxMUIfK3o5JsL1+6MuUMc
+oKrLLFjo584zNaLsstvUdUIuHIDU0l9YMsTRh9FI0TtBcz/sXsoVhTIe4WY5f/botCLc6tLtCBs
ZInLy4y16qDOIYlkHAgInEI6bQb3if+g12kTNgGjc60p1xlwMA+GmyOwWJdCeZYqkYDUaAiVLeXs
fmlaATrTt4PFrrk99Sv0bdoiRRcPq3IKBCUsd90LxQPK4D/ya5KCmALzRSDM36HXqSYWdWMt3d81
2nzBjKlx1q5jnri7e9QVLhvtDucRrLhi3z0X97UuHFdQnpFh/KzVXAUv/8pN751NXMyUNJtUfDo/
3f7OD54aBphqPnrgXJYp6F/9FV3oNKhbK4W7qVUQk5pffm7xfZgXZEOfbCjF+TU6EwN1saehcz0h
ORbXlxA5w7NaVuIQhA6g0GoD3ftJOwmyCFNmuH4OI3GK/6eU11OijJpDEcPpH9q/LsiJJ+HYwKft
12X9OCs6uNzWkRLyhLDOd4NWO92x/Lwx4Wk/LNkkmhq8SZaPifF/Km0hOgx+aseZMj+aBWK74lOE
N5LkCWZ1sZBb9LTjyyyJuptFZX/XLye110JP4DLqC1keuxaSk/CDKFjzGnyWeTBObLhw3Q2QU2oH
FSjbDsDy1FCM0NUBFepraNeboKMqJ/wz0uw6gRIxQxIeW7dqw0YHHmWZrOq7YUneBP2qbU7CNw7o
WFST23OyX65MScapPvSs3dloF7IdQ6hd3TGy03D3Xswnc40UbH6Mh9Kik/Bx0Yvd3gFUwLqWUWqL
jCq41RT28g5QnPZ4Roh8Orqc34fhE6M20OlrTB8D/6/vLoJ8Qi+yKZH5SvbQdNHh3y9bKZoqr3qA
PI0pD3FzUXzQMAhkdaF7ZPX/E/Vgz+njMp+AXGQ7knN9oGUnbWALBRtc0qD7QSdqd6vMUegmHp9+
0LQkttVVAO2X/XHFAK5mNX47ZfXBf2kO5W6DhIAHSRIigAkcepD0WXByNx/sPxbVHri98DSwYWdx
bBzBSBTVC10vp+f8GfWyL8svO5Ow50rbKoMmyUMb/3dAAGPljbRYfUy92Wa1tvGQhvNZvJOCnsmb
kUdOBUX827kVBZ1gOzixS3CvcU6E9amdSWX9Vly/vjefULg2Efym4qZQVjSi8tLgYO4AZhuxRaY+
qfmgBhwQuofilWFf3Y8PaONby+skRDhDEyVW+geBq6mRbWpOe5xtn4QFZAeY9nxnh8HkYGwkRPF3
Zv1bh0u1mHVajCZr61mNiwnDMkeWJp5YwVcpDBmwGM26MzwQGxeTwckGcht67qp7qS5oe1dofFR7
IhKvchIyExxW3YaV5HV+fKsHD0rSa9FP/PaD1/W2FTsWigEoOVk63MFGQ0ipK9oXpapMrGxmxrP+
19lu26njXH4OnCsHzCnWg3fFET2p+M9oVZLzKDHS3ZhufgnI08II3nhELHw+jAfedayH974pcYrz
JRTYUcwI3wxHjNJhboic8tgCbIQaaf3axhZSwOx92GQn6VMkO2g0phRpp0KQvBjnSMMY5Bv9Bb8m
Ant/ho0SFA7oUBrs/nmIw6LTxi0rFJv1yZBnyWwgA8hXcBnk8zaDmNxx2X0CxcEqNUCyxJT8f+mT
hwNya8TYlD2Ug80oMYb1tJ+lQbJtdbUnfMcJ6ZwP844beEcOwAGhzIusxHECws8f3iI12D82Rguy
hAjc3I/xCO2hm79uEhv1NcAljUNuByimqSu0zYkR1nFGH1WU0Pf7DXvPcMhUyIFXXxA2kxkvyfXF
XnBE0jyZcU7qrCao4agJkG3Xs89pEIIh5hIREleAakUsJeOmaSv3gLfEpJn7Q5Vzx8rNeUxVsZfK
Zb99ZDLnPrT2HV1rZNUezk7vim1tqFccPybkou6LnV5e8/atgyHNZjXaEEOWn13DOXxWFKCaemYT
jx6jG5QXZE/1lepvl8iMBEVVnxf+KwdROdM27Ik5i5/CtJnrWSVhywc3MIcRKJLyH3x3Ldv9q43y
Qayg3fCVFxTgRjS3MubKHgxKRRyJiwqj03zzJagBvGL6urHujC7TU8/dLH8sZWKKLcM/7G/ZLBKI
kwK7wG9cvfvUYQSOtWiPBTsOGM/7MnIkvm/hvitCNYI9PRY/DOI6n6z2OUUm7L290rYiYxOrOWyn
a/kiu1CK1IXo3dVq5x6IVjysrdJe9OJQw2cY2JtDGWsMsPaH4k/yoI3riiZWYd4pIyZM7Q65c7PD
9q0C3p76UHK7zwPLtmaCxqqJ9ahFSTBzhm1Ip7FfqOBUGRvLIkTUA8eTK8V/v6F6kHPaA7z6fQGM
4YZoWvhl9kfgjttCqEYgtMvdKt24QEKh8FLpMz0Ka0phT7yBBIrHgoH1paoEH68QD61mS/uCeiZ4
wuSC2HY7oOzYtdLxhwilczbBxrT6cQs0scO/FEKUUJ3JsWSkXP1jNMWLe9B0SeZMY+XU6IbDJbVs
nh0H+sXvDDW93ItxnL0ErK/T3gBgZ2mn/nO7+jQ0QqASMP3sLKYKFDhkxjL86lrP2SvTW4KoIUvp
PPYwZl3zjxzZWjZGZZrpKFQKf2Vz1aq513Pk/RTlYdN1i1lmWKiH1OMtwwU9q3gC/Epzz3P3pPTK
/dbEBuSbA1NzRf3crNpRz6suajzFB7fD86axq1V7RZRw+MJmdI7PQji82wDqWXxnfd1gS4GISpTU
UUKGkQsh9kVzYUT5v1hACZUDk+Tec22eeBTtyQJIVYEX0yIBkB79i8+mYb3y0vM0m0PsxRSbnNLP
jtxOPFhzQDjUSzE6n3I4WUSf6GyLJZ+ykyytuB/LGL0Ye3gK+SduEK7w0fBYRQ9xKbD/3WpU3V+g
PhEFSkGlJbL3Aa03ULOhJemtYcYCShwn/zNa2ACcPltRynd59UcUMlnAZ/ipEtbpbjGxoMkffB6W
tSIhcDdd79obV1gafO4cic9joAg+dJUnlVfUxBbDFjEeZmH2XV8kmW+Ov7EjnPL52yLFhMt0RwJ3
5/DyjTXVyZZpcV0Zthj8RE82Y9gWDhPUhxyp7FK/qu3eFoiruz+YhpraOSo/gVt+CUqq3jE26IMB
lWKMvOzN/UkjdYIcngqZ98gKxvRoynxBhB0rC6IiY5kULSbfpcY4eF0cCgnt/UT3CWIqROJ3HBpx
tKTJkqXAYBugvrKveEazT/qr/V8N5V+i6BHdlQcnMSkAoKjFX5JBNLpGdvaCgKWijMDw0iU7L03o
rnLSumpCAe8S6uSJH2r9KlZ/qNNyiWWymuWV3+rHfeexMZt9KYxyXovcnT7AdctJd32VTsVPGFGT
L9+1cv+7S+czleCyuUqsDjgN/JGWOOu0HI3122wma1lEs0KvNdZEetyvF5uUT+pO+KQ2X/YNkaEo
E/8+j5rJPUkdoiTUB9j5UIEut04OkaEG9+ZCnW3xN/40tdzV33WAAw96qOA/P8o3rmV5z2dxg8Zj
5Kkur4aMrnwfSkIRqU3yDJuH0OXpRTubrw0rYPz3lVjKf05VuPXh+RcUwW3DsNYxKxkui0JKuecU
7Md7Lbd28wEjgE35pDal1RIJeEasHyVTtXzezMfxeWthcflV/beWYZfDkfr38FcFPLXyFmDrg3jN
LuD8NX5x8vE3Yu/+cERUEyKAlYlShZXR0pCusw6YdVnde1yNwFNovIqA9PxNYDlCBkYXZTfGsjb1
2bGhzoZPJZIXJgAGXc50p2RqfqvlqS9l1jcKBGsEl25WOfDyi7HUCHLlxznLYOKXae+wJ50w4T6W
afEvDZHHdEaTCgqnhpO1e4ZMvIWqZ4hvqqCZk1Y3ICw7AsJt8SGEzdFvZC6yLwsZ6htcivsZJYIJ
SwIK6yzAdveeI7Vnxg/1ILRVJScukH4qwMnrlyTVVy5LO+zdfnC7GWEs1pffWkE2J9YN6vRwmWlr
wAWunlgznngFc6IXzBiSCswKWFtO0KMdtY0LfHi4DXv/LYKe+GxTkA2aBHF6D3F+P3xZCawnG6O+
n6gOhp26HcL37jr2nMcpAaAOLgyLsze8OPgzYOoffEg1SyGIMmUKYab0Aw0GiVIL10w8BAMXpghp
4ArsQNp5JsKNDu7AAyemQOcto4Na6vQ4fRk1JwISd0eAp9Tr2sanKOPI8NVx6r5HyBc/5Pik8rel
erP0KjY7uO1K0OEq9sFTFnyi/KDzrnauAOORrMXdKg3CQtiuWcqYiGb9Cb6eVNHLkr1nhHaE1AnE
Jwj6yyjWOO8Xyo/Q8idWDU8DRpXf6lMZTVRDmcF2umjFSLk4bCvbqFDaJj62Wvg+OGix/3AFnklz
MH1+flXYMALn4sP/8mkWVQOIQYE+hUz06eYT160fW5dgA5wa5JH0JvjCV0qD73wdrV3c/hm1rQpc
TrQj4VTP43ibcTXxK0XO3GiChfAZp7kiFMEH2AiNl4W5XAlRUK2bK2vfEXZKn0yM0Azlugl3AwSt
v9+BFA/bBir4q32eWZL3rr2tV1xzWEm1wCVx71RrDFG+SVAWV8ZcrLa524v6C9+mde0An1R1U0TZ
TsJgd0Lw+wM/WYxcM4N6nzlg/8tCihFs370hEOJWlRAHB1DyQUbOpWZ0TPLcol/GDFRSa2PQA3Sf
oWg/tJxTXF2ntuYCXoF0NZJQjA/qC/jCMVITyuG073mZck35+tmSCig3l8gwsvyxD4LuCOLRE2dp
NezzMH2nTm/NcCsYJrcXX15NjQ9hClpnFaxMrjaulI00KGQOBCScvcwYa3RqzahMJ2G8cNltopLz
JcgIt5ks0DDt1yzVYFV2Kk4aqJUDV/dxyFt6cRfmcx9qCjqEegCEx7NbmgVXS1fu661p3o/Zx2jQ
p+Czd/cIbJiQTTgNGWZQ2hXCDD+vFbfYVj7JZeoxv6GwpJmUsQUdznib2WXhVYiJbWjFuAcXgIZC
0MED24W7hdAksMbblgTNusGcScfqXMvftTH2+Q03FpKKBV4gvxGuT3F4d5EtUIRp2PlLhlvuARtQ
BB7UV/KUmdqXFF2OGd7+a95UEGhx3qVF1pDuVa8MVgt2YXYZTz/iW+r6qzdCuuFfzSTycPWIpHtt
ZDP1mzM+tKWXrIONL2UlZ7oBAftn9Mh+M7mV2bvwjJsF2iEfkpCPkATZGI0mC3tXDPiki2+sNMOq
tLcythfjhqnLuQdjy9dxIWvPYy0gL3dlHB9xTGiiMABG5qlX0fQ75AvMJ6LX/MLbu+rNDU8JX//p
BdOkkPNDCfTj54vgQr+34jB7IEyVOeW+JyXB342t6ssNtXXsBPzlJ8e2hou6O34v42SRQ98hI8Pm
qHsZ0jTVuyq/hdr/WgGxVzbbfD7kp1K59OdxBbJJrNOaBsGi+q2oUN3amYjtEeUu846V2UVy7ATv
kRz7Dhmne6pj/rZhriV10X1E0Dj7LWFFC66iYSgpvkOxKVmI7nyv//ST5MGHcqHEApftmM8O9w5j
kYsAyqHOf3EOFK3HAO3VZF8FjMcOeT8SOVSnxyoSuyh3Tfw3OA3RLG6GiMDyT9QNrOe4za4gDSEY
vGl34xIv6EmxPV6WyttOgeKhmzEzuHtuljZNC9Tkm7ASZadzhqusbtzqmBdilANknIZwIbNRexUr
36HQsu80BYl+1Os40uNes8Sm1VMTwfRgozt9okxJaU1F/rYaCLE72yjAiI1vUV+abdmZ9mvIP2PL
d1ptNeU63KbMqUD/FiuGwpUk8xBgbMF2zUZ4iO1bhnc2f52zcx4r4bHAeH/2PQ8/X+ZeqgSpM8aU
Fp/R1JfHtzJrX8R4/QKTVmR85/8Fbv5yfDZnfmoEE2EILw9+DYevvTFhgKYSyp2wFeNzY7vyGkBE
AnY7qXyUGwrUSdQLd/fJA3Qwer6lAMaaLcitDER028s4rG7XBdTJ16m+u+I3tp9tUP0t5p/95KVx
m0T5baltNs/h76zofiawfI6aenhVsdi0aMxUu7ZyenybdfWBT9s2j+5bGqumNrOSRW0Z9NcWwfe4
eB69TAQ2PWnfdJ9au0wstJu9WKq7ddacFKafK2WCqMoj+JW7R5JG19a71wv6IggBliP0qPO0F5uE
6Yfhg+PMwGclzMcrWBsHgs11mrIFBO4YnpyF4jDKCtma8kIHoiWk4WFeGdOafKVWSTWtbziKRAkM
r0OHZ77Patb4kI80d2y0XQk7qyACR5Zk2o1qOgn5tu8hPauwsK26CJar2Q2xgIjm5z/mBzr5F5cP
dUKUo6/qrSKSM4iE52jsbNtCHB1gnLH6dTfEOLOZQby0xVm3TvrfaFZHSzyU7pjjiTjmE9lrjjIt
CbGCKGurxLzMn6QS/q3Bo/dGmKh9ICu+JvIYif2sbuc9D7pzi53Dk2tSSXy/Ii9zFbHwmoDtygZC
zsQhljpHd0jDjFyXBoZIejb8/U4QuRxg7YdeuxnBBHU4XmOKnvfpSE2AMcGsBYuB71ccRSp1MpnX
5od3fD2Yi5zVyf8hIBVfrXw/SdFUcEb9AZQ1sTG5Z9EdEf691H/fBe4hA/5KBFTzITJijaloOURL
PSAL4BkCf4BHGpFG/tDQkZMPfdqvPAdgyoDYTE/FuBxJWG4eRot7ie6goRW2mQz7Vs7gbpu9fGrk
LvTvoQmSMeSsjc8jgLqN22Wgk/uO1EAOyJRsbRHq12ixj7yVDKTBf/EGXC0mulicP8BOn7P7kb2R
ok/9N9iBF2nOjIWYPGq+nQscGjaMLAaFOLjthhYPZ4NsifhRX99NzIFQCnBNbgMM0s0EzFkaWXAS
cO5weCXJH+FaQFcbNBdlcq13ktwA2KF3DlyXb6sKg4sqtO2qyX9QN1PMivs3Xmaxo0c6VJHs8iba
ZoYrTqvlBerQmUENJsFXT9+X4lJisKHFsYzjSmjCkq7JSjVzTPzewz1f1B4oDIuSB23Ghj8z0xKI
iKL+6ctVofZDuDIN0B+r83uprxN76gCRSpfTUrEL0d0Z7rIm6+TX/wBBV443HfYAtTvn1QhdZBAX
fhWtH1p7skr00BuPspaqFCvxO6q5ornK1kKtR0J9+TEO5jTfaCzFmS5v9LYI+Ps9+ReS7a8KYdue
biAkFgEPDWWNKf4qUUJJAdd9YSlq8xwqps/JkHgZwhBFLA+GcjPKfE+gRjCJwDDg26BcASotS5I/
jsfpQAabmY7YtTbMIo+7xw1L1Aq7o+fxr4MtbBC65V5YPpzWoDcVM27EX18y+dZkbVZtUsYICQ1n
aDtfgxn9IO/tbAeDh/ZFljaUI8EIqyKtH8nha1oVRF+dFEfbZQYMqq6QStbVox2tAOSHeQEvUEvn
us4xBlJbhP0WQLDG6svnsN2ORHDqOn4B3vL/BqGJ/HwxD3cuAqGYOjI3fbSNlbwits5yFxAMoAsz
4q4orqtEpOnGZivwyq6zKaAVehKRfuSpAUSr+Q7UhjIyWsvrz+4svWP1tFGV65y4jTbUV/MraKYE
ghwA39nx9V0SJeK/6p1lt9z1kYXgoe6LnyU7RH8/U4bB0vVte+EtIYswBYMAZjiWU2RVegtbpljF
LoJ6Y51ONrK1e3dJpaTz14jcSyCmf3oeMZZLhuWyoSAl0/s/fLl658t4+As1W+yUQmWiQXbTRe+3
uvmabibDG1Zn3afLn/1scNR0EYH8jSAlQv6wUNJ0JM0cFQ0zeirsRW5GYu9TphzLHj0jh/sM/qyc
O9T+FJf8IslYEjASFRzvSrMa4hHtioFoECjbSqHUdCjXj1hPbbpjm0duY1016KsKfqEHTMLsAlpY
kFyPPLTJciyUNHdgVarkxPsuuYUj6o1v7Lrboa2wzWUtsQZgBl5L37n7SQ5xUrYQlN2nJCEmKJfr
Hoqccg/NDloqzdGGXr+wBtu5tHVrQ1Uf7M+4o2ruRfZzGThg53RKfbBACX8KgytSR4yKVWnzWGXP
7Ekp+7/IrQEVHwkRqh9lFVZ8jrV+HW6AVYhEujr3AVXoPbJXhPhkWezGlKHb9bQDbKd50YXRp/zz
n/AMvE8+2TfjTUGjrjKCOooTibiRmYKLyVStDzFECSjU1OtNvqIuO/b71XyiNJXExAt2f7/Qi6rJ
4yX9Cko1TL8QII5JmTmxaA2ZQJH//n8SL4XuEelRH8xKAqmKl+fuHQw0z3NEp9ogIgfgZO1K13Bv
yy30WGfaCnR2QLOgLQTaqFTfXOQBfbUNK1lrkPGf1aYpT9KmOEz8J7DOZM8e6x/3q+Bk6KlN50d9
MzK+vY+cXzxhVUxGeBfBmbpMsT1qNPkgUrp/fsvqQOHq/YDkjB3/ayDWQsXh9+RdzyAeClLMFyzM
Ylnqip/BjlxwpAkGGw+K8Dg1WmZy1j99Q8W3SJc3VjZfEyxBSLPIDXAAWep2r+YNYkfWdtf3Tq6q
kRkTQbbUFLydCNPkpwkJ3zFZiuODA/OHHDm3bQOhNFx80avQQcNZZLBwlsoIZ5JTaj/kXuFiyFVp
3bV8g/pNvG3YPTLaZfPXPw4D19p+c3miMX8R8emFhod3ZISSWnr9J9PxJTblF9DVK3vvS1jmQ7y/
x+wJAQ882G9uwoh8zem6pjVZiZk7MUCY1GP0DreOlGRUAOc/gdrY3x5QXfciouGlonW8FIn7YkwE
W0XA4NK5O+vzmWWyB0RGf2mwr3KFdLoWUA7gWxM4LbaT5tfiq4s2/eb4hxlPnzF+yGjNw8QHWp4p
uuDVFm5MsSybejN2/7UjtKRZblVd56ngibRLj8NRm3hPbR7bnazVeYzLpyasrda1nkdy6O4hNNK8
GYpMzMYv3hqucPAE9gtrUJ5+c/H6b+ugS7LJLwNZADqLrL4AlSEzhIBwgwQytRVWQB1pUMy3DuZO
R1c/cpuR7ik21Fj4HC30p9U4ONd7q5dE/VAT8xiawscghakNk07QmWQHNMs2z8zFk0lOK1QK7JtP
VcC6c1mnHsvZkL2Wh4eqpQZz+pZP8uaIZEWNV4P0CcRS/sNpvJF+VcWGsaI1DAR/IgEhUGaKqqi7
yKlUHG+qdKmnMM6XDiOGMUW/JI0RlgHceM0LlestbcxYv1Y0j8qHjGjkrZ/8r4ATNZxVExNvDsbR
vho30wNdq/nZTR2Sf4E7LBdZIxhr4t//9561lFjdYCuy5kol8WwMu6pyZkVZ8zCqKFsNjzXa9A0z
oTQCIXStji3wHsB4iO9qKv2NgeqU0EqXMK7apWewVa0rsbbigQ1viQUEdQ0bzJNAoxHzvqprN2aK
kFA/eK3Res+smYEjeRv+oq1wk4Q7p12P3xohJW+I6AKbo20pkzXzq0KLGpY1/xeAdR4G/nSS+BVT
PZhJdyQJRw7jjoP+7M/6MMQ+jgEKos5IXBTZEBJdtDd0+idTTL7QaOCvCjcs9ZVQW3nTR9P33rS/
PyGADfDdh8ba+h7nfbLuxF8Vbyx7xcM1DFpxj+FVmWFqfeCg3tIuor+4/IJM1cDG+5XQ4nZJ/RWO
kW20x86YIc5JpW7JOqnp76Sml6hGAj2lSqh9IQPl7Y32qhW+ME+pfUvqZfJElPFPA0Ta0GhKGkS2
dI7n51bWgutoBDWYT1BV5TlKEC1NwB0zYMhHb/PvrlCJHjjfH0SDiEWcAkhtTjw4RD3VHB8r8pKZ
cOWtFfGY01bbK5BixVjuVeesf52phKcWN5lM9fcGWsxVbluYMhxs/ujDwRlKfXohuriA2LzNcEl9
xLWxE2vV26XAp/KevaqPCQvkRDl+OLK5LXDoixvE2Vje275v6B1eyU6smtfux0SP6o/fXbKlSeay
q4VWOgW+tlt6Y3tZwAROzJjX2cXpd7RM23UC+oBC5hoy/428O/NAyfcP13R0tcL3FjlfU96jHan7
mO8iiNSsPHgoM1zTnrAj1eHBJ/xMml0E0vpnw05+hfpxMvtbpNbXdj+FKEI5jrZ+rAqCnfcnFNbP
lZRoIF91F3oZaD30C3vNCle9hFCl+oRfpVuamnxR3lh2/7vMW3Yi+lDyTpJO4w33IhTVF9XjgEtW
ECxGPdFg/Lp6Y+Su3PBcQrZc+NX4tnq/xYZaKhVp/MLEP4Exb+w8MdjtTADtHvFPLiBtkELC9BMu
Zyk4lyiJmyhu01tdwPYcHigAiAZMV9pUrNy8E/z7ilzvTGtQFh9KrMKzPcPfKhq9Da/CV/iTTrJc
8HLFam8XS8xeBJ9mdKFvn8AkGWSbbAQHjgmDdvL1AkNrTjqwp8tGt7FwgPY2+W3j5TGB9BIqZ+XH
EwSxZtGML/yACNF0s/UM3XQj5pshAgAgV9/Wl/LZBZa4+8Z/2SyJermx/Q6TVZijG9q4UXz9hDMN
S10WYKkMMcgOgiF9dgiixaeAwkwBMfrtB84l8Fr85zbj/KgnvkLhUXOZ0FEZQApx6V334a2y8IYQ
iLXX9MHCTgPVpmKUA4OuM7yuOmj8AMqTeUmI7936bXUBbeVTikm0VcTiSCUC5VnU6GFAPjdc4xXT
MEpsdyniR4MPg5WiSuLST9yiyGtgrG6xxp0U1tkq+gfRXlQCVg/i696PmAokCOzauIFQBsbePB2s
U7usMO9YjPIpdIqKqkjsIvFnUnk4G3/Ru3XTnLlNHeERMd2rStNFDwooEBBAs3XPlU2M7MDpKYvw
1sYJGeMH1jLbh/J1UocUuziF3VVqItR4/PsONwoP2UxF1gkg8YpEgDJtjWwnP/2plJ3NaCSfAfdE
MZl7kGPfmzCvlvplyVFpUUzh7j9fb9+bM8u5is4A2MwjnYpFOpqrDereikgeO31xhjMOun1tcEUF
IQq5tagO33T61itZpnrlg3+SNCNJDt8ttgbN4zF91raZOSSznkUhBJ1cf0yYhwxBDoPd97UAGWN8
qP5yDOfybPqW861mQrZiqLZSAHSR9B2JmYMACoa8bbuT7LsecrbOY78tioXvgVNQPqUpys/mIoIM
2e/muW2paoRmP/dp4cn2OTupy0kwzuv+08bmEiSgBlylDd0dcyFnWQh02pBjw2yknqnlIWNJe/N5
+NIzmLGeMU+fBkErEPd66gnUvlfpGgfrhGxs5BNonwO5+eDxXN3H02ibBHtMWmlR37UX5+kI4WBq
Lq9A/rhH8nsEsZ4CTwh9dJj0kaEIdaC0rfsCj1DyJS1SN1sN8mt1XqyfNP7DCD7rHR4sVaoku4vc
37P1pKZkAqUle5ZGihBkDDSttFper43AnoHC7u82B6f+XUbBenUKHnkAoJTtJ1JtIE1qcv9PM8pv
0uNrb3EVwud+htJtyNvRfFn0j+gyIYxhD9Rx9/boZOS5VBZpJiBo08cAn7oTVJNFwhS7tq6MfQPs
SoH7mWUK20AZYoXiJIh6Wm/od9Q5hzZwkOM9YTHBXlplLxHpyi21IldYZEC7Jx4GkfmjdIIY09vs
piwYAaxpI9rriiise+XQqFg+YdNTwDmaw5vo7SAF/6fX/R0WdoqueOvQIsKqfUsykR5O0v5iJr7V
oS1wZdfYP6Fis62Y52TC1nx3AaBK32sn6mLdTZ/JspybbQ1yrlPH+SH7bZA9hMFkgLpO1rxEMjTF
eAPFG5MbS4V7FHf1BOODhAOIaPI/LsG3ywkmagV0QeP5aWlNLOHnMnTbzugo89B5DF/23yUMTzOn
F8t1CjCas/+U8l0j0HDXR1jIFccm8x+fSzzUEtRqg+konaR4Vqz/fTEa482ir29Nrx7AxmITn53G
MHj7CyQlAaICmTZo2AfD4y3kx6xsznTepqSEk8r0lIaWehx2xf7YVWwCrKG9Qx9WsZoB3o3AAJjt
nJr4MEUouzQvg5ZFy2+7nxYoNUvUIxkv7zAbqtc+2Eb+ux7u70ARrtuMUVOOCwqm1UVCEbcXf/aC
HBVhtskBIsskPiMLiO5xK1j3yvYJJOoP0cS7qJ2FgWi5g3Ql2VsPtagC2awTjx+o3L0IG2EJRJq+
mgaci9NMfqNoCiFVIym3p0vpkHnfQhPkEHnT/JtxopYK0E2ki7lkdtH5l41aEgz78Tr/iG3qSetm
tKXrbRgMssYFYgONyB4+WSX0g1UJ+PoQWe/K/EShW/XjTCfAWtYFqYFExC1bA8YvTl72cHC9eAFq
hh9ARX010xCP4LPLhMkGVn71tftFAOkV03QCxmhB189HpK8tyhTHNZMooFfR1eBrVY4Dssp1G34W
b77S2+lp1KdeiGoDnedJjxBCa+omgkagq1+RjEfYiw8TiQyJld8bb96TYaDT5wRnLyz1ezjvSiXO
rQvW/VRnyh1IxnFftplSCUVzQn8wRXyviYuV/TrU9aB/7Qp+tK50FtXiaate9F3NMsXbsKSqsO+F
e5b2bcN62/hFthgF5d9Htg4t6e3HTGaiXWlQxj04iJpbo8uoaJgq6X5eoooCwFaLkLaDzSqAmoHb
g5QJGotrKutwsHqK/FArnyA0ELRkfpAo10xxecoj5p4m26hP3s+vl03fk5H9YGS3VR8arxI1tRPk
rGtautLYewyoMgNxdUp5zzBw+2Q3QQGny2yVkELGA6P2VNKrchirEBRcwXVS1XvgioLvL2ND3tH8
m2FoFKAJaepSr0O3DyS67uc2Ji/8pOkUdUv4ggwkKDtp80YsDHuvFgRmy39OY5uFy/5Ov72lRCXz
PQm8HHtDgGoyOPUfieU0AfBbcyetK71ULicp9AeHlVa+F3wzjYVZ/aXfLNmXwLQYHWCTxgkYwpLD
9iibRHl7x5rnEB7QsagSoFhnz93gTWWN1cPDXAKe28pQX7sLBlROZbZT4ZbQhINJPHRA7eouIjjj
Zl3m41ZnTgyw3S3qVLTFdgywA98qjhVHl2lLzbxfwtvN+O/OUF7/kYF/HHuxw1EW5ai+i/K4WYff
+igg1bY2hSru7HHKctJ2lv5GX9RZPsdRC1VuNQhq4gPK+DVjbHSdDKWvCXlps3EdNclGwk+Kq7fk
2BRmHcTxztBbzd4zaDOUeTCsYrLK3pYGEPdY8xJqqwX+uxMuKgulcnTsC/8TI4edIFUAtSZxFAo/
fx4QbdIyjnS3qGPqhdOI4axv8jw+whrK+PHE9E/ef1GpoW/lVns23S2EPpjFE015hj/EJHq6/eHG
3DO+6g9sk8w0JJWCbZCIOSmFe5TaMb/OmM3Yo2zDpyO/UR48z9EspPkD3wySfE3QYGZOTS2jBDje
LB7/dF3Ia/0sWPgj36mCGRJu23chn05KeTD41aafsk3KvDkBtysFGZAnTcoJnekrwIepKHJdiWJL
43JiY2iXAOsKyxYiMkoV6SNJhpbr5yVgiV8br6VibfZ1cnnx1ZRT+EPYAIzIk2w4QNasv2lWswbo
K0lQ3eFbqffnuxs+l7PY85Z7NZ1rmydzu7yPDh7rG7yqw6kTTRSZVUSN5pdg0t2NhoSAF/xYK4E1
7FG0g9mjBcIvJW+l7mk53wEJ9Bir6scq4pR/5EW9EDve2kxU67hY3Q+OOVAfSOaQlMzrPcHApYPR
B3IvYaPIYXA4WfIQy1zoOAbCq7Z311+/sbdD+LBAoYf4xEQX/RXCzV2zOSsGNGPNtGzLVHVIGhtl
7N7QPgMfLQmiq/QNJqd5GE+hvKHAETxi3wNKFjTN5ONWLFJCosDELRo/aOKxjDn138rBVKCSxTyv
vYLhX1KCn2766vBibCaVFjVMA9ua4ecbBDtk2fwF/xYFC1ch6AJT1YqyNqL1nMZTW21KaYVJG18z
D144QWOB+Yw1yNQUy6l9VMmvhAF40VtfKSobN3qkK7/9LZ2+OKNUXTD8/Xf1uJ7YFdg+5bE/uC/V
ODaDSoPjJBRD4NLMhQ6/OfEpPFaq46QiXh6HbO5KeVWgZJaZoe9iNM7b41ftoTcIRsjhYr+M+zXR
w14UlzQRUC7zs3qj80nDkRHR7fhC9T3eCLvcAW7pV7y2hCBBsbRwo0qiyAAQz2+ZCG1YFmfmTr3o
yDS3fDpNyyeAYP8YiZ6KJsMFUc+cje9bA10tQLHOX/srKln83N0EmsPA4Wt5OfQkFGYVh9UgjUbY
qI6wPDISLPUOtd56+srEaKcptSgLzpfphIPIKdx8VO8BF8hFapdRqGNzpHcIWIk1HWmvprYTnPnx
Cks3MNttxVGekohO8WwIceWnXq54cU4TdWgWfzerT/PzLkINMQ8CdbmTr0RZ2Atg/EpHgKZPvtNQ
DZFhyUW+oyOIfzws7w6lODYHFErzjm+zwD+XBR1HDA0N8z1Da+QXjrJU9M46h1lqI/JHKpHDLmil
9ASqELwxnhOQkfbr3XSesANfwNqJnA5zzD8kwvwNE1hBDq9UlZiM7mvXXCSwuCdzpl+DBOGhSi5I
EokqdfEYeWP7pjxX4GteFSbaCNyL3oDmhFfhvBvPY04AYHPO6VreBsu0/tGlrhmxjENXQxMygRhM
f2EfbK3sqmWifA3vtjkvB9aJi6JKl8IIAjln7xJxApWZ3jcAVgTO83rsErrnszGrCPDRMcqvo0RX
CiIYoa3pdEfQiDMTO0gTAsvzlLmsqgfy6sEVxBbQyKGQE3hIr13WUKuC7z3iX4z9IRFmf6PGMSfI
xJ9jJSldkn9b/cXJ0+ca/tUbH4kYfr5vENoAjEBZE8j3oCrj5m1E+yQP37JKITFsNfxDL/rKC6eR
amtQwi26N8crBeKvYq2YEvOTev+VtWOrvx2ABK4xxdSeoLZXi9iC2CRtzQXzEiKsruMQ1Dxx3Rr+
MqthJeed9soc3pK+GfxIAghiAYXculRiaSYgTWsN1hLsYPQ6MAOrjKfHZ7FiyA4ko/aFQw2xVb+j
XGzq7CQdPGQDfMouz2bor0/O/cdb24GsqlCd44HIUBeK8XyteyIDpr2yhI1YryIj8kuaJPxuhTnb
U4zUeWtRo2/RkYRDG6HC61KeCsbdyluVSPNxhbCKXdz2OfkAyfUc1kIJeIpu9cRWOJ+uW0uyi6HU
VXrEXz8MFOyWYnz7iXrYVXCoDiupHPnsliRyC4Aqc9SQWq4yrR9PQD3UH5ACZoDWROvHw/jSC6no
1T5R13XGUd8bxanB+cwoBzQTxSFWP70/uSoTWEFP1I2+JH+8B8Ou07dmJHLN3a0ZMXzgUTDTX3Ju
jUHi52q6EYsa/GLJMTVcmHwZCq6b7cZYfbZCGq6m+ffRGUUeJqRyVNzk69su+Gf+f/NzKjN/3f4s
pjLqBW8zxIuIdZWUFhYrZrqp5AF6VU/SKEs2Dhdrx4fpq3iU7GI2t4k+kaDyV3JyUBJEyvMlvLA9
VPmEtNe7uUctemnzn8gsj117eOO1KBahhRdGf0H0fare6JTlafV7mvtN9jv/LAU3bEPDY5wunG3l
UQoNVdLiC3PPsTQ9zafRGB9QhA8mRU5cuzNJVRbiidNNNuX/x4fplr2FUs/Y+tOkpk+HvhGSKk1+
To2SVY3JaXV/Hl1LL6qg595EnW7C2UMvYeL5JHCUdWal5AAbGx6kCK8vBtxuMxDKtioa0wDFjq0B
/i5zPxbNxIOFIj1dCq2UTL5oPu2NhBIiXgmhVmwEV1gItSup/KD9bGu4LnRFY5xx6ChN1Oe7FRhS
OLq9r4k3rpjl5CuYR6W/LjAVFiZHCVgPlr/ZBjDL7FgmJ5PwfWwwQYNuIxq1pLBqstQ24u35Xh4A
TyJptHAIjyVoOEasW8ho66EvKL+UUvUNyHEcpzQsMe4oizPeMQXA7EunWF5lBqlSAUWbkZefiR0e
Trev3GrcJKFFpG/JlO0gZhDTbZ0wixdy89hwYk/qj18LNJzG3c92Zy81Znm/ytxArvItA7nPmopw
wFexoeXEt4JfbMem7Zjn/kOLIisnpp1yklEjFBHyDUk13qSjszK1TpygpzCXN8/dPnsNMKZQ2BBB
9KkkYMipADFdiG6AtjFMknzE9jYf8619GN2PIVZeNKdOk3PMCOHeyskmE+Hb/zdi4mHmGZ8r497z
J4XuwziD1/8JIcs212GQVbLkgmu30fe3kB6XYRK7kxxvfxh6NSTb1qDwsuWcAPUD2LVjk6egmxIm
oqrvuRw34FqAhv0TG5VMvQg/fuQDeV/0KI9Uo5+QHgc4mK5u2VeNflQedjRWw0DqyzxO9cEp8SGm
HZ8w9KDtyuwH2dnqm1RuZyHx9SW/tleXxfZpIQRDWjSE6U/XPgUEHfPkQcEWUnnJ8D84v42ZYc91
mb3iA5f7J1OC9645kcY7O4juv6bI8nDbYP0zMwmOQuS8EgUfFxude4b9kMAOZciYIZIRa58W8mJ5
wOCjJ2HcSYO9/2jsjKQFe1hN0Ok3Jx1boyRpj5cQLcZGiY61AkyTNXelPvtTeAkBiBhT2ovVEdsf
D2e4c7yRJE0J7SYJvNUipq+XupGQPMcZNQZOwLaRFR6L5AxLCqDPw4+PsF0DmQSXqemGvqsCLP5d
aHg0lAa/Hjcdo7f0wRd2SF7DSAmkXn/+v5RkGatHiE5bv8KeQ7A9jJf6qLSOAq4qoK2iK08hQQPL
/rzh2pSAqplFZTmAop6vjreFDZbDl+KHC5qUJscf1+deCanFVsLbDDG5pxJ7Le/RcBS/SGXF1ezW
Hy2QEPGrvM5rHZjt16y1RgA1sUAfUAh62/qrjFgdvr6Cspp3CpyCfJq2oGISUdYJBcdToC7lZBXw
U54jrgKs+NKMUgSbs9o7rM4PC5sVUxHWT6Kd+4Irri4mBGHx6jqFu3rJFvMwDC9lOu0fI6skYuNF
RMdbKGQ0rDZhXJQMnCPTbX61V4GK+TW34EXbRzMifh/dhXv8GOSlcpnRHiEZ0YcoDEb8ywr/UMgI
uU8cxjRG/3RoCdli3dWXCg7+ara2JioW86DQV1xbNXaRTQc8b8T6NaQO3niZKDv/fvUAgIct9sVg
RSGNTAd2YGZDPPce1pWqga7PXtkhaWnLBr9SC7b4oZqZxxbkvuhAnkMdTN7j/FvoyQGfHrp7WiKP
jfG/IS3Nv8fus9uuWCZJYeTNAMF2pQyPGqW+tEV6+PQETespecHU009cgH2lUjRYjGDNggvj+1CG
43m2fRjxERBAsuuKdh1AvthW/16KrWgxOGFdRGP0if874rMjl4NKmzDuSyC/HnA1TI6KcWsTrlHG
3mx0qqWVi5/7N3c71DjJosGITpDbk048asnU/jiQvLykyPJZyHAPyHJFnpLKNKFx6l0J2M3eSuTm
bzVk6B0VZbtOUQ/fcggT4kqx4CdBJqH1AQ05oYEhATpqhdHGocDkuUUQii3bBT9afIfNh05aZrac
M5rUoQjztr2ltQXk3KamRe3hvHRRn1eJqc3u/F+6I/SoZvJk16NO8hNcgK1P2OCxcVK/Y+BdTIIW
mbDdFTrWDF+F2i3iDpIIB7MtHyXZDwR48UiUmgXkJw4ngsabrs4s7Rs+7meRon1taYuIAeJRo8h5
ppXo0T1tuNsm6gwgQY5W1gCqVDZTCER3d3CNd2e2EY5VJudaR1W4ph3eA/55Qo5E5H1FQDpqgmFN
GZrosEiY2BHuGDCLUpsCjaALpMoT6vAbug7eE+PBuUzLWqFQl3Eq8UceLzeC1X/9Y4zxew/9ZTFp
YhKSMIjksR9hIq5Gf0o1s5cLNpUm2kLa81L6cO1BKAVfLaU9KN6GL42rn5+TJX5ot8NI1JKolAFc
t2eSy17S+ESzK5oqLVGrV6D376++VZnxPZGA6R+h7ed0N8qco5X/JFkoE3Sld6Y6uO8xAJfH3+5Q
hWciqkL/8+n4/sC8VCp1i3fw0w8CKrcle4u0/Dp2Pp+jj19+fY1KBepTI0r31yCX6yYJk9Xtp1B1
7D8PH3XnZDile2X23XpUZpu6bt4WhyyHDbGKeGSAqWF1aJjrRLjwrRfIIBD+7YOjYRLpusnNCZPt
QbU91+8fFfcEeRGubt7voKF4l3e9k7bsHBX7A4/zFBtfSWM/GzIifkSe4RGH7Xayak6JhfyjK6O/
wMbEq5yqjyAglI3O/Yk0zzDFj/iqu7x9CwjS8rmgFqnP1rStetdYE/K8NWFwId62/h6X5OtcJOlE
t8veW8GSQaIfAjSrlITqBb7c3hVVxDzzEmY8YfyV+/N5jC0PSrpWcXgUzNCkBOcJj0WghGs9UcPJ
vR7kcw/JkVy75wt2+lQSvc37a3wy+G6aA+U2UEFF44BFTVBK8Kpmje2rOpzK2Z80IjDE8mqlwGYR
qA/3fFgWK+nK/EV92H6UR3vLZNRrmoONiUNOb0lxsIZ5EYTjzKi3mwhHQODJpa4o5AyN0u2QhunP
amdab1hkN0fOkPCR9FZllbxSzBHnj87LYdOEpgPnVbVpqd5R0behi+ArH/ONDk1B/lU1XfVVu8bz
97qhGif52tUifGkCdPC7IP6RoiQUHmTv72cz3utJBacwMjysNKrqrj7OGcD0pPTuZD1+7LIX8Y4H
vKyBsqwJ+I4q3L4Ha4JJXNSvKCnTzyMY3B3llZ5bdGsCocFXRNaM2PvstEz7Jksndgk/M6tCHg4V
t5qQeL1rs/I0hfA8OddLlBWivJytDuQGLtDewL8BEHqoc5x8lTsyIto9MWPrggZUezSpvJ85qaDO
JiXHN+gjAWhNNKVMxgxAPA8s0mnRXMMqqHzfNRiVQRnK5ra33oyPn5wdgLZFhSmVZbIUsoLl9Ekg
a11uqQJ9p36n4+UeM7v0J29JN7bXpBvwmDgBhGEyfgH9psMYDpjl60KlZlMQQ8cqtaPtorwMX1S9
s7TdMBsm6DQ3fdQFEsQv9pJUg4lzkvjFqTSEgmRX2GhE0Tl5W3qfEGAxXA2wE0aUJNPETgQnyczV
coRxx9tCHjQbqT5ggk+NkvydIKdm7piBLm0XoyV8P+2AnniuMfoEWCWj2WbjVyhPxzOSgIal8TGb
wVGZVE29zgoHyF7fp3qRkv0Hg+tideTo2FM0ClfBHotKhtT6FWDVjFq4JCpfBWyQsqWywZ0r6Lj+
jlx9RvQkiBkKfZOPocOCnEQFkEOP4OicJAPViRhmL5fkqWQxZSIeW69eCaxk7o2P481Ydtfb2aEe
NQis/9JpdTN8/+J1CJ4os5vFOynOHHZnVYY8JqKV+AyKtucDt0Ebkmp9wrYVJRH54F+XqBxkP+yU
jyIpuUMliDDxknlDELFrfbfWUSRTreEGgFcLYcurjPKi0YqqoQNRfmCXw8QsOqja5wXtzg3QDLM2
5eRPj/5om2tiZmTBxQi8KlBMxFreOVt6WE+mE0FEzlHj1TBytnGyFGAiTqhtn3D0IACx6SD5tYML
6gaNDSXFTnoNg0zAsiG1i/Er3Fyh0W3OuS2M92piB/PrunJR36EL74CPmctbJDv74SKlSX2hHppg
cslgqUkHG5uK3YT+ZgcvHUsViocv68DazpatMmyskRSpyecq07y/Ctk7yVNYo8oWzpJjM5m4n+9j
kCvtm5Cq4UOAVz4iL2n748m6I/qipE+SFel5EZsgJBf8gszVmiScB42VW9S9XgHNJOq7GiqMBK9E
qFOxKMz4R+UnwmFeo7yCqqvyPFusMooNZIcegI0TCFWvTsbfnK+sZtyInelttH+r0jymA07IkFUk
jPOskpeudrEvlruKy3JAGBO7Cb2MAxDZS2Sne7DD+HqSFTk/wlQCtNj5lIbvXgNH1napdxYJ55wP
L++SKeuBZVci7gL9o1rZkMIoC+jbffB1sCGVXXftMYkMDchbqXRzlUTgBXJE8V+fsqFBY3rhdiRU
pcV1gWw9DT0UbVEezIWWfjx39Ntr37ULpSDuyUCXQglubklRBEpiJ7FdBPTraBTlIX0WtDQzWuW6
FAsyHPeDRmM3f2uRZfm3u3S1ptMyNXrno9jt9abnUQryigvaAPGpBl4KVy7CCRu3a5t7PH/yyO8y
5JKDGJ25PrDj8ejZZ+E2g7C9BmUvD7P+kONsFftH9E08yH7laz9SWyPpolqfvdkCBQC1bSUhqF1G
nGcOeBdljTXrxY5Vau+P6EZvPTcVxxAXovfVXgRxP+obP/rsoGMPKRkHeSvVpmMW0u2hKtKYQw7q
F6mt0DtlbcvUxR4IoMXYwZ6pXPRkOL9/yav37fsN0cMjAw8bMCorKoO7mHLdwQF/XbSIu8Lje77b
CmZy0C9i+FRyWJAR21UAEzucpTFDPAPC30uR3gvw76eNhW/gQ+b3GT5oDdQnNENLbAG2+pzNyhjF
Bomxs5dYEIEbEIGqNMZU9OMIS72P2mWdN1bkpKejGBIhOHsxoA8SeLVziqiKGLF/ltfQ/kNQ2H/+
qzzyodM/LskgNStkJ9Ja6e4YajkOolN8K1nr9v19z//1/EEXu7nHDYQ3WsNMybO91KKWArrpSqWV
2QL3xf412LH3EPEa9V3NqfG6nvVvKpYz4NaJA/SIETzYLnzgeUG+dzLb8tPe3dUBJmq5l53lkPZZ
tweqmNfqpfcaRTuJk4GmOeMNSmERltJ38nwKs5G95WBJe575OhMPyvPhv/YvjhO0mcGK+vwO2JeT
OemvnJUJmHNixIKLDtiCTpDU1SRIAOVXs44t+VPVO6dP9hu3EjdqZz/iatKkjctYys4dlNh27aKM
Jx/gCp3eAkrrRcP/fCV/eCHSzfdQ5niILPnO7NagKcXgcD5rbeJvyebGJ6BRYRelk14z+wEZh3tz
clF5RYIlPIvn9GjezrT2X5aWP1ObDsV+FKSNAbYR2xPRbOBGstw9Kyq786DErOJJYcQ6Zu3Lqx3R
SztPvwjvQN8vm0u8/TBZPt5hOdD17vW7QDNG3VF8ZD+FY03DsSh/8qFpB9LCpk5yuX9k+9GP1UlO
SrqnhhUC1J6etVrOW7UGHZLd+3xNy5WYqMDstyeMBKOkM+X3DvRN81gPOiOIZGXtPlvtc0nHX3tM
54NmaKVRTwPb8W2bbYPGVcN51H84E4v2Y8vunmaA1Bsj3rGEwLSsk2aHzgrNchBt/5B34U4/uiUY
vjTnNebtVTGUvHksO9vGtSCn0MBmcFWFVhTI93kop19FsMA+gYeRkw3/EUbt9Udyuc6zTPPs39kU
L1DzbEdI0MTaQUsRBL9TR15nUe22rVQjD/thk7MTbmRLERcFFsb8C9nl/YMhgfUSAwbylI+9C47e
I7LRtSMjfGoc/60A6KPQfTf0HB2QCY97NOhkBLk+wBpEqO18n0d+TNAWMxqla1t3X1JxMzHmjT5i
QtVEQ52vLMIj0yTnV5NGcTSnkrgpRDYi6bYZb5PsqOaSp7kdylQsdHzSM2i6eQ4LY4QuoNLfNQQv
xZc3cTHpkbhavfZcJy8aJgAbg/qIcuZMnZE/yzQ5U8xgnKymcC9gIbW5Hu2hhC9ftyvgiIxHYDKZ
GXLWSKtgLNeRtlfEhsIXhjun7qd6eEwY+JCYsM4u1vQj8M0DWp3ykJ/8bMnRKmykq57YqUSY0MLR
d4+eaVDmN7iaZz3p8wQ9tIXWOhRK/m4dXUcsV2dUoWG1w3GhHHgwhGKYH7kFaE6DYY/IL+R6Sff6
wqvkHFFJDnBUTBRgHfDGs2jFVHNTlobdY225RzJ+50crzRvFqUerhfQNlb3PbpEPC3xXxTJsn1h6
PvkKlc75TQUgsyIwSARM8UJflRrBtTbGAiv9rIxEvryCw0i057i8h4D1tDjr83Ell3gDqFj4zaJ1
6Slyo9GsNeNMxOcCXJAfyYEOaNwgJ4gplOPTvarYbraYqf4nmNaCFiQ241BvzvF6Pz9xY0z5EF3e
Lsg4ioBMHchQOGgV8CYUCWgdlA0p+R9L/BUxQoAP3GmgEM0Q8qT8gwhFx9GWtyHJRPibOnocdjcm
ojLAs8wpqNAf7//+r5lfR7HQF42SFpmetn+YW0XQYv/axmYSsJ2D4Idafe8VhcGK3cOMuBiETImA
Q1bt7G9x5Rjr+Yr+986zW7fnMoVvAS2mzY+pQMI+DG489IZVRo5XNs1Crln+VXkeYhTVb4GT1W6R
Wdn7UC2+BU0fEEmeKUe9znUcYg7Xsflm0yPEtGiTPv3bEn3cppW85P1nRNazbLjdk+ED418P3RiR
tNNY6YBMHkyA3jNjJg778QCHopAeHCbWniDrcM97uqq9NhPck9J+yuqBIgJatwrBEDQt/ygKwQRC
bLh/3FRy0CQ3BQTsT6AAge6ImwUxgtbHaX0mnVicA9DdT5c+hG9ApFaJ/c6MZZc9VcmUDPpP/k9p
HxLnB+x0deZDeTnLFBFNWSqfOLRX4MF9ILgWjWru6v7wqm37Tpzs012hge0jmlVgkQGToSHwgrbR
vQT0m5pVgiZsOvEyEWHYSh3kfgWpyCbxUmnR9nLhkHuRpbclT/mxmn11eDL/1IBEq2WKRN4J07PY
2nLj017mcTAHBVfXpv19NUT+d6cI7eAhEGhKdojVrlVmNBC83t8iqOT5Fr9WL7IhcIE8hh4T3tlY
AeUqYl1hshwLxp8zovY7IBjlnlO0oCV/RK6T0L/jnL7U4KxVmLQ7Fa3JUheDbYAZR7r972uUixpl
PN45AmjCQkt3NCw3/TZ4NnUnEnS0HnOgpfnBM/Gwhivsjj7kewntnpB5lOLYKgZQW7l2l5//9QzX
hCalwkPasUtCZRHwwqazuLgJrdCF1eoc8/nXUjXpuR8u39sfhLlZTRB4K+nt7QuQwwBr9/zE/4+A
7xVQmY/fF4qazbDYML4oauNcykPhC5S9UpZLMfPqWiZT7cU79J6Q5gb9Ee5lW2BNI3mQf/TvNh30
Azg6cZu86mw5/dZHJDvPzYTdIfxOkjStOs3SI/MPDzqhqlvZHPsGXXTXphSAtl6fPPgPh40QA2mJ
JFgx0rYzXDwIZkWyIfOxKITGSevHIY/iTf7Gq9nAadWFq9E6hIdjA+LGlJGfgEv/QiVWx/YOqTWT
Ehlf4BRIRp3foeOri7F+P+XqArg+uFO3eK9eSKl/YUQiwK4UL2KYRpY0faDIW2nRsESy+gK/K5Ml
qm7aLzc2dOsTze14XXQVNm2jFAXG2QTAscmUNlc9zFYsCmXDJvLUlbFqIBLK0YYhehjK4qQg74UW
EsmABsc63QlcSQPnoKRm9fBTnN+pQxuVgjQ4vBKeL5GCdI8Lg09eiw4yKnXLo0poPeVmFBlLwm4k
vs42LMfZ8N5HffC/e4gvbeK0BaTPReJyGTktyzhC6bz1w8gRf3nU3INNQgI+K9c47tPlcvzU09GC
6E+4sD6U01peokz8TPdAlfuR0Kud6/ZTTKu7feD8fmo4KR5pgrBxRYT6tfIQZDQvLE6ot5Ls4R/O
bkmuIyurYXBHFbYFUaMExigvmFwjfB2YA8pks6DVAvWHtLp8Ap67rKL38OP4QG9DXARo/B4u9JDt
qW9qEGlOooeTSDqwOVILK80XBQ9IfrrVjqD0EJhn4//DicLscUOrf2ukU8LJoGzopxHuzK5VKttb
6u7Uu9DZeV/PMD6k//jgmC6/u6j515XRqFvObHpGLGj5x/oINuZNsrazC4YCdda4vS49/CrFBsua
e8oNmrdR8aD3aDiUH2ngXfK2mH6mSSkeKYh+EYvvIKvcv/1lnUpyKVLKvg5KJtovjBws31ZPurBa
hbNcwAftUPb//as2V1hsri1wVlX8jAQRL3mhLQ8xCh5ORAFhqKmLIZTdBcG6CHSi7PyrjuR1471C
pe4LntIOJ+BEt50CqL2UK5hHWrRJH8oubx2iWp2EN74z2Kk3LOLVRu3QStEODJLLxl/e3HEyoWfR
jkW4ckBhdAZTJNDwlXLOkXhCYJmmjQBo7amaXzQXwBD/2R47qWk9gHVA7d7gL6gqeSR6XpD0w8Su
nrUWAvreRiuymLuIZei3PIT10XjiJ3nvLWOlpXrzMoJI/xYSnUbtWHrjEuNCV+9SngV8xc+08wya
PV1wHXRXZIVgMXqX8PnHyB9QmsS7If9S4YN5wDl7OTsQsmBpjTofOF3C53shlFvqn5VQ7KFE8e6h
1uhK1XaYBnHwMJi/A3kUb0IIVp/Y23gwOYrjwk0tBUE18ms9ZoYHOwDlG4cIRcjYpDiQgY9wNmph
CzVVc26HLdKx5NjQZoHvYJL8dad2NI2hy2kS6POGqaiWYBWa6dhmazsB+TPbMgMk5xn/MDXQq+nl
B0Ngvx9D1VHDcl96ONExdrIsHQL6Re9GVz7kQv7fU+yPzGUul2lO8i2BTVkzA08JQAQdW/12Lx4O
ytgNUVjyRnddbACwaRohr1G7A5s9ti0ym/V0Uo9A5gnG7bmLHpCNd/+4NMjhT/YLzY4zCtdL1vgt
XBriu2vq6UUShF0RARccBww3Wi6YC9HJv5zHq3wa2JXeB5ecyc0fKsXJvn4h4ikxQamZK+ppB9Yy
eg7ii1mKr5Ioom8fUFoexLGKW+fcIvaoA3p3t89YlkPhcPVk6APrZNVjinV2WujC8MNpXRxXKUks
jwqi7VCDaUk/9xCLAFpok3LcRjyBzC7PW2u9vjmHKZQk5JIM0aUaocpOPbkPyrIQJpVlsvDOIzdt
7N/fqSEV8XGfCAqOHFHT7zQFBCHh9IJg7n1LpVEIifJ2V3eOMOUU6+Ng6pzILKWQx2Ki08Mxn/je
doF9r9AlMMqtl0R0Oe+ylMUR6voCT9FxLU58WqbpjGgFVgJ5CjYxhVxJIZJXWjAk2ixrlEe691lv
Mj7qFTdvhdhcmyKE+/sqzqwLfufdF0UEeOZC3AwDpJCk46p7Ajool1wF3Xy1YFYnlMX35fHZp2w4
sWzo8aRGiOZbFtZ5b7mE74PneBDmR1DHmWk0cXdG82MkSc9aGF/xFjTZRCUDoex2OB3016oO2rDw
1UECIK19+OiZj/TmNorzqW9evlgsJAXQZWgl2PG8Vr68hMYfAXJdbbjZRHNw7gJ4zqzoUnFmgTFK
6+RPv+gD9KIwme9hf0XsiBCT6sGRZ+ALhBKxjLPmnjjzyM25kby85JMJynwdCBgdu/qZEnncTcpu
80BkyytJ3zSc2Z0goAzRvOr3m57Y9/Bcv/gcufMbSq86J80IY7qe3ghkhqwMUH2qEWm2ZtI74Rhf
mndfSORy+hllC1z05OylOHkIlXzHzuFYtKr57fVRNUR2o912xbqFciFacx1jYXWTfIHNb2SGmRpf
L4Yfdr0pLGEy6axDUYx2UbTaN8OaCvs+4hRdkkLPepsNr49OmdwAIBBY8lwQX6OWPsEHMjPRg5bB
Ez/LZgqPBDMYUTYnN9hPDrRfVhUG04WigL08sKCwFfVbWJhQQlwcEa/oQaPWtcMJSclGMZVFGXOq
RZAnp1ymDQLEi0Suneind+D63ss/08Uvr3LZvyWvhl1Ny7v0pDJhBY9vjlh31hoNzPIUhImehPeE
iQiob2IqGjQXKYeXeYvuzTEBYJMlb4uUNyFbUcOEjEcJLnbmJMffo6AKhYn3FhAlXgUWzkN0kxZC
0A4/z2xU/btT6ECR4Gv4eNQXsn5aoc8QdX0bphUGu5eyZ2nq/tA7EZuFktSoZb1+hZwzc/ArSb/W
t8SmA2vCMoQ8urKqYE+zq2bdownzhI5j3bg9dqzWihrVxn0MQC2DqJe4Xef6wrqS67bVAItedY86
45IyJ5gIOn4OXw6tqmtZONCMbmrfdZinSsrNqSsGWI3kmP13isGDabJ1wgYvkdvCSKKkI0zxmLa3
C3OIJuD/EmRkOeYr8M/ET90Hi8opLbcgcXrr1TVn382NxyohXrRgqjsogCFST/fFKZBdyLpuoiu9
JskiMA6nY8S81mGG7qhJlQWRVdWA3iKjk+oc4UW/EEUi0ZWRUXWmrmmGmbYRf1zqjDpoBir/hvGs
teA7KvmnCtuZgsShKoE3skP3+YmlKUeZ8npOFjlmG8tmnzCkI+j5S9Q8r5Fxv4fiern6H7rKYrFh
lcB1TG2KSu4dZki6zubPjIWitUvvB6GjX/OKcyOC0tfD6dSqTw4u0vl4A1agE1tOQjRpLXPGtQaE
yA8sZc5GmZbgQbc8Po/Ge5XmnfU+pyYH292Wd+4fn99RbcqDpOc3tLbDMCHfHdgn9SMQngsI7kK2
YLRXreIeVBNEWtXRxiHpkZKIAkrcu1lTRhJ7DX71v0SB0uxeP7C1ai7Dj5KJQoiCZS+fV52WYEJt
PFlo/AM9Ztva/yjOY6je/PQ7+mICLLIYvOD2Yem33qcgBLmSkkXyUH9PmSkbsIQYUkIf3mDXGAIz
DjzQGFYENVGOHUhGRBCRw9WNgTx3HIIfLscLGrsOh7qgGlp24lnnRFJxQQswrCI6WUQXcZhT5Uu5
3vhFgFivzFvTJ3mT5Sya28pErZXZpGL0Vl5wMbZRfryRMEHN9/7nRgGj23vymqd7Sco5oIdwC7LG
W/v5b5LSr6N1pFCMKy+4EmR5qiIfdunlkTNDiqoyyYMImcUZw7Lv7XbNxfc6JHO5srhY8DpSH2Ig
yHc9d7vqOCVHqo/Ru/UaONkpbO0GZTlWrpg1VEsaqaKbjvFpI8VdIrXkU3A/bWqHaGvxxFnhlXFO
LVpdhOBPIhXWCexEHhHrbYGtsELwDgGBgLGfeuTdpbOhMBK/5rp/TuaOtf6GcrWnEJk1ji0g9Aey
+Gu5aVlJwN+p9nENF+rRuqkh9bEhuChyzkL8D3ky8MwBmmsYYHodeP6HOH9ys+vvpkbgW5jcv2p6
oTaL/zp7wdHSWQiwtKQ+eL4benYm+v3bzOu4l3KXJDNuCv9OxIdwCvADhyfwGYKjCfE486uvwWOT
65xP9BJR08scK2yUnwtznxHsNsGypELuAjUffzESeo66eU4lccyP8zaKtF71rNMZL+g7Jer0hyVE
+cIQYu2y08lk/UbOpaQeb7Wp+nIycBi9PA7hwyA6FXxLtDMatW82e7oJeSJzqXOYz0ykp+l7GyTv
X9Hbp1mFXR8+u3ttWEFHzX/1T1tXaOpwF5bSZq9oTJENYye69JtDy3I0Mmhhtjchc2/4P3Fohuat
LJombFiUhsY14mQXy8DmGilvkSlgv6kihF3ah2+qGaPL9gfxZbRbx4eoPGjTmkIevgUai7HNxgcn
7BL3wZsTreAOg2PM/bAegqHdo+KqEPDRg6oD7Yl+jPqagdxL+kXuSAXg7cSHgrE+nz/2tRKFD/aJ
nt3j0ohxi9zUGG802MLHqdvcwG1VrL9DmRmDQgoixGUE92rBf7qlcjcJ85BL33qYqIKzUcuj/xYf
8rNJVioSg0mw91nf/hwwr+0YPSfjrR6gzux1ZEseZGxdMQG2pPXzlVXJLWbwOWihRGLedjDScbmk
xFc3XjAsmz8sHqvwePZj9NVEd24kTujkTHyPvS3xY7k8YoW9PTH5stqcLDH5Sd0xCC9/H2BVjlfC
lSopBKvkE+9Vum1/1bcz87cp+3uj9LwmWiHKkCv0SmO7mRoOoxoMN1p/bBSRiCVR5PRkJB+unyht
TLke6LWNpqfxgtHwwS4qWMsP7YXN1bx3jjDjiWuKbYfnubFEFSwnf+5XE6FWY0JqH7Y9qM2gxNc7
GzaTBXa7aKakFedkEQ+/BvsgLjnPPsjIZsXj4pjjYhQZb8H2pMj29fTYCzeXudSBUA/XT9u79rMC
aNRu5V6vPP5kWPG/chGZDM4ShGWQCii6t8HfYi+liMc5ozOJqLRtfpBnnWwUPOkQrjNTFPeibhYw
7k/Qv+MZprQeStMXegk+AcUwVaACpHppfRlWv4ZR7rvGG7DFc4qTdf1HoZsmOM0ZXyjfj7YexTB/
zBDpDxCHJnHmvVt0YoAD0K5r1I7F8uDhVUDxUD+2coUAY+26QktVoOnLsxgVqFXAOWZAayLOI5d1
BISp9PjdDAMFJ48/2SVMLrpw9PVHUS1LIGRU3TvGN9eHhmElG5I3qzPHzbNtQdsQavtiI9ooLD4A
+5oEBoYury3kcwCDatu2HugaALibFx7XWxfSeRTb2QkrEbYYmWiVHb7nw09dE5GB1cO6+1enW9+0
HkAr/pX+AdABUl3AA++eiS4SvdsqctFr6ybHDy+k7l1pBMLstx5SYJOo+BTESsbkFOq/IgxF2EaH
y+FBjuVzjn0OYZil4qg0wrnR2Tv2owHzs+pZCYQaaMay2ajh57+emSSwTCQtt1GbVtedOyk01e3i
p5303Y7Suy9HV0Ivnpc3iLDp06MeCdW8EwcjQsGToXgge2u2oo70VOkeghz1siVe+l/QX1KM1SAk
K9Kxh5A8dEIS9vTnrdAc5KDI5WwNxkxPIy5wV1ubVaiT619JggF4ixj51yU30Dg5hTV8pfshuNwa
JwJdpXOHFtCwXSFhko5MNuawPfbcebQAieZOSEZqVystBto9W27UxO8jP+KGw3cNyc5AMR9gzc2Y
j7VLs9e/h8GEqjmnHl4u491W+tDqcTSVCagOR5jk3CZ4NqwFlsQ/TJPtFQdH7EgcWmArJtJCL0hN
k/cGO+4HExn90bIO/nah3o2j0WR1MVFVUMOOxQjUO2I1m6wrLRqqd0iI34f5VBIDbkZF23f3t13q
m7XWJ7LSRg+6eVE6miCX1rm0yhOUjUZ5yw5xe+R57hKHloTikdbB0iAb+13Mmex6W6azbW7uMYpG
Oni5MG/7S4SOOjT4NZrrGJZk7TPNz2htSQxZ/gemAeeDI9vFrQNs8XY90zTpeRN2kOKK4sxV6WCf
v5yHhr+clhQdJV2mVr18//15CBzwy/knKcGrHKLgRUp4tApMJOCJhbj5ku2ncESIlrpQKfpoumrM
k+wzKj7gjwkD03gfpgpsEMzRcBH0WOCxnRGoE64KwiN1MpMMLWnjcm5KNfb27I2e6we60ASYiHN2
3/MYb8Kq+erpodq+iNGw1MuPZEs890X4h2vHFU7wmoUTRsGIjzQPHMmLwNTyIfG7SAsJQpF66gYU
tKHXGpYsWuHOg1r8Xm8Dnneo3Pxya7hFCi8ZFO6qI+B3oj2xtVgzfaFPki0hau7F50B62xZipkGk
6AfIVQFZCkB93Tdgx/6AwdSxoTr60jUS4smam0QEKXd8nSuatrZ5aUGcCg3huBY1ta2+xGkNMB8+
sGmwPcwTmwebqOyw28Hrqv7ORdyJt94fZzbIfQdGZ425KcNlr9PvSoLJAIRpfgCYmep0ZabFKvd+
/VEvCV2cBcBH34+PXHtyl/Qt6igyDFUrxaDwy01bQqaLCTvM9q1YaZZ8hlVhcbAHd54ukvRbvfhT
zqBiy1T0QJX57LBj0sv7jCVfB12bs0QoN4fjZKtehy8D2NwQnXsdDWfBMGfbblXF9QOkkT77B0hC
awFNGXU+2xzfHNvBnAjhZsCCqMVWChLecbb5bjfiY4ImUPCn/auCoc0zy7FIHfxmlrphehOV5vrL
glZKN6GugYTbg8nP0Un9nuwQIW9ZWOzw+7jwan/TYz72AKjSxBlq3+YUPliLjbDpwtvngAQuTMVs
4qH8PA6awtNCPhWzBtTpsLu9ugsM3091NnlSFwH1asa1Zy584gIdzxiFl8qLIdLsNZUmYr9wH815
tOkhDcS+14JXSyjQgnCr1m8F5janmmIrkbAlEp7IfdKuqqhSYAkhc9bPKHnbX1sAgsFF/a+A4eC4
7i7qti7bAwR6l89dx1xUEY55CDUQJe4d87ldjF8lacCER6PHQojB9OLFDTI1kFbQmY0EqJVWpz9b
zq379jRNKPHPc4GqFs0Htj1G4v4v8gFnPZVLz0Br6i4RGQU8gT1fJlaQ99wdYs8KTX8wfaj1mJg/
AaCMDr1UHDYju1kLtapplQ/sfz492DqsaNXrozss5YQGeNh1PCIRHHLf3UYcChqwmcKgp4iOgl7P
inwRHu/Fh+yZ2iwlkaxLfDPmO1PZo3Ae38gng7xmevSmoKV/ISDa9vZ5laPlUwHQs7sn6VoYS/uh
+Zv7ksiKXe3XGx8lo1o8HIIl9Z8T4QKxeZFfs/vj3P3n5iV/lqpRXeDy1M/DeBUCECQEdicg1MSI
2Zn3D8PuXBgo2bUFxAslMqhas8W5KErm21pyvftE1HAeAVtKSSxJIuiFfPoAZ1T8dl5C9SZG8p4b
u1YbqueNCDjdr/6TbQldkDtv24Pbt4lCj1Z9q/avKG+yWl1M2qsnddoztu0oLSnX/OcgdC55wq5y
Vocchvd3NMMTgqUGytzqk3n8kIAkLgk3/M0Kz01o73fdUmpeR5RmSKS1SnQakk8zKAHxi70/cc8h
IugPEJTpzAUxorwFNtDl8+mxBdFyolIEpMCDNwiB0VmdxcJKu6A3KC6YHZB4ZaaAoPlpojHtGRDC
Hmks5ASxW95sUbs6nxQVgGASaXJDRzqbkKtvD8p0DNmXMOlB/97NQ1GzACksG8RM7ePw7vPg/b6s
6HVz4Yo9/devt57+3GabXrnU2EIhuNLrpvf4tXZocJyYW+2u8bWwPgHgY3FFh/TEErVI0TYmHSRX
D48dobLm60Xx0WQFBv2SlosKnT6XUdnoqjuRKFfxSSmARBRmZOihjTh5c+1gGkTAF18pSX+QgqEK
QvmnxvTKy283rdop6jdjl+SPeYuE3+vtPADZNFlBy6+hXHfgrF5CCox5fcIwbzy7jChtXM1CLbNo
IoBx3xGZtnFfla74qgruurLOuxc6Ej3dC2BqO7vsJKzL4sk62VWFHGBEb8QNpTtn2XsnHrPvZFkS
q+P1aAKzo9dDjArwBf3+lyiQEzDlPaYrNQ69oAtpilGDmq6R0MKIFZyxmR6schKt9yucmbS1z3ks
u26vwqyYleb5JeRQdalT50YbtRx7IpgDDUIW97WRr+98ZOnwQE/AGGmlBbyDtLR5ByVjG6QH6yk3
LC9C1EPN7Cma3kB+dlRRiBnqwyzjG8cSm04AFST3Ekzm0Ptff+w3ow6jQ8NLcOrrGmYM/aparA8k
uRaAUewubscUEmbFsiXpKFOX+szpMm4DjuCpgWcfkFJggoRdeNC3kqhaHcqypGQ17AD6ewogJgIK
nJeQiatdeHiinmS7wSzYAJPQyaMCThEv56RqO2PjW4sXGjco+PxxLjCP4Id+JrPdzGiXnxuegO3k
GsAU8FAsibYovq5n0hy7e1X5K+gAp6LLGPwbO59twywUqDUVYk0nkfOHj3p2m+z2TBIkttk8YdiE
TBA6HCWQeuvNcxJARvCS/78zfB1OF3S7Zwi6jZWl3vsS1TeDuNfuoBHEDeBHMJWzI52Wn4QAH8YT
34M5LagTGzsfkq2L16V5iNHJ2SYrlt15aSNLb+D88sce8/ea3Q357UibIXZ6teqxub52tD4rrTIX
DKZkRImVAwydPaXcNjJEDLzuzG/CMc4SvY/IoDmqrQ20m1ErrDOdMsoc3s28HYmexJ+7sinoXa9x
4j+tlQfkwZqzSd46X4sUoOa/OZNy4u7IaVPfGLT09ZxyjLTGP4rQR+gZbXnXuHHnvTG7ZyURJDs+
CtNciOF4irZqEtp7RLf3Qwgj3SzXQRdpGEVS4TfuREabSCbkgyBjWFHpQLQHvhM6URIK2p9/lLG9
9Y3wHB4KG/cHbS2dp0WdKkJMdzgoCEenYHQtiZzG101eB128+Z/cRyHKShQvhZlcwrBS63JiHr1u
BZ3Q0d8uPqNJNAOgdA9QvFWQqOfoDt7GYNa1WAMaOURTbBCDaTaigtSbaHwd2fhOkfbAU/cMWQX+
lUnoaFbh0e8fOo+k1ngZLXjvyPmFIeBMd9+gQSql2VZWJ4yYjWLjlekQnGN+PhbMZrZZSWBKatqT
6PwHjZJ5vtcIko5FWPB0nAj8kVNvAkKLc0NJxdyEdDuQjMRfNwx742aXzDQtDt9Qmc4SieBhVEYm
DEFWHcxKWPYzkMahMD1TsSSGJq7W6ezKKDcNyD3KbeGI3cD4RQ4btVIQ/ch8duPX2HitlhNf1mdA
GhgjXB7X3xLNylo1+M8xOMAwM3ZE545d9Jioi4l2N0zNU5u3bRbzItps4ggMuuVmKJiKEwjlcNcd
/uuAdAfzFuKTwuDVWgbZV2odvPcxrnVI+KQ3gaVneHLEdOBsMca7s5VvKUsRJIbBGq0BFYS5kRMv
68V5JTbSHL2jIPy5YpGphT5BvnnY5gpI6XjPetk+wZWE+xvcAEK09HmOTmNwmFZP0ha9WhjvOvvp
CLB4Hrpd7NX9sw3RFtOND3ucm0eR4ZpcRy7obgBXvzbpFnRLrvp1QTZLJTSujnCvUAwIpDVqnoc2
IOsj7yb6m21fDuiJiUsRLXgkNG2lZNg+jrZlG0AVkImoPhYge1Fs3VGHuYR8faySw037BgtKpj+H
vNxcJjG3SXwxQowz1Q7hnR+OJ3/E9vMn1M9bhrOdSWh/TItEUr4rDz4tI4JL21Ne9RxL2B1xwbF8
6402yyn2VpwG6C3SdEGXb7H+GIckJ9+vdosYwuwg0+DEVjp4YcRh1rn9vfnUMKRus5VYy7QxqhoP
ASI8YBzac1XoJXSrHb9PlYDXCOuVVhUazMM+PS1XyalJyNW4bbefeEiUGt8LddghQEuub/XfFRr/
ZBm1X0vzrZKQ2wdCNcHpC5JLUpOgePKgVOXk/bQcdmCcrzQL4yFMvRNuegnLnp8Wsgl9dInQisa+
kkkrAiiF/CxFSlKA41pXWxb7kgFVkuPAtoy2oykzyoyiAz/S1P1CMJXuZKGTtzVhvs+g08YyWsGf
iYPrhemKBaae6Drfaj54iNimXGBUohz6ePFeylUfDlRN9Cv6sdj0EtYNy6JkWQslHbpOoU4uJYGG
d019Uj7jqtRW4Mb5AGpNkpGe7nGTpJv1iJr5bcgdQi7Yk9VNmDIZiALaN4PRqCP+/5n8uIDUtw5i
VN4tSHa/6zBAmcgQek5UNWZoV8L84rJQvGiIHVvcYGF6rkyJiQJQ2pWaXI5g+enXfrtXc56NMIuo
qg/5qDA5TGSFmRmOTOA2ePu3ylucAAcyjoMWUlpSUm8LRbtgwVy/ci26fGTVQkFgs5Vm0K8WkRnh
Z81RUAGBAnzMVRGuxnhfZjY+46IAJ/rLJ4PWmq0hIviYJoWedmxaOw+tmeCmVJ7HiIBhnn9NyQvV
m5AXDFW7REDIXIHBG36YU94G8BoAnTA1CRpk6iZriDpbGzOHHMn9kCFOrM5574lrIgijWWVInE97
pg7xqChF95gXK7/gxPAi4G54sv9Kl+bh15xb6sWbXPEKbOcvZHRWDwMqQIPgg1uiEEycWXEt8JUE
aMmEB/k/+LLJQHfpizBPBSCNpvuBOFUFvOugM8O6HeAq68eUnmZ1Ql+KECHqr6XcRgvEOO5YwC48
AcILC4GPbZxc3pNKjQRZXmZ3mivVXPwajn7AgZCK+pDSrsDTjzFHQIBtemnF8fej7Q5j+IAQYVki
WF+6WsZA+Pif7VV7HVqMg4zTigcGrz8wTGF2EkdJnihaE77JMfwXyTpDi4+RcuM5MHrMsepQfw6r
UrR6q+NOV5KVyy/KKY3VLRRpHQI1BWOkZ3HUrlpZowg51nX5uvcW9NkB0Mqe8jhItMVbY98XOTI6
m6P+lHH9xXdnc9/0aZl31GfkgjndNYTllq3NKskn6YaFQ09uW0IH2kXBdWHQ/FY1FewPikIXhcq2
E5bU4amXX9PFBmM/0FhYhg5oNZnot4QG/dNc2jOJYhoDvKyF6mLkkDD7ywMn3ceFVYqqO4ms7c9R
3Vs3XzKOIqq/9nQG8NKQIT0aTrPSIF+JxwgP3gDlARkk08wlAnNqiWd4Pn+1/wA1yBcMCfvNsfDN
Nryfcq7qiEpzISOD4zUqyTLqfEaU+7wS5tsodP4BUpzNezITN4p015AOhQ1R8QgmYnOLluds+KG8
VkBTpY3vLe1UGeQnoK30ghTgMXt86JvprNjj5f0YrjyaZ+JJq+WpSUp4cvT3/0gkgqjtA3EERwRx
OmXJeOKNcq2THAtZsCivbSYd5x4QDh6swUCnV3QuPCltWbFICAEf+WVbjp0e9uJG50wMss8Xjhla
50xFgtVg912vLppKZ9Q0kwKGpgZMuTs3shQzs8kdAQkfHGOcnirAmv7pYnHn+/+pIM9iZXwn524Q
e2WA82KkxFo/lHhu35mHKFGVRel8S92AaJcuif+W53pQapmyKrBZbzL9AAoWriY4fHjG8HNcfNJg
NTgMdeU+JPqL00ZQExwLY9EbkdmXpDbt9NFBPwiAOxYQuC0ReNBNc9xHX92vrJLm+0Y4EKq4FQor
MQYUfqKAmrJ/ih8xCaC6tsdLZEQ51msG00tFMOk278nw/lfyvlvHRFJdrlWyPPY+sYqcalprkWrL
h8iBCnQlgo8UvLjjfb88b62ZA+vyKF3qkWaby7EjtKd9zCQl3WfVBSuveRo4V98yMUPcE1nJdiWC
LSM71yvZPWdq8BKy33R2YvxJl8ADE6wF1fU8sK2MfUNyF00ussfzm1/4HUbZeoVKCGZwp/8B8IAb
9vIrQPsCeP5AhSbn6wEjnbb6jug6pBsxPLCA62yVzb+uFaknsJb1z2t3xsM9TQ+urh1Mm2j7F8M9
vfZ5iSkN1qx3DMsANZCMFlcfjWN8u7zlg8nsPhi/PA9RtqZfU/lpfeHheGxi1HkBDUsaaq1l+N6o
Y3U7GTcT8/8zzuv62hwfkqWjaep90z/aDJqw3h3IyzFbazv2HHgT2vRNc7Ev8as6t60xwPLS8r7t
M0l5rjK/1UbHO09pjBsmOfTcO35+UCz4c9bijs0XnTM6ygN3/LvMuRLBIyHT59soX63ei+wHa8el
ZOh7+5uzWzj90t9jiKdEi5H/xHODJaxf1YoYaU9E3boeFKG2tSaJtl1ZGVYz+TK3+aG6yUEWMuNI
90ppKFuMGvXfrS2gqN75Cdrw4nwQQJRJXuJJ702562DZjSf+fyf/5FnBpdAqFeBGpHQDKf45pdUn
2HB4UHwEus6hmRhsu0PS4cQ+gAmJWKWWNHMX1cxZaKfl0gBajg8OFuiPMOh6enlPtBZnlD0gA1EY
WKHyUeBPB5RbwxUeeE+Px3IQxk7dYPrjSG+acUN9KX2KdMXkcF+PeWeun/189SvJFBIY0yA8ZOJP
Qot7Cr9FPvITZn4muncNjDEk/CJC7jissBblZ4WIR26DhVfeStoT35JpCN16/xx3UT6nYiMiKu1u
YMu8MJ+QEAkMMWGpQhYIQwoCJYWxGYSvj5iY2e2loZhO4chpDdIMQCMP6TPjRuUYGBVP199DM0cO
eNV7JWgGZ/Oz7Vj2AyotLLpdGUzdmV9LNdemP6XnHpBTLjsUXiIvDvRdt45jM6/l2INNOwUP44BW
efxchwZdaLiPmbrcUbfAixbg6a4rSHGpTUQK+EAdelXZgc1jc0nTak6OhBuhBCxXix5AvXhFzFh4
SocNmzrIOg0prQ3YSfLmavk7kPuV3q7AB+LOOb3uw9PE55vakPJ4oQQMRkpBNJXUtz4USEoYqs5r
tWOHQtPQHQCNO2/i1xpIluHASLTVy1KCEaylodlGPP1QeCeeey7oqkRwhLMlocrfhPqAnVPghUnQ
aO5nVQawoywnLxozzr5sXBiStnAx1Oqg83xPRudW4RBAuLOzlNNq7ceajuGyhL133PNFbYdvuI7G
dguMzm+tB2h8Bu9+pNKxR0ptcdIQ6RW3m3cKv4Jy+Z99WBAB887QWJRyVSlxOWH3HV04sEuNqZKQ
m6yB9TlCLWTl7TXtBp/DfEEAUBzHoI680MBp41thHVWZBuk1gqY5NXXONbKC7MVDJXkKhocKkHYH
kOrD0y0C55FMp0rWp3cVwFOQ3iQ5VMU7lWDXul7KnRaGG5Y4qAmElxG/JOOmPV5m6W6CzL+KRrdG
9Gtssj7jA5/1+YPDKyMaLnqNPhjyvyL8Lj2am1HGXDhbJdPSNlPngAjSZXQ627lxXr+nZBtu336v
cjoe4iKmmUyjE/NPhV3cBDJpU7jWe4KLflBA1akdOb8ZnUyAMvM9Kg6onjgq8Cz36eeCNh4WGLEN
K0C+E/kVfTqIZ9zeTcxeYEYnFeCMwjr0yaYPcJYbyHZkVAIad/JWYmDG1/4O42TLTTCmgiAvdXl8
qPiVRyEYKIJY8GD+IHCGEj5jn4jbQO6bCcNOP5WdfOaq9rFtfD2gldUV32dBLfH7Fj4lUHSe/37n
4z79DpMJoh3TTZomtBc389c+XQ6CX17yQbqeh2EZThknn7tt7181fCSixd5JEewo9LrjEb7TZmmp
Uxj8yZkXvxmZxzoAq060+ZL4gXbzbnf7hcMGaZ1P2cbtEFFBaP64UasWEDvu9IsHUC/g1nd4yoPK
XOyMSh9LooNE+5rMzatWOljr2FtvZZROuEWe/GADOfVLd7qT1ZISsVyORWgTjlwh1jgP5D0TIEiO
V8iPCn6iSj5ChFnJK5BY93qmijTDbaZE+o+C1VVAmPMqycqrBSwqt/l0BpIHRE0ftLCVm9UGmHf8
kVhdCF9aQXNTVYYiqrseWzpyXUYJxfU+RtaGqYVNL00ZUCts7db3LawjgUDQEn+UmdXDKMAmLOm2
KkJvmFb5dj0HYPfXhQbMKMkr7VDq34V3LGnMKLpukQCZwyykm59yTpXnQhK4gmJm5DUcP68GkAyW
kkXquPc3trx7D4KCltxUA05zlxSlyVLAaJ6W7J/5XEVOAP4B5IfARlK1JRQeIn+GUE1hS1QWkHZ5
QEgwsgXMj3QT+4W0bVPXzGdUOtH84ltHZRA9iP35pW7iA9WJ2lrfqnjeImqdO5qNF0Z1xdZozLjV
JBQ8+uEH5tGhlFgXRLONrpIRs5uqXJILdnP3ewb6x3tYSnmeMKJA9wAHFvDrB8Dj9mW+yYzqT1lb
7hMukt5zJqwUWeIYw6Wxsadg3lnmgRgvfNY6Di2ugllN5vAZKWwiveD1jJxPSdH5OKfIkOhadMUr
b/MVcmFc/t2fWki37tY528u6MJUlrhCxunlTwaG9yVlqn5F9pW5hXOd9sA8ovRKCs7r7NllsJ3K0
KJ0gxwTmqTpGj11KqvZ5hcFeITuSGn5P9uk1uFBy2w+RqmngBBDg9RDGV/RULT/ngK1ZqYWdKaDm
xy6tzEKKaBhc45tPomXyglkcoBgxrQyv+vZSNM5ODvjZQfvg6Gs9J7xMXlN0ikoOq6PIewpxAG//
KDQSk3x9FQi0szN1sfFlFhHB38vu2AsUQF0wGcVn1uD5Z8j7ypK4t/hx+oIDvuslg6huRAydpvFj
L2yh1PnRktM9FP0JOTgg5sHVTValg+CSapnED+UmJTqtcoU8I8Pu8kL943KnCAgAi0/O/cxSAywQ
iECU3JX294S0OXEK1i709idH8KydV4SnZmqbBSPwP/lHaWn6IrehgyZsVztPKvR2RxF6i/tfGUTn
ZGG9Wg3nrTnE2aEpwFJb4N2xNDbU2r+bs2aflgV0BdqUyS4MrTVdxxLFhX2jA1f3Br5WLJijSmC3
H4YoKMZG7f9sgTTQqY8/h6E5gZCJp/EKS+YVTFsFAoY57Nw0lMLKn2cu1R6+JLO+ydzjhaR1KF7q
GclAvP1HFFmYo3LIIBLHe4AaXhxCt4v/94ZVyY/R2o0GcyDf8kNZ04L4IO4BimP4hLiFMPTo9lNF
zxgGHpcCn0cHVxEVJRD767f68VHb3jyWdBq0ajri3qNAUu5kvw6cufr4ewzFqCM3JSVEI8+DS2KC
9k07jJaJkFXv+1/SP+K4l9tJFsxsHYhB0akkGGoYYwb1cs3F+XnhdsOiEZZQRJiK/krkog224FwY
U75CiWRXhUQBABIwKndiiFY2YEwRC0CN+AnAcUmINDUSpLSE3+2ZGgYAle3B4Ghoj5pV3l0/AnAL
l4bmhfISZ5uBWe5dyqu0EyR24DR3xJKVY6N8lrbAQb7dvbhVGf8Awgg1GSYFTUZSo6NmsqQQMJKE
HdnRx544dfNNcIe96tHYnC8ilVXrYOvmYq+rLKayh+4YnV5HF6ufSzYqWVIImWfGOn3Kd4RebBUS
oRsD8PoJ3UB+MuaaKb3YieHEIPjiZF1P6hdH7XEPRAGk0wwv+9ND6yec5aswezw7FlZ9642oDV0v
8YyQUJhSW5/Bk+Xqsp2KMQDMAu3Xhh8cQP+sEcIwgvq/0GGbMQ79qcfsokSIRjAsECBJ/sZzuUmx
oFnxXSa3uslNEAlRcLlrMkSY0MPNnkg61+g6TYowJmsRhkUYfy3ljeOqycQZG3ip0BPOhF3sHkbt
bnYgeSwN+xZokHFzLDGoIlAK/ABTSzd3Sm8cFTvd/2af4CJYLA4xpewzw+FPx1ELWWHGAWX7W7cr
/htTqAt2+TCdcT/WUuDZKWc7Yp2VCt2/x/UPtVj8+X1F4OvAsm1zd+NpvhOP6BA//O+j5nyPrc9e
T46TpyF4qfvVG1kd6rIH6J5SrrS81RaUGJ9jkIb3lN2viS0VfZ1rqveTMfmNuXbSU81BEFEznUpK
BLjeazNV/lr0F9IJrinakE0/iLVC+oM157bbE+14IZec1uWjNykXWMrWoOoiMpF8UZ43hWO8aBbH
T46zoyA1lJBp5bowILX4LaC5Ck+Ghok/vt2SycLp+M5Ugw4avLcXXQIrqsGB1EsGwJ/anAmfUfq/
JhfJDjOYdDzwIJBjhvjg706ZGnGY+c3KdrC9jtwt2Wt6Ac17MBHzD1I1TmlwCwO2d+S897bAhLFx
y9zd2V4IVL4NP/pfqvS+uDXQRaERqUcnOq3LzubAMi5Jp0Sgjuf5p6DGP0N+b5lytZTb0STBQz2Y
enNuqR5HsCZiorzwtfDzClHm22GbuIFTuqISRRnApJMt6skNzZbgGE1Qt0NJCWDdwYSrQqqXTanw
g1T9AtSkJNFYpnp6kO98soSSMgEyMvBtLgYzfGq0IP1wpiAskjZRxvXSa88g8dK6edXLhSE4BJGZ
bvijTL8GoS07YjKVVmyZO05o3tdEiNKQm6inbGyMwb/u6QCQMW2ytXjstHymqEO0zENpDN4uqOMT
Sks3QyXNw52Ph378lVkKkWUHLkpC9c/aQnCanlF2uzwNjw0XJD6meyHQAs6YqFGLw8nAHyQB9feM
CrBak1z2qJS/l9nSus3D/eXiUinJKaXAdIza6xaCsB3tSIyYX1jqknhYfL3F7vx7K4/+26OToy97
Nwt3jSDbbLM+PDhl0w2eXnkYqDPtt3S6wl6MZKqZ+TA8gUejHAvDMKCb2wR6auBlrmnPDoT/wQNO
OLLhLJQHgQH3jca9P06o0o3dyvrIQ/hAyxBmz4GgcQLTz0NcqNlSH4g5iiYUcPx5LGnZshUtlcub
NPwce71dHqEivSQH82qLNHSnndvf2ijTXMoWfYU+KvN9PGepdvg2iDT25pRixMuCJCXRGCn0dQYO
Aa1+1tUlwLG/TxV6xp+cmvSbRuW6JxOjHPGZ6K2vNQBCPx4/C4PLzA9lwFaC5H3IUc3DuUV4GTDy
D1LidoVhPrYAXFFxMBdw/Kbj7MR9UJ4xHqPSJ9mEsvnnW6oqylN21pYlUXdvNDMiZRbjnqLFbVQ4
/DRC4fkfyRaU7LlLfnss6cY/JZl7bCeQYFfvcW3E1nOGZ7CBPamALsu7CwdmuVuwrhTA1iYvWlhC
LnQsNHgA7aXCGJyJFcB/TyMZzJZfC6bF1oKbLO5h2LNM6XKuIqq+B5LVlRorPxOYzcF4NMK0TE8x
++OjSNiWhZY9ZNWrfV6IfnpQ2sr5oLwJiLQyYDGugTq6Zq85Cny1ZwldCIBDp5na8R7dMulBM+Me
v+tu8FyOE8vieMdUKNYgsDqmVCFkJIgfDnuKFiXL6dEkqsAzdcLI1cPul7dBbfkcQDWgSI2+XUEw
hV73/P0j6hSu46DX+aMyHJtYw5MToGfH8p99Ni9yymeJVe2HEMihIXsAMz/SCGKac9FH1BXVxGE6
GPw/ashireMx+xDUt2eRdysvGUnmJ+uvlTn10Gkljbh1B0TmgSRUKvJOzEWqOnPk4KUgjnD6xbql
sIwU4FBWVRiNRzb+4tdJ2Owa2svkSlGIKSFStWyhKs3VcnCTYgxRcQsIjiZaDNrL9nmWfFOyDMQ8
DiNQvKj47QyMTRY3J/GPvGBU1H75LuSNK+FiEBkZHyOhku2ANbhS04OHwc5LukKzzUd9kDB+9SR2
jEa8VSoAlvwCTdnx2EKl7ij6U2pas//oaE0GkQU9DMp40lHp6AZ8XzRPIASlNksgb+jdtUe4tiKT
Vn5e2Gsk2z1JfseB2vNim+5VNmpxE8NgOjxBJBQhUiqinaFT40wVy56Hmut9alx5u1qwqyGifuAR
6lQUHYyGLo3EvLglio+GTgpeBYLHuwSYg5gE62x+q+KnlowCikf/trKBiWPc/a0+h9OSsvCmSZZ5
5awkAITNZt++9EsLQvrVtRbny4xnEE88masb1o8DFctk3o5nx6RGt+6m3WEWNY0RHt+ESZ98/2Ib
j2qi0dEO2bEQ6HaK8cTcQhvM8tQUk26xZ9EjENNcR4iwb8GnZ9Uq+nnUwD0ZlcMkgW1AfpvNflvo
LABnVGxSM7M6nuuM7/hPY626dN4s1776O3BiDMx6xNPEtHQXNSoLJKvjzGCYuV0FPZj9tbpi2898
cv0TCsf+yzY+nw2l+XOveHa6JDrBPLXKDH6hsYCPLGgqv6Vs5g8BIb+egRgtjGdOsg3Em7C6k9DI
TNFlPoBo60RyreTpzfZSPC9Jcom6Xqc/IpIdks1RbqzOV9aQE6joEy3rdsgkpnOdUQnAL8hzqpim
OXgxMuOT2aTEVWNJovAHcVQ77h5bwaR5KkWonY5adPzqAA+wr9AKfdhApa4sDBc1D/CeJ639NcxU
LZjjAt8buyKMQDToGo92kadHpQvE7/5AuyvjFe/EKSs83is/eo/sZbzIwxFWzsTQh9TVUm220+Ov
iaaqBQyG/glpupqYNbAfTB3s0befHsk7deubwwvGgTV8I4/k0d1MVFi3EyEf+Ei/zm1JUQFf65i8
8QCph7FtEGytFilKroPJ8/tQxN9ho1XwNp2cW+cUuctXeFkXIbEpkIQ+F1tEWrnh22Y4hABQMZiq
16SqZq6h0dfu8I/rTp6Wd+fCOYWjM6qVGRMezLEnBow7fiMgkvppRihqTiAB3kKkZGmex+S11igf
SI7DtJmixSfP6xsEsafRr8q0FJL6UPHTtJEIZZrNV9n8LQ4Mv6d2RccPfoqMtVfh1WMTfl2YXjwA
5vc+wktUFWsMyQN3A6YwprJWyzG8AWO00LutNAXXcpHXrff7x2KJyZ9oyuCjmiUKzdrqX33YBOer
byaBAZ+3hZo4hgKZsZG6naMJ7P9KE6cBeZkswmI6aG7bQY97wRVraQkVKMGdQ5LwE/Pe5zbbvTXa
UqKITXKqqi6o2iCY/2iCmOyVARCI/EPZDoVRrFHYdhtvYcy7g4IlnjapYFa01b+te2vzeYPcsep6
cgbCjOPHA928fkRhQUaH4mUI2C5dtS+oEakFJPkcG9vWdtPVrXgMNotvAByajy0K0coQbpflcfHQ
fA+tPIicJ8L/WY6j+lsIpNSrb071w4RvLxQxSvSJKTH9OlXJbKhgtpfcuwlYynrL9fs1bl6juqFC
HUbmqyZXadiioKMCppVtWpghzMC/ifAFWYHdyzi1kmgotYmuVRNXcKQcLLHRT2K7Y7FmpOnHDKpS
XW5P0aKpNgpCZYCiTvKLT2WNBH5icMqJGBv2MgUX7kyqGAEsnB8v+QOvMdxGtkBhWMwF0WI56Tym
zIEr+eO1exMVgKVjVKQRTt4pd025rFLWB2EWNGAMSpIdL1GP4GrIQGxCaSWqiBCgJLnVqJUpXlV6
UHfI7BfZzBl7th0wqaYBGeXJdC4pHpSujHKGUAUsGCJd2Iq/kpT5adImQrJy02hCsr7W/u5BSY6m
c6ZYno/8g9kFeN1KCkpmcxU3titY2e3wkW9zwVGzophz2Vm0XKzEowjcSJ4ijYHkOkgzT3xWl1Ki
ydObuTM1SSXO54nKN//vD3we/5QN1Cq1MsfEfDxw9BZXooJr05y7cnHwiX295sFCYPjTYBEGh8xU
GECzVaIT6uOZUJmNIchX3cBtVpDRM31wif4kY61BkW2DDiuGrUClfMaceYtt9NgmK8/vRKIH3RUq
CYxfP5KLMZNzByDD+fNjmXBPeZqxays/cHsxiIAOTXIG5nBsbokFfaXWueysI8TcBHLYW65CsHHt
k+93ZPVGOfLTycqaXCwf/DzTz/28ncIcOLAGMXsiHKKr0rt0cK37HXL0JvxoVcr3d5IT8/XQvbFF
NtyEntSeZRU/by3d5p7QqDpTnzmz6I/CamGMXggNQ+0dyO20YdL96zyv2yZvBZSKETDV1PRDc9uD
UBFZNr0GoSEePNE1wDM7pLShqPRbk10Q0NdDhe51r4mnjnaCM5XXPgWJcKlNm2l/Fg5y93ibG7Wh
ivfHVUYwTTIspvptEMDGr3CIJb8hfPA309D2HqDGYUemiTqKu5XKYZKg1RQoUmMovuevf8gb4J9v
DU9sTEHsbFuswuULmWUBZruJHuiPACVq+zBUyuBPNR2bBdTBFJ0MZX8dWT6JtBNKQvQjeIlAQxWO
KR4PuR7k0DSWvyu+NBaESsiQD++mqr1WO+XgA96zyMYzIuckUr9qwiTnHQf9yfR2HjsVEk0CKarn
/6/1MgOj10epYcKqbDQidzLspYqPmgHTsuR4ntbj00E1fIOmoWHzRMjjz3dBsBwl6hqcpevnSEER
VwTkAmeNFGOJeDxF83hKxVHKZlF/XULjnlT6c+DSGla5/WuRQdd/COLEpE24o1Y3XSHts1DcVRIT
vL+gtxDB9YOZ5xlEpus1dY5+sUrOWocbLfJmFWSTVM6zgH3+VSW02OoKUpH/oNHjRZMilw/+S1kY
/nGdL1RL7AS6c8cbp4J0oMDRJ5aKxWHMnGiwe1Q+mdq29IPcCdK1H51rZa5o9QksDgfJTfdGsMu5
m3M0hSd1jTdOOXayDfp+lxzCeb0kQfmG2+81QY0tJNMr7Izf2z4HlcsvDlXx5xvq7kzABTEZxke8
rRbhUTUjzUk0w+p7P7uuj/rnedufgBiGG2U1IO6qqaqYS72VmONskDrGNtwqCX1iG6H0oC9Q3hky
1S1dndJpcwgqj8Fzv6ST5r3CUXNDBMkfFV44EysGOm/y3AcMfv2XD7IPqlRD1I0MMVQauYFS8dUo
k763mX3sqSevB9qol0oeFh05mhf5kq0G7Cs0BnMtv6Ud0NCOs10QKpZ/1POopJ9axpB0AFv7om1t
kjh7+phmWni7Ad14aapKmlk5qPt+i44B4ekkptSnrdy7L/GY+7YsC5dsusqAV9xU1kk8BcRB7HI/
Gj3JzApbDnXzgAw51Qcf+9RToSZ7IgM65LWOTB7sTqIv/ayeZAsBmjGzKcLX7EjGs4C3X1Icbcgh
5RDUWBfv09RoZ4/uvFyfpgi85cL4aUFdzOlsQ4zxRw5hfYS/ERTUmE6Wn11uyIyH4e2kInFoyGnt
lwMHwpo6I9j7Er3bDHCX4ghsxjM3pn6eqZkDw6gxe7Ac2pYjKbg2a0YwPyJI8RtCWmhvyHZ8eCfV
6S+hRo5xxWSinUPUZeKYMGlN/Tl8BL5f+iSd+iViEhoXZd+4hQi3ocY/n98+tjlbFoirVIYJ8ge/
O6QMVCLWUtuqBf/7CNm1F7bbeF7J9tTT7MqiQlYBai2imyRUQdzYxGQxRu3yVemw1yY4sotd9uSI
popX9u7/Ld8xHGGHtYxchNfi+HzQPwDGmB9I/HWJ061R84NGVAf9p0NKa1fQSo/h5tA+tbI1g+oT
Pm1fcWpFofYvV6QkKAzkcZc+zzwaHjIbn4MNZDkKn679WNC3W0YOUwAxVaH5JxKA6zTdBBpWUY8P
yUBhSMKTf9N8PvUvIoUItdErywgvapQa11bsRWvvlnUo84UNS4Y0hBt7nlUyqXjlvkTsEeaz9GcO
D361th2Eb0pa/3SsGVmOR4L3KEbz+sWn7mvfWZVByuNO6pxpz2RSBDM0WC0SRsrpku5jiV4azKrw
3f2F0Js2tDthxk67sldd3QB3RgAnrT55DpMmuoyknTYWe1ZKL7I3y6MAUiSOal5gDdNxVmkZwaIX
Tp62C9BTHW3UPBBA/Qsm2kMQ12ZHv+1hDkjAk3E8aqe+qMgynE+1PLJCC1a3nqroRJZwjiWNLSES
jbLZcmssdsFxXaVrWyUAKXVLpc4C2h+3x6aTbzDNwDBvjoksA4ORCKte3yGiZXrGCxCYwyT7+5dm
h4QAj9Bx7+bYIPYWE4Jqa5OV24/4+4wvSv3vK8aWg3N6NNYWOWqBG7SjBuPw2u/8j5lqVBCrz7ed
ABd8XisFyWImCL3mdXvqBhe1DagaYMvOL4CxMQ+ghvCzeVXfzulEL5KNjJQWPbARUWAe+vJei1fT
DQ24252q1shFFC7m/OQuZTDCkfSNuf5vv7DS8BCCy/nvyi7vw7PEl6nLBd/zF85lK7ymsUqv31Nk
opzZFEuPrxkK8U6+khwAL5vJadGOBX2KZ+jmzDSxmFisiRxYvQbdxNAQAj/0u14GmV9LcAkTDy4e
b0G9XvWE4dx9CWvnEYKgXjwFS6rYmUQ7eXnnG8GBDJ9a8AYKdo1tGwgHUdzBPORNW72ubiDe0Ypg
SVDYPPh+h/R3JhSkUXQJLkqbJt65vh6S/yI0LRmdizyFfknI/FeULXzeaxhE4VUx7YKY29O1UkgN
HmOsAic2JG7/WjxcCxE8EGBuxmJHVteOhD9pC6+VxEgh2GZBZfjcLzlr8G+XExBiN1t0InXTpkYZ
BH3CwcfpqbamjNEhbrU4A4/uDQlF6sf0LJpvSHcq6z/y4pq7nAqYmg7ao0ghrITFAiRbbdqt7EFN
bytbCLjcIed0kjOHtWq9chDVmlyY/hVKX7c1O+1mT46s7+SxqYIF/yHggVjI/bz5VUTtwBSc4BzA
vTwxEAe+Jq2Fn3Nterc2GcbOvZRh3gCg2UWWemxvt3+CpD1ZQ9520OxrCWe5FqrwIuLpl7Laf70d
YtGbmBUJz/QZyd3YQTwCvssZrf2nK8+icTBW5m6Mg1aCrbd2t3z6CYf5WnD8EgemYlQsofjGro0O
m4vuB3rAPt6rtUbNI75CriccM5aC2sfA0zHWh8opV3UsrX/GTaAHsNgoiLnM2caOmIV8sCayloK8
DjC1RvD/dOhXQnS9inxzPt1/i6d1qdsVBVZBGoJzQHf53we6O8Oum67f4vzdLYkGnNVIKx2IBlVj
G1IBV17HSlh/D1kGBF+wW6U6d7gCXqfnvZWSzQJmYdfffIYEuE5Bz3gHXfCwWJ1Qea8chiWEd2V9
y8TDZYl2qWT808yndxqv7HuyTXT9rqi82Qw4Mhcx3nF81VgvPYz2W10itwgstHmY1hoA7aLWJlr3
FXmwkkPYiG3XrXrzCAWPyPmCxc47PmQaFLpm1k3GAnIw4cSaxpr7vJFsZwBu9zYvfR/e3tmiTwdv
5rpWBtI9hhQ/uasZzGTflfxZ4LyRsYQlvLUXKvQX6gZ7PHomJPy5y1CQDGvDi5aXINwbNljpK44b
EcHjwA6G6zsEY5D+LJIFRYlHcU4IjMviMlw5a1b5GbUuy5GBHkrMUWwgpRciVcIUUHwovk58jxsT
9p+r+Wbdrzm4m1OKMdgk7NhQFuxdfvlJjdMjFmp/F+1+n5o1NBynOVKOKejrFHhgdWjsZN4CD397
iMm5s4aOWRfFF6Ph9dC+R0bTZXWl6FKyL8UQXUCO+irXexjMLPzkh9aep6LDReZqNHIw5FL/RoHE
PhC/+UjACKP/7S8uMaohQe5/mq+J2OoN+MqXzJ0iqg8qmB2aKoQbLJM1otqn960dN6llXd7LD1uW
ZrWnkARQF4CN3/XV/SBRQ1u3qFJS1IeZ8MgJDO7eRGfr5BVi/DjNoyQTtOOZ+DmqKRl61O+l6FqY
j8isEYUxcaayfgT/B9qtCJaNFrUj1EVPBXa1LQ/56SIWHk1PeombejcxYCJFzUXg/zXRji81TPWi
w+H4C/qfogxr7ks395rMgR2jnGqSiiD7T8Ltu1tK6m7BSPJOUV1HflvO0Yy78VG507kB0jBFaJi9
ct6LzopzNEy5ZwWGYagBQvlXjQImbnZYvxzjVR1011euLfMCuURB8CL0dFOvgSp/gVQdI8ylbxLS
QHfMSu60HBcf/AdvJQ7j99B1RmHnQljEXv7DX90mSIjDmRXNz3UOWEGacCPGUXdCNJF01Wx+7XJ/
0CdkCeYfeSez14qB8WuTL/g1CHc752hiEdA13EgwZI8E2DQ3nqRWaPkELq4k13lrmNtpdp5IbPlC
bKgg2t+Out/66nd12ETQvP6va1YMINQQl2QivWDC7bXvIuGFuIs/4JjSCIfCe9vc3FL7d/16huka
77uj95yTHFFMjjx/rHPrldDDF3DTv/JZzPzcjHdVivcKH51BE0d5Qe4AR9aG6heaoHObKLxITrNW
mHeauA5ve9o5XbuA3tTuELoZQ14bjGWjuwXlkdYJ2TlYH9qj90I7SReCL6WAwOfTUHxZbuNdWBZO
3Q34PNvLsxKU609byxGCR1IXG+X2gJf5XRUB9oouRnfNXmSvaXol3gSTYj/gcW238aLw++NqEsq4
qbshZuxJsX56JuIzrCg/rfTcqzII5ZVUnxl8OSEgt/LoHJEgFYHCUOHHdfHu8CUQp2bAGl9nslvM
Ct8PMZq7eUQRkSYMxOJiwWrJvjxEeyjYsmcMWHs5mXDg2qs4Bt2NBfKbpuBwJv9JqWgncZxi3ztt
F6z+hUYjtavtk5v6UnBDJcc38ks5Kcx7/OMDIn1cXw+3A9p16SIMNdR6ePZ1jvT704swJi7Ot+Mi
VI4U1QSMq+8+o8Vi0EW4fdwaqGp6md1K8xl55D5WwJXY+SHsMkbNuZ2Ez+VPGsTUHgVtI0EHHIt7
sznATLqBP0SHM5yCphTm6HQ7KntD63TPRAemjBbhBL4HZWp6MUFksWmFvsGeS2bJlrXWFGhFp4E3
JqcuUTfXGv4kjUwj9g1TBVsvIZNt7WKlAiyuYFk63DZ5UFiye9PKWwX9yfiSukly6UmrjXkQvZRw
e9vfIZ7W+aF3wzDCyynixVdwT4dQvc4Ps9Y66o9HKLE/A9mES08jhjV70AiFtfbBZ7q0yzKPnwbc
86hxJoZLMjMBSI+IG49TAniYJSzf4D/l7EV6QJ6CROUZYbnOiEtagQRTCDqxWJFN/gWJR+9ux+n0
clWmvUZDD+ELLgxiJechDtWl0FRbcVFH+gAPXb1wUW2yr1tTkwpmM5JaOKz3knU8a/Kh4e5VBk2S
9N6nMm4HewO8Az7tQ7yXFquqdfE2JgkM/kX0SHHy9cIdo22LcB0YVsj1dC/kHqOE+i5/EMKRBoeU
TGQVZbU6Vs+eGWQkqqGWLen7BzL8eCQr8I57PQnEh5K4VRllJsNcyNSxqzpnMTV7k0oC70IjT5II
gvNyGgmdmoVsyYfMDzta4CjZNfyL6nzJRkPQMWqnxtAIPhposv+hMDM0mO2CG7JvJUME9mQ34Lnx
D+nEnfberxXN4O2nTrToMJkKuCo7NO82FaFjTMGhlvjPDH0dnmq84U0QYFkdeXk3VGtQFA/Y9Pjj
sHfSJh7Ezadw7Ye+gDjk2bsQgDq2lqJdYztwg14XhK4K+5D+y4B/tpSeb6/eQcnqe26yi8gdFnSs
T7eh/z9GUFNI/3wW6ieTs8qS5eJ4piLvUqE/a33ml8NbnpeE9JGPSOh6gP9hxIihj7VVaG/3rmR9
O0/GpEzIaj4Tl+jYSUiF8mQhTUI6q61AmOwAXj5Ktth6r9ZpLNBB5vUvU/XPZkmYNH6L8n1S57oy
7lfi/Mx12PMY3TF7488nSBR+3O7Hqycl7MYylAHvp+jrh9s5iP/UNDNF31GnIyJiozOM1wcmoeN+
AqNpL5a7YwfU1zQ2hR4L7/PdH2AppSA9wF/5fvQf/ZIJW+oIWViYV31/CUy+GiVUvWiGelQ+RJoi
4J4IvZH1ekqyEizjMB6e1N/CrCwkBX+xzbrbRVmeadMdpQUM4TPnGyDkScg9eGowOl7Xlj4c6TIU
b/3NT5ufOLTHaA8kO9QqB/8Fw+k3sd48Bw2GB0CbcCmhIGtLDu4Kw5EUhCgmU/9iz3QRLPaCJREN
ENPRe7tHSouqv7NYmMqHYSqCuR0PyU/ZrbMdzp1g2gZxPqn/bdzBLsviB6HajyHcd+iiSxR3G2iB
HduZe6bABn53B1Qe/Y1wLk/dn2mrOkMy9N7Tza/zvC9J2IPPTLFUYUPIm6QeXW43irMuSP8Uayv7
i5BEmFjkDqY9Gmq3aaIEvD0/US8Qa/OGw4HP4dSSAVlTtHWdnN2x8uhvsbzlKq4uOx00c0XctfhW
tucVLumKflCmhAlfdAiX/P13qbTvMUrFfPz7UGvXrfypyfmBSZqDGopsVj5h9fCjhffherYMirgw
ijW8HNZf2KFVIHcOs4PmASQBNiiooW+F2+LWRnxo28EhyZs2vgdDKCjQtHJl7xULOrIOVrcpFR9k
AAyU4In27jZww+2z7y3LfOR3Xjzxgg/WEHOLDg2lJiR8MEBeh8BXUdfTyWTObhg9RgAJHqbN16sg
nQekbOXru0h25RmGI5nfrnaTWh/Nl/VwnjQK+zQlFDNdht4JpAZ+mhyi/olbUI/xk0/1zfZ6JzCz
AEzz80sa6bFGrfq7J8eU/enjZWfKV4twIR+gKOHd1ZHYU/PudFenST/VEyKOQP0z5rIFHg/Qor1Z
/DPHueuercnffzI0ymn88OmEjK4bWkqtQAg3FvxZF3pmT7QjFBisI17yPDxYZc2XWGusdAPzwlz6
T1nnUEfB9wv0Nik8oVb4tJZTz70kfXrD9RyaPK/CN4D4CBAObSthMxI/WJNMACfD83j1nBnk1p7J
YIRpKeHTQeTqcMq1RhthuC2h+AzXl6eqQWfVyJrlW/Ol+bIyQizwoUsBPaBpJoIzKQAhR8AOzWN2
fxkrsZuJ/DAdKM+NSHwpenYPVND2LYdzb8jfXVobb0T8nPbTRPZs9gbEBz36mmbwWPB45HLeZ/K0
fYVhBOI0pLdiX1o39eJVjv1axLT+w0dTMXqff+rpRAy2ItpG/RV/oW+yyW5QgPE0ostuMKje8URS
gI8tvO1HocnxTZts9wMqI0Q49Yg3+mqQ99DskBi1a3RKi+4kAs5qypvime2uP0OgtVE+NdQScqRD
gopEMRcNS/3UJCKp6FY/34S4hUg6UKSp96HHv+TkKd7A5Ow2eL7ztjO6ufeANFoxb7NCUkZacD+n
mNyzBOY7tIxkkUrSiGrtWmangLN5j72cE5uwJS1VNZ+x2ZYCxuAMmy89IGSS2W7XQvPgN0XgshiQ
Yqk91jWEI60WcAsR0ZqlR2kSzBMH6v9jodvCe7q5yK0KdSs3qtHnAOmWyerccYhFOCmB/DEEoeJd
67vAi1FgBNtlxnvwOazmDZyNUS8xOA9np7hFrdyEBRbc4vAqpvJhhNgl0Mi+WhDXMv1d1fZpGnvh
Gtz8cPbmoXBHqAjJMsYhHVt/WL3avZ4TjSXVLcbuR4nmpRkfdA1czkmXwjn/Qo3M1D8p1CpGso0P
q9e23lLvn+B5VJvOiBmU9bkcIwg4AWfUhD5eNKL9MoYV8qZtK7Iiff2m+E5PQpczOewfswKBMrsT
sxqvNsqdUNqmfHRH5guZFnj6OUbRDENkEJyjnu8x8sgLHkJxBNVTw4JILvjk59+p1uX9t3rjNVzS
iEk7pbEjT0JncGbGvuBQeEbkwjr/ECyRwXMQSlZSlgOD87vDIejSxcW9m3gnnntrBCZm9/i1ttaq
Bk7b3h9L019NyKZuWzb18q4zksSnFw4v1nCiI4ulegLreHGbDGkAYyd8+vEKFdU0tA9TwmdPUH1D
wSCIPF5W2rqx9U0H5yrgHeB9bcnzd5+Me7dYFQyu7Mbu6ZU7iAVtONR8U+0HIBby6lAEuKlR272g
nSuJdceGAGCifAUbO9MAGKnrC++BjE65rOACl/upJcMYRU0yMBBTs7NgNreR7zsQS/N2Zg7i5ona
B9s4jgtQgmj6XoFhLlza6CdOIrL5GPGBxtJfwFpYCKGlJmPVME2X7eTnqNgrZLuJghUdE3uRbFH5
FlvLkX7khBVCTcbb/bHov85SG01nZf8UARh7k4x4gMNWKwINLisjn+6KyXZSUGuGS3Pa0ZX/nfA7
U8TCjiO7CbR3GV8RvR9tCB640VLlALj9BWkXPMSwpTH4Kq/4P2kO5SnZM+azutm0+3iX8DFGmXU3
wdiEHiZg8OW4K047268qc+3cs0iGIFC4x/cFm97ufqylvtqDCk54WtZeiVpqkyuKX5Oli05PfEiB
XDsxrbT17eESnaKeB4tefPL0BGhmomzAhFsGvjtWPRUrXIzykQvqvdS86StnBPSmiB4LOg2o21hW
2bnSKBXlA4voRzfdoMSpI3tCJtAG6lqSTCvvLX33HSZfRO0bPXKlmP1UBU/iXBEFlTEieS/noWEc
rJFHNgTrwT+fxIGdVzBhOfkEIQ5qXqdKRCXjTVA/4lLVzCbI2HoOgJ5fDMDKRZvBnyyW4egEYy3X
8zb2fjNevCqdMpddOKN9MdSEIF7EXsEQs2mV7xVoYwqa83PcZ36Q9Frr0pzJawRCZo93qpYKeR7+
8nd3l6RDpL16KF+OrZ6vescOO39DNqExflhZZWgL6+CTffN9yT6p4zdQqYQs1n9Be7c61x9dbBax
ROYTrfvuik0TOi89dVhnTJw6jiOd0g779b97/y++44JKiEyFiKsz95IaVmJtzx6dWg9z57mJGHWm
i+V8A3VxtWaTc2TmwrxaQuFT4Gq93f4qvjPhDFY+4TZivjV0lax1ghQ8nRHm4cFvoprfl16BHr4o
c5v1LditZzLNkMZMFLYT/+5b9qj2+ADi9LqIPfAwfjy0QXPZ5L4C0YOxiSuTYhM2RuobOYNQdRv9
vIPkENyB+R/q61lSRNgH+WvOZnZwoem+QqTUZmbEjv9CN3JP4mCGoLZz/yG3aiOFYqmRP6Q5DRZK
ZTyhurHfCv/OeVFxtC1E5ztYxkUuH5oUrJY7wa4mX+76I/dLyUOW3EkrBA/Iz+D5G1/9cFov7Pxq
CJ1rP07tIZKMuVUPc2mBC2q1REPKdQMF+d5+XNQuautlvLMa2JGcVQSpfjQt3Eirgb6aNP9BgPII
0ZeIKIuTPhJfNQU/v1Smbz94c4i9gKfS+4yz98HTK3i6MUBqAOtG4x1l9g7z3kBOz/Nu/fpn5LMy
im1LU9TX4Lfbwh+KP3IDm4CSRhT/lhBIw8DZoQM0frtLOyUJfJlycGc9q/bvrn2PYftZTpHdE+x+
pRUhrE2MH91TmEwGHp7z1JA4uWbE1cz6C5iuqG12wnR/D+MueAyURcAbSw6p9K/M/Iyn2t6dFfSi
vJYMKaIAUm+gqVHgmJ/ptVu6wNqJJSdM7upCZpH1cM1AYM4G1Oh1GEB3fVzwytufUuD+0Jw/jV8e
+7XACQoOgBLoDbeuADYTMCKEG3wwiA2mBmvoZSTEUmh4WmEmQLncWIxpGGFDFnGiu067ydmelnVt
5nkjsLXsQtT5FFCvQDPDgLqzIm/pp1GQG6vk0krEk0w3l/cjv9ikdKxdVLfUR3y6vsZZsSPJJrhB
m7EXvQxsLvT/FcXGQIveDcLAE/odXxH2OWnJhn5ROxgaRBXKgQPuaxDCY0Vew8OWskS+YcIJIIZZ
ut6sI9nFHLc+0LM7v3Nx0jq8rX86MA2ay1xB9d7U37j7ZZ3DWlz9DwVqjR8kqYpQpk21yzvFcoes
PgF6AzGPHRwmMQ7C3SGsNdrFvpg8wQqVr7Mw7V5KRZPappVTxE9nt3kKeIk/jGqmgUcwiHPPjQ6+
00sHl/vuHLVI/zh5Pg2BZhHf7biTHpCZNFTZCUv8LAYuZZwHepvTHS0kL4LL6BhV4LgxC2SEsSjx
DXvJAhi6GqlGV98P+vgLoC/RTHxEn4QknsuiTJqQW8pZ0/iRO4uVtv9E9oBKAzIP1Np+NWi1GqDU
kG1jtTgzKk4WOiWhWfoultohVx9x0cRef65zgCGtnQEx+Wq8/K3dC/I7XubAtsSL3Oa1L0xjAjuD
z3qYhp4ItrcrcastuCaz9NZ8e2P4RLVuel9ZJ8jbQCG1/hxvYhD/4OIiCPv2cS9F2eeZA9DFVvo6
CZQpccWoSlMc/aaVSotH+aXdepNpw07iQ09ifjN7PIYTYnUZWGYQ6myV5M2R75uu+6X4lMJaMUO6
P6PaWOqDaqRrbXSagTCZ4f4tzj1ZQsZtAAO9I39zNgIxW2Laab2Do/5Q7qAdI7jswMZ61tcNrCgL
GVxiNUy3+x95bdd0f18g2pe7geu4CW2oVNcYJvosjcv7r1PXxWcgC78ofJAgRWvFMSZMHT49+A7w
VV4XdQxa13sWseFEb+lmuJNethkHlSmZZP5rvrHw32D8jg19wOJxJCR0Y2uUSeJCu0RG72vQZetZ
WTQWSBsYy4EQf0o8u52y1FFYFrFTvUNQk7Kyte3FlDFC5LtaWmelUNlDDoZ3/h+WtqiVWUceQOjK
YfpeFPevOGnC+m29CFd4jsLB9r/lpderBx30WpGdHG/n5aF2lWf0PRmO7HKWKp+1hbfLk6bvYszQ
xrJp5i/cFq9r+mskgesQKIfWyY24tr222WUypg4/J+RvyIcWWmtV/nW+RkMlWjvuidZux9jUAxkE
JgeGOBjhdvFLI0mHc/Swe8wpIBFO69RopcvdpVhPXAv0ic3i5JkKM91fd3Hws7YD/rBELhOVE0Ej
RXacweWV3ntMqdsA4B/aM50LDy/+759HSA8EKBMIpqyPuSWj1qN4QeMqMGxW+WJuRrAfZqFld987
q2jUXm1Um0Q6/3phzr5yvrR0YoBSs0WQFQhXx91HgE+TxPfnBG6WtVLO81CKuzKq4LQIRrWMMjmd
6nBBJvFlX9N6tgkzztIEVX2Pnk4UO2/dPEroTHkQPeQfTYx9zpt5W8P+u5Hae40nDNKCijtvPzVi
+lidvsbzm9DMt5STa7YasjIft+GjXYpC4MtmTQgrxbNc8Ekc2uc89VGRqzVYuezyMQ9rzbH6ReOn
8Z3jyW54iOCpJTyc9sJ5vEgQatdmBU6/Dtvfi649KVn2SoWeh86ZgF4lfvigoL2wBzr2gFPF3GoZ
iCABR7qvplLIeUdnFLFzUgvW7r0bvE3VRvcym4A4sMPoFbC2nvh2jaP8ur98zox6INDsdrBgULXY
uX2Lq31pJGpghcHgRiPNf3AJ7NJtmUqb3b9laA+58nSYGzC+ca2TmPvp5hMS549dRS/gVqMNqSHV
vFaOq9y7/o+8MdXqNSCyU1OtPZ3OprXHR46RHkQ7HMghvwTHeCLDLUOXh6Qa5dM+SbIzpmfE/PTV
Y8v2LR2RDFDLs59AT/8g5SgmTSamwwCCw2VsCCdGwuq7uPSh/rBZ1BGz5DbsYsWAxLamdAAHxlnN
TcdPBq4LYrLF1yZiwM4jpx7ZNNtwTxEpCpYy8LpULpbH1k5MnTKH7EEcpRW9nvWBjLLtC31RrgSI
SoldEqbNC0DsTT4CpRmK7cVW5F62dF+YX9cYXI8pOVXKUGDkqXg8LMQoJ7lS/bN9tjNGxr1gTWp5
wYXBfSbL4fKs1U09xutRaQzf2qLW/7uUN7LfyRYIA9WNNP2f8Orbd4QN/YviGGCC5Lr6shbWZJAK
JPdOSP4XjrgJ2Ooww5sdFGBeNqCrxYc87ChH5V2Ko3rP7OojrOISieiyz40njYFfqSni2onLJ2tC
PldYS4Tjosoh99KKKbByFD1Vr+3+d/7AKg8pqaJo/Qt5OZq7BnF5uk3vsoP2ns/jm6J/p2hi2qI2
b8mDwwnWlT6wrYxvTCdz03IzpiKVhdkKlXs3MBmeXsgVEo4SzgZ2D3Yv/coXpfyBsuSft1gUO97K
ymIW/umkRnUzuTbXl1ZCYf1Mbtku5UmdFS39qjqBMpL6LzCOJhOMhsZYuSmLbaLJyqH5At7+1Y6k
GqA9ofjNZv9qTjobh3zME3ukdxShun/efjyvlyl5kq/g7y/Q2Tl6NJSmQ9t0UhhNB5y4DlIeF63h
Mk2TZGuBioqB45kKPo1YEpZTfS2L6p7rkmQibEhnXtoheQ8PcNux0uFP+qTgLt6CHvLuUpRKN1Ka
nHty8CNpR89Qht/gKebb44Phk7c8+HXXr9druVQX3yHY+McqsWFQ8Pxi29q4sANCSTGP4xm98UE9
wdATww2rkz+NrWxVKr/5MJ/NotIZ9EcviSxZv9Av1OMRngZ8vPW74iNwag2J60WLM7LYUA9/9eQH
r/w8rHlIaTctIVeN0eR9kvSm4CYxm3AMJwEj/t4e9mHifKCzrc07QSr+PTSSZhoQWqWok6S0JTrh
96A6yubLXfzWiSq9XkrvoZA1muz8I4Dncw6Vl0i8yDsRQ0nwcteRrRLzrH744q7gzBD5Zvm3GURo
jOhnfxdZIz50lKxcmDT6V6J7iRfASlt6TScV8zpdxb+MgYw4n4X1x5SOJq6mClUiMVV5n5EJWcRL
Q5eODzW4Nbn4xf6gbEjIsN53Qqi7V2kQ72KpRCzWdnGYOscdUMZU1WsPxmAIqyFsU87JpedPMmXr
Ca/iAF/8Y5byJx0EPPg/Lquy13iPwenXXmaY5sgrX/SUWmUY3uqZ1oRI/BjoREB0b+PqSns99BHj
KDKAQMcnHtL+eTAhJqaMzAm35Lpnffi9rkz33yIUWOdr2Ocpy3fOLpYVa3bApdIOYNSxw7dyMqK8
PCkZ77URdYDtSnfgDVGe8Zl6Nnf3x+RBRZhRzcK4ZFjddZWSjVUJx9EFO5OhEJlu9yMXj2jIoLde
1KVfCenWSWknh4YZkLDeUYI/wBNqy+eBl4sju4mPYqM3f1SQ6Hu6Q58lT9m43kcRV8d5me3FGTWk
+CT5xc0AU1Hk99cMuHWrI8S1v1k32lQG36IkXCtgW6uj0Z+8x3TWJ19/6gXBKC/ZPi2MjuER7PZF
LzUbkptW5W5V0APiJR0geRARlXEqzkVYn6d1WD9PtWyHBJ2u3iUFfotr4p0jxlMXcTnrK2mJWN8u
pkNUQ1TZgrRDCkGLnlaN0aHLTvCB4PhdgCG1soS2uMF+9eAyBg4l2D0YsZ51Fp+j9XmEscnAA7Br
kPNZ9Ykngoid43br5ZyFU6GrctuBNKUdneKy5qbgMrLjqNQDiERENQcxZgg8CveH71Mw+BQevgNS
b3nIDI0Q9Xd0HNi3sU3ATbyxbGPk4g20nMJaA6kylCrjxRNPO3J6uUa3xhg7fLF2Nzp0WCWrjuQu
Odou8NTGhBfscmz99MWnQ+lNSemt3O5z8JooATuGDjMIL5pdHWT7w40yyIhPqzH6CaywKvaRwPmZ
TGhFIGJveACCyC8k3BzyCqMNACF2cRIPboMEZ0d4JigDH13ISYhw8mYMplawGIYjGUcCo8t6JY0Z
b/Acd53n8u+wBicmg9iO8EQPzf2EPHbKvdUCZQRE4duP51tNyaPAaploUFFNuWQc2za9M9T/4fWY
E5ohRSRnqwthny3rXds0mR45wkKc4KdM6wcZFueE9uJECcP8krPjZoVjeu/CuTDBBMaIxX5DiyBp
9UAYZvBluvGsGLgtIaN8kz8MFHUVugppHP3xbDxETU0EAfBfffAPyBKygwxPNR2kkNlOwbV1Ei+d
+NKtv4YotfiQDyAAQ+DcmKpRbfOr51+Gz9Qi8tCGDiqWHuH0Z5d4fHguqKfLleToUD+1loHDFoFi
LTS2bpqcYGfWFKfos/D+ewtV3SmZslyz+0ULL7IGS07e+iAQ7QNAaAS0nNdwW3Zbd3oeGzHYLN7E
buwIqbLQFPHO4Z6DTguStZhV1OVjnTp4RrDZbLIsYmMsut3pfDx0HI+/b1cdjHYvFgmFRN/EtFqr
Fqwcx/cSMH2jOtq3TCAa9WAhaEdFXVz8Djah9l1zGiNVceKGl4umLTsmkbATSCJgJF9kINo7mfNR
P7/Czy9hQXwIho8Bb2qoensSQNEMmhb9FNhrWHaRMfWw7KrMcnd6FURtWSM/x74w+iBKQ/tb4sS+
p6jTgN+MDva6CzynCFbvPTQJuc3vAjqA1LeiPMqlzwjgIGklksB+Wd1bIkI7qjZwA90k6Xx0onaJ
C2VKS6WE1I/eMJB6hVmWz0jqqFGNieZi1P6srqCQf48fgfvpfwiaWrtp1y5DFVuY1l+MomMIrd+d
totMbWd0Zx1ljuJ/92jX4Dw9O0v2FsEjYSxLgR0BBCx7nSZN1iagKFEmdA+dyxwOakxknDATXv0O
zrqt2Za6gsv/1FvD++52w2JExK47q5Fq8MlTek3hDRkXoDBvJlg738nWNwN+RvLNJzAYAJwEtGFs
ErjQyVL2ZzsBrfGIlJe8wxSIDBSGonb/M38YtNebdLwrEAe2tR/KGt1kvq8U5owgE7BbuMNUzFY0
AG8x3gwmAoAJESEwePnajDIjjpjzjDZ8UrVmiQBVULYqLYGpWzRJfyNp7b1385qTnTMtnJiSAwVM
o0NVP/ot833LO4jYjtRYVZR8mSzijSy0xnSenfvEBtTiBwRv9XBU1tqNepwfZ58rIkVEOla09LRk
OrA+A/Zu2gVcGz7wNWcDCcpq/cxS/wLSR8Qu7G6H2pCav+GmRcLK6icNjnRz5fcknoWXDzdYNkNt
Dd/TibjOgYH6OcF+ayiz7no6lB3kNNWsOZ2NJ4wSaQqnjgS6OoLAw54mjEXQ0t3tftTf0po8yI/2
kqmfN0T3BXiFnlOqajczVkdaPY0weqqJiNwvPdEBdMob3+dPc2TiTFwvr95KyX8IDcSXMq9KCtT0
oQQR6JX4NBGYLtCur4Y+VbEMKBy9U3u4cCh5fmG/u4lPRUwZ1BeWV6gw6WelsMZaXJUvSBxdUzU8
P7LBx1gQYRdgn0e4yjWwpbMr8XR3iCZ7kq6NYu8lxchXwbTSgPEJyaPGMM4Ep0n58NTqPee4QOw8
+ecNSaWlUB6xxWeJ0g6CnP5chA0Qj6Fsa9jaCJZ5j1bgoztI1Q9+Z/ZZOYHWvdweua/D56U1vlgH
iBZbY7Dbb2pmGOvue1LpCp8uA2Fll6u9tMPX8bVpvHGsEIRCTTSUIbVX/Mgw0kElRBb2yYsuGsK8
RQ0RBDKmQvF3zbnI970ejFfB0bi3EAxcpLWDfXObjQa8iSrU63rM+LWdtRmeY8MqtLx6wumWK70h
/lAZXcjMGF3Y/2vWJY6yENEBLpL/03EEGcXTsmM1jTbOmYurVBi8mnlRQHwUolRx8eBZ5c75LgEx
6nJJgUOoAzQ7zcqzDwCnkbm7XNivGBJi+eEBOV5irWJo2wFEAEui1JWiuz9i6lxIIQol7VoSFkpm
igsbzYJbTp0iMUGgYRj++JKj5vyNLkhd6/3qkru9QxyYG1AO2vz0gi7njjhIFaKyfMgfCp5aA7Sr
JaxCXn7UEtYTZ+cEkSgJOBXhymq/xZvqu14UjNa/OBqy60o2K4op/LlUs68eB+Mw8xrB36BZyjve
H3P6ZnfCE5KpCrNOgtXbpyCdeJAwt7zzNDMTuYfhi5s4geOT7dB94ZfgKatBu6+erMW8UCPIly/s
ALH7T325hNWIA1Du4JxJSL5MxjSKHtrlTep00I06wxQb3eFsQS+K6MEnrKqFPAPV2hkzdVNGFhEe
/p+U0jvdMzgA+o6aZI5IjfoTNvsvkozyUQBUTm9dI1l5sEkc2Ukn2KQVeFPuckZm97XayHZnZOhx
+bBNBM1cyD0aOpmNmzVXi4o/6Dfq6hsI0vbLVBSadeHD/F8gHV8KBBWpSjlqoSlSCOSJoFTfJG/h
CDHhVIRsSpivDDcVUlhs66Xb46YUzLvhHt99v1FXfZIHmUIulWvQY6ZrRCCzupT68lFFMaoIhtO7
tFg1x6dXFoBl7VHUDlN39QB4UjBF5eG/6MMck+U7TGddLkvGZBDC5T2MmMbxaNgCo/jSolwSRI0u
tzC7U09Q3XT6mViA9it8QjS9J2w9rukIwvGUf68e299tfx791JQ3ZS9QzTXlLs0YtIS9EtUB1LSn
RrroxDy07hSbvqtny6qv9cJ8FDnq9bCG8ahkti1kEIwfYeU69LoUL4x91ymS5WGYEG6e5DAq5rd3
s5hOEQ22FMKUhImYIE5tVskmt6ubO0xtPmw+xFWNLIprPNnqfw9p3/JSHSbuP6W+ny6cOECd4Vsi
64ZabbKKU6459hc/Ca9E8Kfm/cWuiwoMUnEiWjH1Vm97PlEs4N3+kwCW3hJdo2OgAVgVAr8zyK1n
dg8eqUMxBDcwjPLEHMHO04LjNzDpv7po8z5sjip2G1e0ShcMvdgF9lpniTBkh+SF7rvtT5RrlfMx
clUUqzIW0rp2Qwtyxd2bUcWR1VzfQXlel9BWJEfRnQ1coIWEJRSSZ3he6hbetqXwnOX+75YEKkTy
1wjX1m2cTAtc4ctEORdGBB/By/hTBwpN3NzCTlL7Vy9Lk6Z01Itkh8Phqj+gP7bHSfwk/LtS6ohT
KikQ3YYVYgjNPjyNftEQ/xU1hlQp62pDTCiV9JdzAcJ8I1iUu2g7UQ6Uu457TOheplPQKU83wSfm
zBA0qkBitkwWUftK3FpheK+m+fP23jfTuTeSlcSUmsT3K7lxX9F/6JCNwkFx/0XGoH6YKW36RKJt
Z3je3qaM/Qo4+mASFGtbwu5JDyMJ46y7JY+XSojOJQ5UhajCZh+Hf63bHgWQ+N6ChXRJiY2uc/kE
o0zr92KrupTPfTOce2GLoS/xTMzw3DY/Zy2/bfxar34DCOD17hzpMZqK23HqUJdAv1WI82zX5NmT
n7nrpSvVXfZ8nfFrfrvp3HiavV9zzmu9IpEX/YCH2GNTmhdTFqn4AhMrzxYQZPPK2dlqYjyegmVD
Fs6V204o4wZPbQnspKjMRnW6sW1Wl2xoHTU/k9IPjIZ0buPeKArAYZarwSFGlstblscg87JTKS+e
1q6fPaEpZGtYGjK/2C8UPbWLn+YiaOoCZNvRPCTK/tnkPke6PIPio34UwbwkYmOPpDgNJaFMWoef
ytOKVVxzhM/5Tsx4GW7S1sF1JoEbid31fYfvJ4/FfD1qyYcmyeNt9PUrr0Q/VXsy0TGSEL6Gged+
8ieHfII5QCs59Vl9BoVohCxKcByRorKIKtkRWdtPvYa39qcYgIG/74Bex+g1hvwUQD3NOh9HPteP
0BlnByghBsUsoX41+rRC6pfo5BwO8sjUvH0EUNswFaRpNI541Y7xRDE+1XCXwliWQ+2ACyR8jCbX
s3RGTkHZCWYCguP9OKx4m2xAH7xqJjQfqsOaEDc2QNV1Vrhuq2jpytPuamfFGPM3dfz5ISr5ajbb
60sIzVP9DEMW62WiUKvSDeg68EHoXmnUOMLwlV1OuC7fMIP0Ulhb815UgkfvpLcxGLxlP2WLiCZW
CIgTxeEhtoEvc5ZgFVRtl/MQQzg7s3Pe5lSSXFfUQczvBu2cQE4NohOxLRoB+gd2Y+6UG916G5zf
Pgb5Biz2ABqwZSU8NEUjqN9gYP9u5ifutmwX4M848S2KRPNZ77uWPKQ8C11ziEQ781hLKRr8UZ3i
5NhtKC4rsEkfNf9I/WZlGmr1E060PbvhycKqsuoSMRdOijG+peqXzt6USyLgRIMWCvH0H9jvbgpI
3lndjI5nZ/VQTqpovktnkr7fiReXv5zLyR1x3703rAjDB3zBx/4hpouagpZ/40s3YAy2pSDQplo0
dwWU2ujlitXWMyJx9AIas+skgBFeAlTg24y0eIWjvB0hlqtPShcDgpiKb+xN40SbBa/YdODcIe0K
id4n+mJ/0OpG9LUoHE68c7VVCGrIC3nD5xoQ0A0jQkDVlUBk1RinE+wI8Y6H+TSWLif+ZsWIt24W
TGuwJpuOAh3Nh/k2ZwpXoBRvyD+GjHZnrOGo+mwUwyL6loTFzcL68RvKuUiGaTH73i/CIdEsykil
+b2hYSwu93ARwLDz4QA1Ncmkayx8ZoBCiGYqoHuwYaX+0HOm4GUDnXVFpiNVon7965Ekgmd/jvwF
Bg1rHenFZleyIVTu7tfcIxLFG+cq6YmaYNGr5M9fe0sY65idPAQjp0AvNjV2bQqKvC82b55CujD0
qDv3fV+1e5FEvUAG5GTyZtccgRAk6Ey+zougJR997H6CzG0Jrhh/2orPBORE4lhG8WY+R5Cl8+yI
8GnIRW6OmlJfidR2imxum7tu4V0AiN2JB0zp5werIo3qWTE0p7OM3ujxjWOwE4PkRvFn91mqsL4k
ShB3qKBqtfLoD6w3q2zpRV54V9hQWqwZIwtEnvfxzzmARdp5X5v+8UDTu1zZ0B3j3BznxM55Vmvt
Ry6IqNMqC78nHY3YAuK4iZ6TNDaNPNZYQ4loLIYpjg1lMfDCMmOo9BTU+lIPmJGUzpWwrF5sI/+/
VszPyZ+VQ1fZBnvjxpNcVwdRpFY6YmNKmDR+OvO5ACiUR80z6Awh7E+HIOgaqqct14d/6f+lqUdc
dMzBn+eflm8zdQk40iDxIEJ9WFSm8Fme1R8V/22R57RQJ/eyYfdBmGFIoFInJUftQSQrzuru/hgO
QLx8gjMMVjfQu7sGl8mfPW5SIYRGIvlOIHKVljiJ4647A/sw3n1QxW3N7CkofxbtGuqkJSx+Nkho
9SiDwG7Nl9xt/5IzZVKIe+HGNbx2q/v9ndf9cu9zawMFY+QtSVxJLBgErHLBO1RnwVCPATBzCma5
xjXj1TjEp3zC4uM8Pz0NliD/ZIRJpS9fCt9zrEP83jDWatzjlT89ynONJ+VzfTqWIU0fk84kfecQ
uHs4m8UdEp5FUziKDi/YoAgmY0CFJmeW2Uzvw1lJisXZAt7qZc4WUwI25AlgvPZBvRjCsej0pxVF
icSS0Piz1uVj5nUytGY98+7dfL91v+0UIBh5vY0iarXFDmxOjlgx6uBjdpyk/wUbCgTdQYdDr4Tk
ytQUcsp1y6YaewQ+C1QHsgI3mIbkVUoE9fu6D7UvggfTHeDFtipfZ3sPq+Zc6Q+NUV0r6XoUWnpG
6ydBnxyuvndyePuodYKhVtDHHd2N+r85q5dzp7S4P931NKE0BPxeXgVtMLnaF9KhjxaBI4L3/2au
hyAqbW/f0XXQvRey/usQtTh/adftSkgsokxQcIdFXrf/6byWc/cCrB2lAJ27Ic42XPUeQE//Yqx/
UW+XAZmNTFU+k8uSXLeORfKtA12rxGepa8W9ghFD1ANRUvhVExwFEtrZqIVKoKiSVMV51s1EX5ZS
iDCz0Xps987m3xKZpza0iu43F/9PfRyEqvC+Q4fOefseDw+nFTXqFMUiXOzLcIPpqH29UM4nzzFS
v3BdFGjTjfBmQH6QtP950gr8fFEOqAV/jf8em/qsFpsuOww3wYzkwqPiIoPllf0H0gfMmOgQliyV
yCSn2P+vDMOBbuZmPU1xhPjSqSnMhdXPe5Og62CsgIp6+59XbC9SDsDTxEJdG8vj3SsNYfPIXO2X
LkNN3H+QIo+Efh/fz8ZU0Spv8doKanb3uK4p41MApgYYhQUkmuG4F481qRw60bnt03l1HBMr/iQd
ZcBTGEAE9Ibl7wzfPhxeKaif7zE4PdA7Fn4Mr5/9FthAfrFEMqBog8E18BGwUSJpJ1heF1rXDxZ6
7A+MYSE0kjIrRtQ4sE/pUV/oMRU6Eo0x+B4sdmekikdAA5DoCKwXdoJQf4EoQSnEC6DeSF3yI9sS
IuJ7QgcBYyQRp3ls25IxFtKrHKion/mqLHotp3p/Pfz/hL6kp0s0lpnH9ItSUoodM4ZyqqP8MV0H
X66hTS+meR0VQPvCAR4UJDB5I6Me8jtHEBYVKjgWJ80OjknNUzEgOlikPNq0yeTI/wWo3kq7DVaO
PF4pIApewccT8bUFpE9D0oeCh0AVLpyagElKYsRSFGeGPZ2pezssf/e6FIAxnQRkK/bc4voxttDo
Bntb9gEA04LyXcBwFlvBZr/RPVrPVmCZJiJkSb8N1pkvt6WvglkQI/85GygzbvbbsM7I1nObWSe/
I2opalQJr+nNi9Dab5z1pHBcRDSYYTwHgY+hkC3mM9S0IbS8Bib3TUJhDzYP4gUkyZS1+VRyKpNT
86WgDBOzVDMakFRs+knNAZj2setWQScNsarsnFHxPH8TGfk9V8MgqzP4zNu6wOOe1t1oShPlkPmk
za763r782YRXKsj4dN3XRHgezBI1ATltSXhvC3eoqsdBR60m0d669SxYuvagN7K/OXmVd9i1vqvE
4dpwyLpkGiBu3I8QqA0LvKiq8PZUts8/JRACJZe+BELlJCdNmCXcuHpVncXM393rHPmHzzRPBuiB
IUHebxjxgMIq2Qp/a2MXcFCilvFcvSMDlqCixTMoZsLcgMUgGrmOjG25tk7rleuprZBGz7iLcfqV
8Xgj8js3rU8nonBQ9MdBNdunpP5GEveBBk2oe3nEUK7kZiPF8J4ptPH+vJFYv8RuRaGiX8n0nlAh
AXDHFcWgHtFfiF6/e5aUkgd2yn3LHdZ7naoYC7DyBHw5IAeB067ByzPRFACyyszc1DpPd33nB3Wt
0Mmi0yQduAe5C10ozXrMeSewP9Q8vDB5aSmSpD3sl+g0VbcGg1uqxOO5CxIIe1Q+4pQnoBpTudy0
b81d7zT1F01aQMGSl0xrup5TTuvgZADcCMdo3YkdYsx0YRhTODcJ+uethHd5hctCSBsG6T7P2XoT
RQN2nYWGtKLkE1TSHcXd7RX3zRaXfmPbHm66wTJTqKi4sNjNAOyKNaKbToKa633qiLLH6eeQwCAT
I5Pf8nyTg5RHawJgtg0ifYfyaGTjA5JaLB1GoeycHG1IzDz6tMr/a8y2CbbNMg4+tS9VrwMw5P2X
TqD0es2pYQJsr5/4Yw6puMJhOalyriIowO2uxsD4PjG4syBiHP7f2nD8rIjJJJhoitpT9ziaTwRB
fcEHHulZZF0HxqP4HZi9UxLrOtRBRBcBpF1YjsqgiOz2MSLycgnoE9FoRzmdcySkHg/ITfNi+ANc
xj4Ca12aaQ2VWlq9f1JT2W02HXpzvHiAgGGv1tN0Nqx7H04M58CHUvCS8chtecDCW6WyA18HSlaR
6Y0Lt7ibYAsLLmME9JMSi89h0xMOobu1CFCRBOhPYwRsXkyZUy6Ku7TB4yxQZwMuUBcFlhZjO7TK
hewTVdQZswLMCWgzU/4XqWTCxHDClZTABZrlWtekBAqv01wpgtSu9ETSOUsXjZq/6ok4I6P9D4IS
bRyVCouFYbZB41v8SIspFLXdJ8SrAR/4otZmdTUSuai5QaF0g89vG1OTgyi9kNfpPuynL7LupWz1
n+JqRFAppEUvJBDSmVKQg0RmNL8xuJz/jeaH3qlon7wxuNoYgEt6gpLYBsJEp7BP7SzCmExZ5Rcm
dlqSEiJfQkAQ06/YprVdYDaPb2FDZVkOR5B/WXHph2ncsOui2+QPj07UAMunnGwqpwQK+E6+P3vN
OUAvg9IelOBmuAJpxj8EHnUexoZTZ0PKF83rRaJhwoOlx2pmQeDOdMgWS5lOSNrh45VfQ2AHCDXZ
K6LgLp3eK6/imMn1acJ9CZvuHEqqs5r+pEwcywTA7fwP+6PtZjTlWzmPyAQ4CcV1GKoxIlj/DIAo
uFplxYyXNh+EbmVVrfouEm5/mBVQIrawmNEIJ/U0N7uMTt7y6U/LHBk/khWxQ+accPAMu9qju+GD
L0XoY6acTc7v/hq6YDV9h/WSuifFT+oo5UcOF5PLclh4DUhkOMm/C1RnvpKEdNoti87jLEDBtwgL
LLrBn2O7mDuV81UdMOPIMb5nC5TXwSZSfBqXeRAN7OlUry+ox4UXuC/J9+L+CxLIv0f4JrASj1WT
d6YjLHa59XRXf8/8rwI0o/Hz3/V9CziHhhPEkoz0YQiiGn8bPHe2hxEA7Ry2kFYP6rMwY9dyj7yQ
ozjvSsMS541RgnG86N5LSNfvQBs0Sw0ZCTsinsADuy+onLowAps7OH09yKyfcvIuYbg4QZ5SgZ9j
7EJSfShMsb1om5xjzlvZ+sea3Z+VXig0GbNk1RshzP1Dzebf+QM8qQ4YdPjwHryJJg2Kjf11CAsg
UozFhczK8/WkmmlpDWwD/4VQ2HWb11f3A1TpVtLGvJwQSrkv/hVM3OKkbknSxBeRnTNlyQFLyOMd
6uBROLNmlqiFPr5ym/iRvuZZkSSYid1PcN5Bmw13w6qsHtR19kv2yt2dGqAliZYAIycZvMGAVg5H
Eg/PzBVss+aCAnNa7dlxaPNn8azW5YzSoGKMgEQ/rMTYCnKMsoi3x5hPSsSxVDibqQ53uHodoFuc
rp1RSeQO4uvo4bpa+0WeRa83p89rvYJhBtpufBF5+Hq1m9STRifs1N5CejsrgSJW+Tro0q6bIcCg
IlYW4XORsJQXJ5Xd5wn5TVtmk81wuMj9CGgxksMeBO7r2ET5er9mP9SOQp/o+I4UBBFy7VP5fmK1
+8dRhDcnCYKfEqHP7gjDzqgooH9HXH1EM7x/hrc+bxxxsiZojPD5fRcGRncU4i+e3g5VOCTD4n7a
lKN7KXdx4bPo6irWz4U4RITiM6gjpqiNF06NhSjXJ1UGBy9ZIo9PBhG9gP0KBozZk+/jP0acdXxH
ttl8YfhIV5m3QXxDj9J/vH/Fecs2OutNm9KDofhUtxn66XcF6qE3oF6P6jVyc+xnqOIp+ofwf5zY
rRdYQ206U2isMzSrdoORqdwwLE/X2q7C9PwT7YA3cdxgHVc4izWfA+hfWzxdCd2AF51n6Gc21rPl
6Ur9UhSiHKfa/Qs0ojFo2wVRA55BO0Ly60ezTc8iy3aUZ7kgMc1BM3XvWczJJavn7elVaCZ0tUon
8TB3ztdNgGQN7h/rgiPYCBdhevKEpT+Ez3kRQ6yHDMGonOCvlmNMxYyUntZwzI2FlOzJZqtmT50z
kIpFasmFX25fbyYWI7s9nvN+vef7FEeNB5UIxhxP9oQ/CHuuffoBjuPdJEjn1DTu20vg/+tOL7LQ
y+ahy7lO5p9DcWHULXLmARRpIcX5WCoPXyYVI5xo3eKgJVyHooOotR9yNwSMcjSQN0OHnXdU2jaM
99FOQuu6ewF+1ogYjBMlRUbyxeGuRlM2WvFkRtK86Twj1Sn0xQ38quU/bky5s+RFBNd65S2aHbLF
LQe2hkZVVgSQCyrn6/ajBY2H7FYRGylY3WXs0ko+QvsLKlGO/a+rU5Jyy4JYBDrthZvxxVVsXpt6
8DYKaow8QSTcgWMGQGp1+h5NqCUs9fmOGz36OegWmAkKVpV6RdQlgF4RBR0wFThAmRSBxT3JWAus
aemWoBVwR8x3T5mEpdnO2AjTADlbgfIuBU9o4ay9AlDC2wOVs8uvk91G96Tn5VLraeGJtOKTzD4e
9EULl5CeATplZf7aDrXrWpf37TVg4oZQZnpmvCC3cyMmaAk7sfpQyhw5q7UtcaHRhz6/Zg2ASnAA
PRB4ZNL3qo0htOmET/pxcI2x9Iug+hVeIl0L89234+okkdUsSGfAu8Vxh3emjqV8ff516r6SbGbT
Bq1Zswnyv1XoeqE5HEuNiY6bFjtdn3xPpkcQeC89Tj+kYgulKcQoBxDoYGoDB8cMS4IusHBcXM1H
UHzQiVdffBgLVJCoqJLrnSv1tfrgeXFbhFV28ICzdTy8Bm5KTFy4CK6Sp5m7uRPxkiH4FIfLsdhF
yFKksMhrpsucjba5AfPWPrwk8c4d98eF+k9MpMi9ZpIPQTM6LWWQHeTcmRCeT9uXl6sVzTU7LGch
+5dE10AkbGErMs+tUUN9z6LO2F7nPQw4d4PMzvEB2SNpSFdEugP4jNzS04zQZ5bWVltnLw81yeIt
PrStJmxL9qDQIYIJWu0DkLJCz4gosfssJ48KrNXx2v3nhP0gaVFResZVQbt+d1+aWHFmbSv020D/
bEJNahfms8mi+XXDFNPM6YeEdQSx4PmO8mVIQ6qFTFkyyoXKnvU9AgIGL6/RzYrpSwNRLVuJrTCP
N3QUqblCrGHtSczJjOlZSX+KpZexPp6JeF9MvwKeN6w6mNxYfeVz3XC3veu5qKoIT75uw9gsyAbr
xsaoDifAg8K9Uo6vzYS/t+4fn9lc5tOemGzJulqwBtCB7H9MrcOkQo0LYzuBi7QLunzn7h+Qjv1K
ZRxtG80wkE0S8DjFsmiNzLBBwr1YeFw83bePxSomeAdMdYClLSZCHDvn//8Qg9Fb+FDWMVYyXmli
EF1mW1QM3c4dADInCTcNg4K1gZnEAo2rrnYsWmnuqUrmr4YSxspWusNnLRVDj8qQhG9ZFxpSp6SI
wMgRuCYPBk022Xc8vXjAL7I6KNL4u3EJ0gkl4n65OJbSQMVU8Z0ITGqfy4ZGDlmz/PY1nqC3m9oy
YvkBK3kR4JYJlheV0IcWq7xiHp9tTDbdNRoIYKm44ooHxAwWWDB7Qfc8EEZgem+F0NiTbDEIfrL2
CgD0V+mbI+8HK+0ss6mBq0asxV1CnsxOtiE9zdx+cGYe1OnG+Jzt7bnYCoWVj5l60XOZtr3/HW8p
nxaDx51hqfq1jekyPnH9WW58cJAJAQkAV+h0m3mIzBIlBiozRkiG9jYYJw5glAcFpTMvUCQttY1t
abKiOXSWyo11o1pUczjzHs3+U3JbCuUTmp8/AxxaCTEGQkDAuJ2FjUUjsi2qHbvCn+k4j7rkQpEx
wX/cfPP7YE+2QsGmaiz2tygbtid5o0wgGyvOiBSLJNvmSWhQ+0h6FWjJ240y/9a3/B0B/L8hYMaK
0N1Rj3txn/kRoLmt5/MDyR5FJ7+U/4UfHNyiCsSI6c8OGiElDL2CC3e3Pg5Xdy8j140B7RzJsgli
TPKkUQlS4ehFMKzqHZxuwAhXmlw7PYeMqErzDcqllReGuauqEA0N0qCwCxkx0EWRgp0tMOLIkU4g
E5l1moKM3fnp3sCnuSEKTHRItupLzPjwAy28smljDzhvkMDwcTVoi2iUFiDLh9b5X+T+eI6CF+ls
IRgG7hVCQTt86muDyuSdY5X9nGnwtME1KFV5CLq33zEB5sAkfAIvS53S2tixZNlHvXT3c8zdO4+w
/osogRSvNeTmW+gcsaAXL1dhqNegY5ECPumuCUBW1cvkRjypD1/dJ/D8aaGYTlOmwXEQs8BLjkKv
D954vxakd4V+hREdFSwwflLFhP8aTPEBCDf8Pc00oJiCKfa1nX8+7wn1BL0fxOqa+gKlYmPIPjL5
SSc23UPsgAFAdrzyaor/0Z0jTFFsm8zY4cpygJ702yTlE4yIx7AnJxB8Jvg13gSsbTSBs5QBv02L
JvB0A+5dHyUzFd0qqPqWk6txD9zKy0dnbqZRyZyG85y92VAyHVNan7I4fXHhnw7UAuvg+3rBzdbw
5wtmTmsqcY7TyhiI8o7jc0M0MeeGyIQH4GEtH4OCaUpkCN1KyTNdD55Rhxv6I+XS2W4EqFEjpBnc
yXtT1NXW0BnnKnFaE6yq2+DTZsj/UFa/88fU2bTXQjNCznPrURnopenT0P2wOeWeh5ERSQARazKT
TbsnO3/ke4AByGm0v3dbyzT9TvLvZf78Yt04dqxSBZimSj3rzTThkT+n6Ei20AvM72uJOJ7UBqlp
j/VOM7uhnTtcfDUu5Le1MWrQpQ9+IatNd60wIJg8UkepjzwRdr0MoVcKPofqEvdqWWL2d62Jumu2
ugefZrXNX7HxhbFZl/oVT4ntIabeURHoCKz6JOXZQSTxu1JZzoN23yfrBvuJPgjFjiGA2ccCq++s
Xbbr4x0Q4D5T80TEzLycMaZ154XrhWpUnRBVSnSeo56eIFLhychbHFn0eX6OKDxhNPOyVed0dqfB
AYKn6RpTRgsCC9gaSTlhDwnIj4LVkx/X5l7Plss+BFRqC14935h2yYSAhfxuphsDqFVe1CuGTebI
rVhApjx99Kie7S8oHshPBQaIReBAkv7Wf/DCWGlZnpBR71mM7Ta1Kn+My7MH13c4e5G9gyez+hy1
QAlPUFgoiGCMIVHdZRWIihoOPjVZ++YklbrIn3IH9KAe/M4inS8I1Zqr49E+BQ3G3eiRtOpWuNId
WNngefZ+Q0bg4e9lJuOXutCM4yyNyiBWj+oYkTv0Aq69/Be2dYBMS4LMjGZU2nEcbjsj76Or+JtH
QhP7cSThAIlsUQSMs4xVajfyJJCWnII1+PPgD6+AJyMj9K/C7TdQdfedQDvez2UKyMjpZokW+QGX
uoZWLTmqRlt+Cg6nt7J98ambZQb7S4jlJuN1JNHSC9IxrtXZkswJeMAvlmz04KMiT9GMoOkFxa2X
NYgffqDXqLrvU6sRCwhyqvk+yc6RjdDFRVOb22bhcjmK+8WoheCv5jjj+5xXCHi+OXx03ppBrqT+
dZvtZ+9ah5CtivaV2vmaYwfn2BF+8kwEEmvANU5IL6gIGdyN347mO8Q/fpp7+KZ8L7com33B26JD
ysoCxihy2HYh0RZW1E46hjYfBY7FEFr1uOTi06UOnmKNHQcp1IowDlrTrMQ6n0b2BrBYepZxEbHw
oIRCbyFPm7qPMrTpw/T8BsBaI+5NO4uaQL729thY7/rl72AWLzdwQvwJpeGT+Y1K2kQYjTk8uZ1v
2u6xq30hFYFcCqpdFvVJDYlpi8qCEPeWhEdbRYmQGnfB6mOBcSEf1BsmVHtclaWaRlcHdCu7C18W
OrzAT1BMh2z4J6JNfGXX20rVgBUQhYh11xecSA69B/X+2Yt3of/PpsZ8zHH21JFgoTktUuOue9+N
PhHM2i+tvtRUrCUuYcKKAU52DLauhbNm+1TqQUQ4/pxBCdEajQb+hiB9BMNsNOOSdv3qaGrGGbnG
3DhTuYuJeIyP5YAbhUQUGAhVq+ri9CAMgsjdBvlbIGr08EVfOETZuKt3BgjvTu5KGU7eYZzSYKbS
73Ie9xmfOd37TkLsj6M9yzPhYZ++8blqqGZDcLEIDPaHyh3vp3YUMrvCsV1fxHlmkWPg8h8CrfTz
pQgLuaeNLMTY0DC0kZ5f1ViMbajsB9TPLd+sFmRuVPf70ZlJgS3OU96EhVMAni/cgx53DiorFNHP
1YX+72SNcqAyq8nMZILaTkUS9D31huATde0/7JRCPyxKQp5Y99IpToY5hSOilCk3lkTp7SlM8UNJ
Ak18zrB7aoMmsHdylUzhV/KDXOgmm4T43kzoVr25YMoHYCXepKH4WivZqPT6nhXkp66WiW5XQxFJ
kBfTw6YMqi+ZSv+5+9qLkkeZCUlIKNcPDFBZW9UQTTMfF5RD46L6jGxsLM8klFuvTzjCZCSQXxPr
X9VaxToK/bjHAkIJi2d6RVNhUgKAu7VFfucxKuCoRzs8jCRKdS6+BxfI5DD6OPqCI5VMtqusAyUG
wTselEizI+IYlVlc+NV96sxizcbK6BOhj/O03PeXsBcNhKJE8xYwpy9VrcSaRWOEvSsPcbpF8Rjv
HCV9AP5CJRf9GCFyJw7f+Xkuq1ABzU/aKIewikGxZ5zEg8BxSWP860p0Ks+vWCdohcNW1K0OplLa
FziJD+iofNmmVHPFjRbn12/pGnimt3cYh3MjYOw6LiStUHX26rbA4f/BecFKLRsNSZ1qakdEsj6z
GfRd09aV53cYU+ogs0m5jClPN36cJvv/3jdw+6MjemnjYN97ezEP774bXgJScjlcOWefC7dbnQ7l
HMZg9M+XNkbw/lWGHoMaPSpcyLe1IyBqrHSkRuanx/xGI4wq8yflPHSEmLaRSsx3XJopVRDUpT+d
M126ghmiLCSagXEAMuL1svBXglRWnC6rT9Yn3X2uadlH9T1L1S89959RHwdQ947281taoNSc5oV9
vyht+ReLYvTxQbray7e2zqSnL9lF0wbeCvKazAMAqL/l6CNuBvI1g6GuQQO28WrIrru0ySH7eadM
dBI8XBtrF8WlHVPXNdZJBP6pIXwvTK7jfttLetF5t1DYj3Ac/gbp/jMSmt2PCcc0PTR626AWS/EW
2Q5ipkBchhfIlxvw1AZcowZKNnMpiaOcqmXwbSzal6LOcchjG5/jQlHef3T8LZ7PTsPUgjV1uLeJ
7tfXGB2wh8uIr0gaplF81/W4urvj6cTXDaaq3c07pC9st+e7Ih5NyGsSBpena4ja6GQpTvjE6/6P
EAP8PF0UHW7SeifD2DFw/30XPfbSAfAmV69ElnProDRAzEKqPEmXxPCB7x1aALc9inVuLuOqYI/U
V9qem80+EvOrIn2cRwRv0zmhkvqgPM4jRlBqvTceT6zQfeFM8NJSYvGXE21cU78x108YaRrP6zEN
2qY65quH3fw3AU6Jyo12omnHMSLh7yVxzxJXy7N62Jd7GS/DGCGVFxl0Ar+amJIMQyET8jJQsKpz
O4TV/Eey92EBZ1jp+dI7w1vWYhHDDusNVHtvIl4CZDDpsJz8j3DXIr6qClbnDNbCIx3oq5KEkpnt
fz21Fjq0lH57lNpkGkJHaTC45E6ojHddauO5W3rxpaqoe1RnahjH+UMot3lWiHzckfIwICBiYNRx
+oQf4G5eG+iAuW/t3xppycsTjUZmsmo3EJFm/ClGsuK8LU9UWYxCuuvrUD9rBVvA6tPPjA7yHmGi
b7Fb/EEYlth268ApfiSFQ4sTnMhCnkcabX7RQxPeN+jFAArowW4q4rpgFnMN/hGOdJq0Il0ZCicP
Gyl3k0H+QH+70JVeWEqbDeAVV4aQdXejf2E6I66A9w580/OM5iODV1dZSnRDthAk1V0wIkjRU0fU
CbDLK2LrXRdxLS+ft9iFpT7tjGC452pp8NLUVIK68sRnsUQXO5G6mkkuX4t8WlEnXbPvFR8AQd2v
GknKs4G1LuPrhHeH9TEOLGlq0LVSbuzVYeEcl+rydKYWy+J3aES0+8g+vOCCR4to3TSE6z2e7I3X
1cQpLL75bspiP4XoXMg3mBb2/5RKJkvGUhyx3ex2RszZX+0n+76cW5RTC6lEq7UPLBqZJ4G/yp9Z
crex4rLbFyBfqIWiM3+6NyhoGBx0yG4AStfunePSW0zdfaHRi9NPZbnJ9MORuGhhirx1a7GCD82k
QrkbHTSOl1DmI2Rn6UPRWKizMsOjCOJia/cNNNtDBH5jwru/uxMgkUY+vdYOrILKODuQw+GydvXk
BwZ021tf5lg5+TIFBREaCKDmfvvx3hnyaZg2O4+WcE2oa8dbcIKF84sTTWD8I4SMs6CI0bqBaSWo
47kScpHmSb9uNLf0vtFuYGtmPKfi0pWXzgWeVieoXdwVVu6Q/jvmAXXcBSKj0pnfWVWm+P/fZnBN
kb/d3zEKsxNovJO7lIxJZJUvZ3/Fx+ck22wFFRWIqFGL0a/xOTWVXlmtkRo26GW7sSG9xFw4kEK7
iZ8869eMiahZIO7f+4hYgX+urwzCUv6bJP3L4ITcVlD3zv+OhTRdZ0lszNYjPoEVARN+XqlxDjYx
PEJwvjUC/JrnvXaVj3shiWPynN2MCefiCMhLR9Cd2yQq2AUHzvHvNqbf/DdHIl9j9YTVa0yKG5QP
K7U+IkGEpNrU/bEdiCFaaHaz3gioPeGIMoEYy94CXD+GEKbO/R1LlHGROlQ8ce8xroU2eAS96jkD
7wv3y14t5q8BV0iEOODLRjYb6adIK1ZIR8ngiEwQcrgZ8JZcP8vwaTV4lpX00+Ro/gbSSVlZSTAA
w8U8qs+dUD4bCjdyIxxJddfKma3MHqjn2fYpPz9TKOk5IR8XQOYjZOLRchWx2SVzm1mbs21vC1zr
Bjivw3uuBd3ujjK1aNr/eSJJKplJHMS2TECS6LJR4MEv8W9+HAOvsz1Yx+6HmpgEO4yIaSfAHPsG
C0ppOA3+Y7XY10cGC9syqrhm15Ce1sfdIkLps3CbSjJ3Rer+Opn39uodjMbdQnmH6bQClQXjwRlQ
0A8HbueXHnLvWlwVodRZ0M+EqINsz7Eou4O1WNPZ4w+EVlK5YDvwFpM381vSGjq7YnZ+PZLO1tL2
Ul0DynPq+WKrYxF4EAYsp5NCoKsM4a7XBTUpo5hmkxi3UOdbwQKpXLMHq/rZCd7vlPh4o3hL716T
jGagIovGIW0HZUZOB0VxpIiorF5y98JxEeFs2AEN2t29TvkDSc46GagfV/3yAtA/YCTPILakbUSs
Hlevx6LCfIPFrwNwh+3B5V0a65q0JQQDrXPW7qPKX1ndG6lQzkp1XNIVWVQBYFRXCBLOOAmJjD1q
kHjgQ0i3MpYUS79U6g3swMn8k5OLUyFjOmHWMadgoT2Y/PHOSwyL1trKCrFlIKbC9pl1xGXP6oIt
Mc08yEexJt6kkxasgVXpbcyDG4rQPUC5PV0a1uzZ9WtpmxM7FAguElrLElUBeAcSq4hyfPEeVQqu
Xksjzx4ozQrvm4Z6pAy+8Axxh1hjJecqhA7tRz07xd3oFcAK0mMny4Wc9TaLMDI32No7wzWVri92
zTYOcp4+zbGBj5/wKy6xPNyggfoMRmISw0iLcA6RLqrw3f6S0TLRQ6IV7qYGZq5wITJxw5KJYbHi
9KjqzGJvK74SNpdEnd1sHmxOC741StoOqCkTSl48TpPUMcperPthrxddcxsWf57Iy7Yh6THrKQen
gp+gmYXRw6cBBce7c151mYar36wQ7IvpoNKyQhFVy94YL0Yjx9PqTSCr5WERXmgHPX1dAfAzAhdm
Z8ScVCsh/LGWsHWRfo1PGYb+MjwfeeQE47T4cdS9gTdVh1Zitj+HnyaOoW+iZn4mBMsRxIwnxuE6
aXaTdi7nd26xETD1p5c505DTYAqsbCRQBxKfCkDuv5dBq4hsI5rAu1iu0Yrh0rzLMNcRpOQtp/fr
mmpUyA4W3tnUMTh15WK2hDZnYfZyLs3R40rP6scnN/bZQCBHc1fTXNhyu8FoB9CBgIwidTKVtY8X
64GEWHeQIrY8YnLjDOkne8wjl5FzLOXxlpo8XQLXFeKKaUfdZWWxavx8FNExZDvTbI0OI+QThmeQ
DhWuP/7woSGdhm0/3oHoDdqx6tqDcEKofFA2ZAuCnOiYc67d8yuGSA/UzfkQTNIuItBXqtxShYzA
4z/LuJpdWF9IEKe9ByunWmcQbDrDNF0tvJZzu2R/3NyNtx24+Q/edg/AvBsujeyqzGAA7oza1oWD
VNDNK7U6lJ+M6YYDbbrjmNw8HeNCphlmiaZsme+xJpK9ZNdqaBw5N6EoOk+hLaIjgMOKcHCQhJi4
VpjTEr+i19zXGUr3RLd+M4yJn53SlCoH9EYVPW+SknmwqAqoe0Xz/fIm/NGuRIE3KTKIq5cTHqYz
lKrMqDJ0RSZiAU/L5mwWZSea/gsCBgLSn3qNIWagjc0QdBg1W9WccCrRjIKXAPYfY7dlyNowo7r2
D6VPPZq5rSWa1BWCD7GFF/WADu2iqXuid/HvhAzt9OOuhwuxBOBVsevZOc26yZUN0olimfO4lsbC
PcCeNJfRk8z73OOdsdG3gMgfqnxEfvm4N5LOqdcOsZkq0wVBznvPVJKZfF2ShjdoRobp5JqUIs8n
xYcyUj6BWnutUj9wYgIcbUjDsHONfnHTZAHqKtk/vNHuK6VbhJbF3KpYpQv9CaC3zC71WT1+Rn1R
XlHYDT5wSgn8rzHWNcSj4EXMldTd9zd1gaIRcbOe3V7lEnzyanJxHwzGMILLRwO07+Gz+FuRYgzd
El2fvPXSBerjTuONXyLnvvr4XKvBtolCzdLyuioM+nToeXIcxUmOrgfTKkCN+lkVPNlFrlyxFhYD
vJ061IHeKGoJk7KNjVAlsfDlxV9NfjM5WOHoCtBPohFM8e7A9D3E0h2SFIJiq5NafGhGDbQHlzPe
J8fGEdFv1tSb61zpE58smC1jb50z5H7NrKcaveyFRpmulCNbzhuy8m18Nw4Ngmkdbl87Q9mJxWxu
03gDv+2CAKOsyp5cCBTjGF90Qku84CUOsEhIdYQEkqJo0MzSjpJItS65o8V2a614mDbt+2BaJG38
JGzJ4So0Rh3FjwMDcyHzJPerK9YWreVY13D0GWbfSYgQFOk898yC7x86HBuBZzpH/8vEgvfGLDbS
HH7HfPeS0iMgjP7Jdc955vLdcoxmjkdjimDQQ94Yo9AAcagb29kDWVBIahVXD7K7Ge2QAXSHx0i7
ZrU2UUnRnPlr7lxs/AB8MzaJmpw9VubhX0hHehG2HQ2+PoLJZJgvp2Z9v8DiM6fOd19BS5R/j0W3
zWpK3hDQYaI2/kPoA8rrvwCWe6Q2KOMRszx2B/HrJE6Dcv64hBULDmgnZ2qjvs70zBoZ/R3zKeWF
kColVPdJeaeUUTqAgFksf+N7G7PQ5w0QHLu4rzRxW9Ht0vtUlAOcswJorYcb6/34i+4HQQeCrAvr
OEHqfslOFj9wOPyj7/klNF3CboT0+o4AkBOmUHHhNQv6v1rZx9+5YzfD5PPXhapmDRT/JtdnQ2Sm
jVhBCpk6MQ0znIccdmhLGhVmhbwyktUbH+BeiJc6N0uQjxaJ66YmttQpW/Z+j56RkIzED1OXKB56
pypFAOZdMQEtxVApmP1ZtF02mgiXP+ArlYzRjTvOyj39QgpxhP/Jcv9RQsliPR30qEFK+FTgPG5d
gRvOGdnV5UpYKxgTMO2llBuhyo7FjVKkXQ3JLWnmyB6aLjI7GCWdUIyCaxk3EjBPVsQgvh/qiwfh
5SPjNUitEiw4lSi6STIp9ErjcOVMJn2t2RKbPm+FkTsCPB3Ns8o4IjiGyxgHQnC4uZtXtpZjbORJ
Dm5RrbHqgsc/YWYeUbRHVpO+yZ+8HPeiz0jYQPShVPD9YormqCU1qs0YtsJKS1RiZYZkYB8i3gV7
wkMlO/MYKcmksFar6q5LHq6qQGmsaR4WLe8ngd78mUJG7NdEKHgr64YDs/pdvV6I10N+v1UcofkE
bo6DCdm9LKCifhvR/moV8/AdxEvWYrAWFGKWwEjplnZ2fR4A4EWJ07KKIca7Tps9h1jqyMAdw7Zk
QJtsYTpE4MLeWfcSFc1EArQfDHE6SPDLpHoX8YkhlQPwmQ/CygJNIABbHBFg0iQs/2kOXvOoe1eJ
QbrzyUVtbJUv082tfy2Y6MRtsulf3n+1RD1mzxJ3aY5PnSX/ZSAhOQEppr7rWtWz7Noa+/Dmlwx4
qKa2tIAytVaFRcfQJ3vdBR4rRpSqfuUl3vucgX7r68p3a8D7tEcI/HjWs85xsKxLR4J2CQHOWt2S
PKQo97IWeLhPjT1g4aaHGst+05yTdVypFLp1k7oZACbRif216/ZIvBj+cDoqLQP2Y7ZD4vweyEMQ
kCS3WiUflB1t7WFB+P0d57MlEQoI95shQYeKJFMxP+zRqAMIwjMQWLUyLVtPK0jYj2QyfJ2GtbzN
9RgHImjW/s009m83RzOzbaeCzfiJEzsq0CscbrygWADqfQNQAMyDKz/BpZE+LK3vTrgpOFmc4Jen
JyZobnDm/nhAplRBsl1dvwXPB4tM66qngNmWpcbtmglzAMOIqVd7Ao/+TuwggKysZDaMlvmLrsrN
vgFT75WI258N9d7SZfhIcLl7AF/z4r5hYlFGCQq8DSV7Q8FcMsGBvgddZdLthokdk+Sp6E+v7jVb
GBlIhHA0O5V2/ZVV32izMpJ2rbkHKjUvNqBHKg1mAdqL04N/QOVzDobhrOlgCvNGImxXtHL+WZqA
9dLBcelrOTHdk3uZnM4W4OKyC/4EWn/A7NrsEcuIFYqGLqUA/TJotxuQErYGngdrrbLXYRk5pekL
JNXWtS5+ivhsjCBmfUBC9lJ6T3m8cxu/Y5XezAk/Ecr+EE6l9P+bkrLeLUKgiTc0REkokvd71dMa
Woe2NOxK0wOyNkPAogPvRmhTOacNYj1RbZ9N3/fpVlN1BYPOWQSVaX/ydVapz/ZOodQZlmXP8Gx4
t6vZkAj1Uzm0/Ucyg+HD1VnIluQwBI0jlicWxx19kIcWImo/d1NugT3T0ho5DOTQBrDnU4AanqtU
WhlSqZGPnbF565jHQkqUjWf7VoOxGlblHs3m1WoqOZgbVhhz1tTze1EkEtifva0jpvJBpv3J6y1i
j3RRRNvRiPNbj3Ab/fNQQN6JjfZ5gExFt06ScoExA2bL3RrclNywg1w4r9VTlYXO5HoygeYu9Nsa
UjpSs5LlsuR3hApswTfgDrGy/9j70J953iUAg4FtblR1Oxdlns7JOzl9k9cyjjrMEP0yqAsHGK34
FqP05Uja0SbQbWxJZA6BZpUZPH04C9hYyBMnrvipEQtxEQV2ntfjCJXJZSXNnPMnDvwD/iLiNZoR
IpJqWIBAqVBATzsetcyjHRHSK1I8jwCrAgFwBxvwA+lZYziWAt7hHDUA9oN0sXs9mZwsuyiClwPx
NEFdAPjdWk58hCpXGJL/RsiDB5hM0r6O1a179WPFkvBvdvoBwSIDOlmI2jSJXhSQa5pCKeAD3Apc
BIZlYR9zqpW8JZaQg2O2wQpAkFbx/MiGTpDt6TZLVPXItEr4BdGOyFcdSMerB/6Hd1f6HiHN/GUv
J8Yg/JqyRbI48V9hUwkGbZkWpJfFgCFZZWziBX1nEH81a+2HkFoZHFje7g7mq10NUP6x05kqUKDz
1DFyfaF9Zob2iaYt6o1D2+gUSSJ6uMdO9CKGByf8IjIlE7QaN6y+6wuM9+TaIlmSuTvOqASuD9X6
Gkjw8ymbDwkgSvsLIBb8AMVJ/ogrRCuzc1VaV91qOkSP/UPXTFenW0t2OmPWIT8wKHLMpEDRB8Bo
yPxd1q8g7rKygUH1uCRDci2HvElkWcmx/PFcZUU7KQvSOZt2iB0PT1Wh1Or8Ienk8OOfQwghjCWl
spue2uIthcRezUcnzHi+/t4hldrjoQH7N4jR9CTR4owGjC6/CNtIZ8XpHQj70/mV4pUd3xe9fEPR
6qPekS8JNvHMDGQMauQfQuhFpaniuzBZ22M7js4jci4+WnaUBefTqsPvdhHW+Sx5aeMCsbrR0+0t
dDXiloddzEOT3DYwXBYHrzoOem2VgGf3wEpcGVMUwTkw+EBT7mny8o9oau0ifhUJeAVxR96J4YfF
8vEz0m1CzmN1BO/GTN+6hZ+kBSGUU7fNkMuRENR6PuofJ5uCJuwCVk/Q1WF0sR/E9iolkPJNiopP
4qXS+opE+PTwq/RmXFsK1adnEPRncpYtJ1c5Gkgw3FyE5EQpnwsx7W2FJsFfl9zAvIwGaBbYBQRj
vL095juRcIDDORUtEip5JDB5TvjvYdPnvJEj/p/fq1uEZNS0H8aqkH6X1C+696LjRrQo6vGzABPt
MuszMPt4laV15eqBeYDSpV0Np25e4B3AiKdcgPYOEliOjnMBbPTgcUn8BAYzWWHvAAZqKe7yrWcb
CZoanFKRsCrTxsxSKtXzxhUUCdRztCmx5GiwqAwyZrTQfyUnGNUWNkxUauy/v2Fmf3tas95lvZVN
1FEdtU5lk9vB5Tzxb2pnuDck6tdGxmtRnI9pnA+3DvDt91kF9OcWneVa0QutKjxZJrwcmuFbCGyU
kPoHyQvr5T7+CbD/lkbkSGZlK6YHeWc9wApUJIHauOGk0z7Hu2aW7sg0sOvO8j/C05Woo7TMRSps
/bvLFFhiMvj1WkWObSCG9c5CNTBOQo0KKz5jFgaWKbO/jSHvggY233IOH3L+HMB+9hKXXS7TVxQW
sslyZLM/cuGSkz1vcQjhLxSurt1n7YP8u7Q00RaHcMvrPZsKKNEa+QFr6fWBpCYfic/aXjraYGp8
78+axVVpZUKtVpldnm3pGXq44TUA99CMbPJ0oY4A/Jl+8gygvDTslTqAF/9X4SIpetbwhxDoqcNJ
IiKhkxHJHnZlFPnPQzgud06jjx2w87dv3/BObscKfc37FOVoOHXw08mU99yjrKxAKq8LIzcbwoxC
PhST0qoaA6GKHe9HvXbKWdNPGwChxfOx2xCuFn1fyJkZ1ECeMy+quadXeQKQb3yaxRvq2rmOJUXq
4HseJNNci3HGSr/79AoxyWkhbaX8MAOCWnZzg0aP0Cm9SxqKKS1ALIU1FMVlCjzX3sLtpUmFGFJA
AUBNS/66taRWXP9FiwDg66Tk0C+ms3N9Atzf8OfFhxg+xnY3OeVE1gelro6w2C3/YXxRA17UCt7G
xsH0QzmcQYrUjbwqPRlK1TnsTmWzkXsZ07cqSllwTA1fGUePcPZTGByd23vTBxY959OYjYzrwB3Z
A9127DjL3gW+E0O5Hp7/T+DH8CxUiBK2iesBtUgTt20kj79aNdejWYhlGLhUZWTPSNLq6iqTXteY
wirHziS/IgGtWHlyMPly98CxTW/z2/aUiAfIGycsMYBX6BKXr4nTMR0eu7kCm40ZN3A9WBwQ/eVZ
bYmmmqmEcP5rGen0dhXMsGGYxCe5eHFE0Av+8qgNrOKMT/9V7uPwbK2FPZ24wY7EGNCT2OMRUylL
5/uc8eFjzf8qQXoIuzNtg57SGzVYsEkP76c5giM/UT2xyFvvK7qozPNpPQ7vS2wPy9hi9k9DZrTx
WFofgYbT5AmAiodeqOcijWmi/2aulwIHiPX07t3ADSJVLnH0q5niT0gZF96ytxcFiGsoj8VDZ/so
y8TV0vLHRvtR+oLFQfChQy1OsvGk0iMCdZE2PZn4tEWoJjyLeYqb76c/67bXxNdT5/Vz+rrYdb6p
Q11iAMbmZoxHwtMt/MdPrp+7zRKM7sII+lJEpljDcfXOoNv0dvxFqbgk5xnGyH7RDM0KTKdUKXm4
W3pV0riZqn+VY2KhrdGzOv/haXn21ylWmh8/2IP/FrJG74BuLwA11gmwqVBBIp7KGcibSXWqIZue
g4mRJpiqOasBLmpnPUdh4OkuKrgaMU1IogCyvtculbYHrv601SzYrDYeg/0OOCs61PdJOFOIecOH
bf+dgLDViMSRR8U2mMlL7feEY117EHbXX4atn396vQt7Ogg+0d/Ig9tu0E19gtXxMYLwce6mMtCZ
RfJ6QsaBwhgAi25wy7I8zEgYbZND/oaGCbChbd9+cf4fcLoV1Zfe16ej3Ua6XvFVHV9I50JvdGkX
7z74R8hUsJhusomzvvIiD3EjyfsPbGiIgZ5AXjAlz1818DIyyw14rKXNjIhXP0q/YeMoz4abhFka
tUzRlPDaLdbpqydbP7Aigpu0PfZ6Oh+56uswypcKeFY9clluvdrhy2FrFS2SpOtnIGbOW+itWPmd
8GFiJovTD9GdbjHWUNFChtAEoZygXD6zNKyEhtsyLtdqGHNmxSPtgHozeGFpmLGYjAtVPR8X3YLX
9nefV31PRnnGDlU+ZOl7XTfi/jZsRncn6uV3jLh+E8A+IVynwZzxP6Irnz9IGjw0N2fWttUopLVV
qe9zOw7ltJWkVhhPTkNtsFRQKaQ5lnGHTKLMBptC02FcRENYtgzLzl1Jx5KrSJgk5O/AvF+Mly08
fw7r2Po7ET+r2GDwlWfhTRsW2Psce8cI675Mc5krj/TQP6WzdY/82aaTf7a4nvHOh1vtx0+6o5lD
JmIlAUvB4c/Eb4Gvl9vth93ANtJUbgDoCvqcf1zTqawBtg/juNl0NeV3lSMLb3UOTPRx1x/pBqVz
f346U9O2OaG8i6Uzl0C/rvPgGHKlT/z0UWo7t5ydCt7svbWCIb5WceHZLjVFnhHGpCQadehmJWOi
vB3b3jx8QPTivLdsDmmajyPTv9N79YU3fW7r9Zw+hDyv/DvgqgSeK8ajEerwB8kWvZlknvY+zWR1
g2TR4GL0VjO9MMQ3anXljfUzs/jNHAmZt1u3BYHYRzyaRU2ssbqK7FfTe8UPQPC0RDV++Ie7eGn8
B9fam5gORXSkPCxixgkq+BCYT+cPtEOCfHGV1AYxmapTi6Aim8/g9OElGOtt7gIS6vxAAjMs9Wzv
YsAxO+gX0/8GkLAH07m25jUnwIesRw3lzRO+o7COSjCighz0yHokrVGW7W6hOMUj8n6vjIAKgF97
VPfYWwjvvmqXLi8QseSRj1GNWwfrN1o0+ysvR9l8ljIESrZOgy3hZtNS8fWPWPUKeGyAAgBdaJMg
0WGsw6E41eE9gu/SAXL+hs92/c6LbjA+Y9L8VMZ0KGns6Qfoh8ATfTm2V0N9Fn5WPzkBwVeI9+2k
cm/TSGC/op5hiskR7E5DbzqrFIXCGEnkkD7zENf3pQyI0B29uLc5phNUv8CFigXEYLqfCLS9Egdb
s0vRXFIaO+1mJLi8hvyveY41OUFXZMiF4m6U2XOjDSzm3Hi0Fka5gbyFaTKauPfcK3FI6+JF0dTM
Pi1lYLc2+uuEPAAZ+xLWuKpQEpiF+SJcsKYOklNR4uyL3QAEfQIJTwYHZ0BM/m3zU/6jhA9SJCD4
oMrsFw0Oc1t5Mjl6KHfZpomF6Y0Z6mDVE9l2TLvq8jv5+AJYxtfYU5j2OvZRtsL21yY2dL1rx0J0
HQPzQxXLpn2hCimhBj8O2rEAxh3r1nBO+AwWgVxDPetweEY3M30D0gSJgqfetJKoUUIUdskngKjd
dVT/Vw7fvgprlDoUsyMfhMF490xnxpDEeGIDtGax9fz8BNc7ETZmZx+GO4Tyf9OlnKwYDpZZLeLx
VmzB1odsyP07EVlfRcbLfrQRUEzrjvN41gXJxWGnCsKiCnnF5Jd8Gyv7AfmXlsxVAf9j0PrA7Law
RrfBPmcXD+UP3/GqMyfRDLz5MpzyhiFQ44I8EEIK5/9kFDXYjE+Yd/xxDW+hecrLVVFJTkAHNCOm
oPbRV9kbk3XlRTu32XnqGtCYrT8X+HDgs5Bo7SoRkyHOScRCN5xaB15XzIi/vmZYUMFt6oIzwiUl
LHtYN3T3KhTRZEXgnD+BksjQTV02wyRkjh7Og/f6+lFF8FD6cPn4lQQovRs9ZELkr/NIQXiFIJaY
CtOnLHURBn6LhugYaXISac+ls4bTcBhXJsaTZRaQfe6tM9WTmJEt7NvJBD+EgQk61/4knOGOECRZ
RNSlZsFpR+vNDApdfrRHDHVzwjNnmmRhnHao2Z8Qi/nQ607O++BXG9hWifJBlBJGsbRCM+ET8z0N
UFr49c4chcuJIgjC6QEqD6uK5zVQ1m0EVAao6qFTTI7FonkdPPd9EloNQv+Vz2v9hUp9Xta+iBtG
+jjEt0JDANR+7FXTRUBuyOzQ74BSehMPWlft/5Egeb0j+aDRueJ/0xaZr2JmfUppiV7tPK/W+ETD
zSikwJPSBYts8WuawRYjqbz7gq112KNGUXmBqBZofNOfQmdZ1O0ny2RYijUDR2PdGiFyua4ci3k/
iEuPGJjcFnI+myfS/FN/axyH/spT9NbVwj7z316In/pNWvT5FulHPO7ALz2kDyoqJ3aUYXK4EO7M
HCDcICLwWkkdeap1ch2YT8gM7Dy4Glc6q9pv3nxTqHF8jArB9K1u8CZwLJQ7cgUuVEF+r4Zy753N
yJXsViQJ4DL/z8xQKlYtKib34kjauIuIPvWJpXNs3GtxzxYEYT9YWUstjJRvtA9DK/QgMqXJUYlb
llpq5f79xQtYeWRYc+e0UbLa/j+UwRTxh3ZjpVF4fcTbanKFd1cXUHQe/j0RcnF4FMe6sc4aQoyz
817Gzeqz+UK9W0DhNqHcUMCGFpXsc7pIEGQVRIBJo3KvGMAnKFN45/6bc33VH2zPdFEFemdML6Cx
1xE1FB6kWlGV2JwDAzcQfaF+nDSc/Vgjbr7a/FR61jOBePZ62wWq9gH6xnFXTRkY8pOOQgmz2SSI
/EOQQQ/Xrf8AEtxzLRq38wf5NGtraSGDz32/ZefokZau25jwRb6KrEhSTiHEkGxghJ5xHssxCobc
W3UTPoDsQ/NbnSJoOJaW0yUdbx/je9zHVrdesSrZuj+ryR72QdzXfH+vpecmugIn/H/wphKmZ1G5
8qxJ+e1uBUg6UxamSTFEhY07P/sn6BC4bW3nIvbnKSOJmVZO47vTZ3yL94iMQbv87yt0h18KkS24
hwzkSLPwESYH5oW/Uvviil4Z0pkSuOu1+L7ToNBeV33JvOHSKOTVVks8Y5kuDQ3zSbMbZxBoq+LC
z9sa8CwrMevCsn5b8+H81YvW82vL6I5jnEJVszR/BaWqZGEKARef4ipTy64N31eIWw3z3vqTZMjM
YIso525VJTjojLIo3cna/7oi5S+THMbH3yt5WpDlvuC+iH9Cf3NhbzcW3RCyT3pGsQPskV3aZ42K
B2hxFfPi/XVoZGYxH9UIFyZa3YC7CSj40m8KyKOSE3tbxPKOisx3IsWDqePzdISj7fcQWw7v8Ne1
HMnx3J+DO9keASDp1i9uKHVvofNv8MrbcVuuRkJwd49pTLwWyQfwuAzPVRECcG+Yz5Pb2gU5A+JB
AIWXWwCXd6tJpdxtOC0VXAQrlfVcWkfNspBX2i5nMt2K8q7y1I+LfTjrVynDXA3eEa/l8n9NL2Hi
OjiGkBL56N85yCBzQIv+9ywvNE9SPHwhYzWVvYb/4PTPa5uX6K42Ew2CX9EPHLLYUibAXVg7REoS
yprrk5iBGRiZhBfaQ/yvZ9m+gbx6BP42SaK+q3qFpkKskGuEgR7SvEgHKfpC2SRMy9hpVEfnTn7G
zI2GQlCXgyT1fzTtZ7FxQF+Bc8fYIfUKsatnYUPjcVRMKfd36r7PBdVqQfLMrYWss7IRoyhy0cX6
DopFylogfDDeyyLpcZOpycp9Z+pnfUF1xz/vpfjiLmlD4tBv/3Yqii24McfUoiZ8OP8OysUwV3SP
sBfqokG1Dfn1lOSle/hjNIN2BKcm7yvxcThxenzY+UfxUTzydW/D1wfKzQ+82KQhdj9xUe+6XEpD
KAJVVvFP5+q39gwXNpgfi8QVYyHKRygoQQjcx7FZEIJ6CLijPbHpUhlI80sCCPPqDxm+PXN1xMQy
vLVdfN+7lsqG+a9LyYcAN2fWC1gWfsMHew6w5ywmXRGPXhLfSLCHDJV/SIz9OOk2gBLWxPEfAXtK
2ZOciJPvIu065/MC3HfoPsw33GsUdJzzE/sb8mE2O58+Il/eHl7iOB2D1EG7Mx9sLQ0iEMqP8UYH
EbbmFkNG60P5JlJ5PcApmjzKEEi69bJIrTG7mxt7h20WQDed0QVycRuTIdjskrPQ2jz3DVxHxi3q
XzCQg2grWpEWCZWlatjkXWIWAmOApBc7uUt4HLyNAFd8wNYrwSdmvC4FzkDwwlqwx7kqU90W5xmR
zBLJ035BqvUHUj7wmHcs2oU2jsqJ8Cy8rgxBQWAO1tf9+BiVYTcyLdPhqkE/em1Y9FKszPR/5I1Y
QkUyC6+HlbK26HStXzp0HGdx2pSgPkJRIjgAJlIuJZDWVTf0NMMKL0F3PnW218+lW6Mj8yVGeFEk
76M+17Pt95VcUKYd0jjjRepqvpwnhqsXoHE2fONtZO7XEe9DPxXyrJOr9MzFAmZfSpmQTbDsOgvJ
rQLob6batJrDg58DEKMDt1ps2A4upaH6w5tHMn9EF2HxSFgwIe5MlQIX41YPLdURWlE4AG43QjGH
qEESkLOoTZjG5Sy78VhCZA5c9QX6G22R5V0weTGKZQkxo31FrkEwCDegS4dsY0cJ9O/xcwa2m8c3
SzsK1TGkMojMlkXUJNK78Nr4y58EuuEFADObJ34D9Jy/EZxPn07BBcG7mslR9uaQ57Js3pbWzsiD
oKbi7eUxJgsZ89KfagYQeJ3H8Hi+Hec6cfCpVJDFDOQhPFngmpj6SKHMz6bP8K12DcLbB9Ap5wOk
UecG9ozNAU5h6+os2cOibFU+9lId+qnzQUPAWEsRMSAdjzMVSSPEFgfeffD6m6xVt/+bZFv0+Gvo
5xZCsCk/JzGEUO6ejYmCO5x0calnEY+Jxje2nuf43tD8hEipXhOH8wp6Q2UWfrk9ECVX0Sj70PIw
uVQYxRTrprsIOUP1Iuz4tqwVYbLDAVemf6cm+6PAIyc+sZeKeo14VbiZVfQjk+YvKl3XBtwjFNCI
c7aVv103d47GtKmvcGnuuBCYAA35L62ns5BNd7xo08F9yB5ujlnWm46EONJRmqsJGTgGJaq5O/PI
e6cxuJ+5ux+ck7mKjr325aOv5NnLrWfbDb4EPQY5FZiU8vmY0Z1Z6ah1M2CSDzsYilSmj8woGjie
9Ekob6Bb9ssbjNqZFuqYogvCSVH2dy2B8grmCn+VDXA7ZtZUH6RfpYPv+y9GXYViv/8jqnaniqVf
NqYRg1zKSacYI1TrMkIggRGZT2PZjF/OKRolcShIht5Z/Ih1+KkbNcSvchSUir1PTsjuDL2X0GVS
pGL+0r2uwzHeS3Yrybp6FMw11D4i+wneXTPeTGJuMAFPPSJCop4kMNf3/XOyX+45812WhKYLghDJ
vcNJUSFI6ByvaQc/BBkl0mW6r6gx16YXIDBTavGnuNqQN6qgs8iBuAEIzgoLxEbjLUVjBirH2lpj
6vvM3Ckk52tuwkw0NvwjHHGJAb6snmgQPdpXJAMLFnQyMR08MaoJdG5JnbwTp8DbuVc4z/Zlp5Fh
qYbW9UM+SxdTN8dV9/dwJ8r8M1Ow4YHsfXPefYaRlzSgZgE9cbdfON0iwrVMpwpQFD4qAGDDe7R5
0RFtUCncWerlaFn4fGd1suW4DysPpHedQScZmm6v2h+fM7sAsSd2x46/1trF2ncik3fr1jod+ikm
ibBFY6fylWxnqwKjR/J3JPLYDgMuLzZFcPsJ5M9Rk9Q3KDWbevnggt6GpXu+oj4rQkqzTGcRnVwu
TCbmX9EWanTej9E64VzV4C+eqnIDvSOTV+8Xxm9ThQMIPtuwHPTv6xMG23ket2IQjN2f6E8hvjVV
u+tQvZaAYeprUyVmfKXYYrHGZkQa3Cvzx23tv1mIQjRXLt4gL8IHViCkEY70jRuaSz1+nLDbWf77
5NfIf0Zt7ID+4IuUk2szy1gQ2g7c8LS6OqL+RN2BZK4v/XcY0BDPQBD7aJv8V+6GD9PgTLb71NxU
ppmoVpRt0IdIHYlnA8CDNXBvaKs9CL4G/yMCjbujGNoQ5mFXKQ+s3U302ym/2j0yv0pxXxA1A8NY
/kduUMx+smcTzQ9qgBoFytFFbMcUOPSiOMnURw7xbVnrRE+pQ4t4HIUdiiwz+uYCCwrxbMMphD6A
pDXYtgNnGR8sFuTQ+oIRw3NWBDukUlOerQLvXhKc3ZqYmozwSVaLmNrMfnA2IScEusVUZLEhiche
jmz2dDxBvl0lkEeDIC0k3mxlCBGw+xHzm06rCwDiXhHwtd6rw8Z0zUyZqDNull9fiDGa7IC7tghR
DpWz4UgAP3QvS4BzOzKGDpjPhyh1AJlYzlpimxdgQVsjdvZUw+NhjM7qvCa5pDpyVXWhIx4LuToF
fhYu1ilKB1uyP9Yjem7H6+mMYzsY6uNR6FDvAQ8DUw60jMDZ9OGd061d3UccAfxB3ihrODsdRu92
n/PrOZJKNHLH+Z3/5Ugk5PEyMAGe6eMbAtXclJb5vwNyppJTH29xhVVZkiLvBSPrBtCZHdV7l/t0
o8582j8pU5vXPnDiGpRkgfrqP1xK21w1X2I+DXmKTewxW3AH2alLH5eF0tAyb5FycmiQKDYNDq2Q
YoeC6lsdSTfnQqA9F5CU5NHKSU9E/E2i2QZDrJrgfnLOTxNGkFpVZbLgkkBhFTAGaey2jwZflZfj
NrPSB9WX77siuGJikZU9wAoHr3EflsV7qj3yCu5qZ1510SSbguf/p3skH58VXOvkcX2YtF6r/pXM
dw6hx54abOdHtAEVFTaGDPHfy7PUJEa0GFKDvDUu4w2kUBnjcgtEnz/ssJPoSVM2fuj76UZ3ZMgT
Rp9Y2RPIEd2RiapJNcUvRo5cHu5MqfJHp79HLyhPmOKSjIB1eX4ktAYF6XxQjFhpAR9btLy8H4wN
eWDzDyP5Y1HfkUKzzXw4ETURsEDgpzjVX6VPHaxKQPi/GtJ1J+CQgtH4dMXF2Sctwjp1Rv3Ua77V
k0BYwCkfD3tlCBDpAQ8LGeUVetcBtNZzgGzICe6XUEKm2PxTwYTp1Ha32TmJ/JQSI6jsnmX5Gi+d
uo3VAFb+TC96lL5VeCzX9TcYtm6XKb+8E9R4Y9jrHpNxhQO/PFIw00dC4OOE8/zu9WJ7DDWtmhpK
VLzkSaFkjW2fCeIBtZlfTRaZRkxdL7LRV9iMjgRRWI4gsLQNpT7Fuqs911sDCJzP6jOvEa2yibl0
XwrhXYE9TG7dLKS2oHUF1+OFkEy8RvONxj8O230wc+rS971cuMPYylFFhfgaJt2Fo7RopLkM06aC
e7S1rT6TYhe5PZujjWfYzO3D9mMjFgWrWeZSk+jXPDutzeWpDwAGetQxsBGuVfIwBrC0qPuSxaqg
mGCf5yDj8rbTnBnB+rF6nFJtsiSAIbt5Zmyo+fa/1Vg0DKxT9LLFiBPovaG6inreox/fcVkcyg2n
sWOxdRL5nT/l2YoWDO6KjDDQbKBfOKLFstrT5jsm7M732RCjUMVila3xRvm7OQIN2b9ibnUoIIpJ
K3/sDGRJC1HT5lvIQTkP+WvSanFAol+6BM9Um+t/HabsZBNnt4UF51qoXywN9XiGr8TDMPk+YlFb
Pn3e3T5aGjmj0t/C7/HoFcrcMj62eeBDkxfdv6USTMQL2Q76rI0hik3pSv+bbxy9rlq6xx39jqg9
5J5Q5UNnr+qVzc7lp/jEpOMIGI3+8ryjO38rFru6m9BNKIllIdWiCOCbbeFWht19uTdpohzfDiQc
K8Mt748GnB7mTsadH1enfqxT1VHtomfY3kSTS3YdJ3plwIyM/hNnQJKwoy7hPL4l/TVtcZk32y+l
gaEzulqlgjKdSHejQhFG2eLi9iVqtGkJ9y3cQLpJ7XnXmx8n4OwFl7M4lM0oNuDYjJ9pCyLRa+Nq
fMczt9XoPjmXE00DQc3UZYc6fGedXEUX8aHjk49HIvJYaC+kguHbG12k6xmu+oQuFdgk0yAiKpLV
dH0aehXG2jIRaOn6r+LrdKTk7VVwiKCtxgtuTPfSZPWkJJIZlMsujXtLXKCCXLapxIFUa7pWiUW/
FxaJLURNpOZocv5LZl/3TXLd4IpfVC450h9OmWfPzM0yzVgK14RopZyJjlcnbl4CoNsJSjqURD96
UOdfbM6Rci+OHwDZd5jljIwTgRG1lBZqAlox/oUBmCl7jRJKAWFmvG5eL4qBU3mXjJ4VfNNs/gJ4
I9NY+cJ3EwcBWfOIUlwnTuqPrGIVFIS6p291QJm1MhZid9mU0uoMICPyuNLbQnVHqWZ4iJDuE3VU
YaADNVrFMRUF+D/QJlMXBDnDNFUAPRa76IZdGrZEDkICG6LUbTCY3/cTohlwUo6AbFIl67+3dXKi
rbjyRG1S06/64m2+99FLombIow2P+lEYgd/1wSscoUamQn9N7SVqutfQXIpqwmrctze1G8PPadba
KoKBvtM5TGtKYNirooS6p/82oyU9yO1MjNl07ghlDPCKMZg6KgvA0ZLLWqXMrKHeqKwDxnsmADpC
+s+db+iLN8/1Gif81yF9qAIOubIejsB+HDhp1hf8M0Scrg8/nv26U1KlGRG6+rGDRVjCY0AtIYn8
WXU2h2N+Gy11rzB437AZckdW6T2izp2P55z8DIkkfgDnqNobhwI17PD8OGABvc/UrhoGGMf5N2HZ
PU4HQBXpzZ/KA92KcGG+3wsCaTUubZs5ni63Q3PqmSOh3nKdenn8S8oTfVZrshQpOjqeShjxCwVf
I/r6hl6moTqZ2eazdVx2mCjcb+5iYnIyPit6Xj7CfzBs/iD3SVAgNAuLL1TzdbqQFjsypsxPJmp5
aAKCwvZSAZUWr0ClULN42lX02HZl3V21hqX0RswtUao3NN1evb84tKRCJ3ttNm3HB+8fWIqYpbSI
1cfxnEMVWsr/3g9CptfHfJyQDfoJYfj94GeJuxPLUxCymazbJm8ORakhAbVkDXdsTMGBTZZBKGOQ
0sKwuaW6+RsQsIrtfHXfAzEAgtymMdULNTin/xNZ8y6sdFr2oGpDDURa4dLS1NYq2sgmDD4RgSih
1rXYGxGLLLthLzDesiUkiTST/nQIBUk0kzn3PMjpZadUJPd7s+Gk77XKvBltN1W2xoLlfdWqVlF3
hRZJi9pMjxMsonqWrLXC5heKZokSGFJVOZKBBAlPZ1tBnM1hORnwOtdhw1I7rGVqYlfLFMVCo6rK
8kmwtvUS8JIl1RLhvuwpahEMeDjDOYa3VyHTP/+xLuLWhRSyweBjXdpRjh/rZYUKGi9+BozyC+dh
Df5BEDuIeTjsYCbq/Q77F2sUBaRS0JGNsD7aoeLjB2GzwImFDYxLdMs5p6t+/F6yAR1LvB8CynTP
KefP4cmP0Ws2hBbzv4ww58V7qnv9Dmf9UKKvMzfs2QcwV6qW6e204UExH3p6ymEHHRPiJA7mllG+
9pt8R3s8Ho0OFtMDnfitqRKbreN5YON1XB3Zhx1VCwA633IHXRLcVLS1zsoqqsuduGj/8Uv8dq1i
x1IMeypug7qJarTlwqcE85idhtDr4i+jh4r90canuInfaz+dKh8JK8IgNDE2MAE1me3eFCLhTYLC
ZEvE6W2RmM0lbygM6nyV3kJVThyMZwmDgQZxhsC6iiSZudT0eljaW3gVWNNOSy+Q3x6aQk8E7YhK
WuY/RSSGBLkvNze7XGlahKTCUiW0a9hxsOM43Voec24LT+D/n5AMF0X8wEgnZmj8jMvkxWvyaQpq
MbQQn5mkKD2E1cfVUD7yFgVKmqvuvuTLVl7+1zNuLstysoIxE/VbwHC2ipk8qSue4riMCmQTpGqD
axxrPndI4/Ma3I+dSkYYFpN7qONk53ZEj1Dvimwx/+jcZ4ITif/QQeK+iKDXWs5gUQ+hamWlViL+
I192KFAFOLT84K337RYh40bxZ0/arQ6k4QQLzl8mr+gu076UbpmLC+MAnM8uwW4wjLp4r9bsHM9e
WjLi6zSN/qILcYrAwQgzfSx9XIkoOrgGm9qE38CG0j3S5KMK8hNtafQavNUipkTkB2I1FRl7+Ibs
FIbqYDA2eEvOcn8w6pSSP+HkN6PC1ND7fwaVdosGVO1x6wJtoPcybPS2ctJdh+Xm+wH/EX2x/vMm
Hqn1xW75bJrMhRbDgV6pogp86aWVIm/sZr4bJZtmy0VzJMqIQB2DBK/ojEfG0N9q7DSEv3Y9Qix9
ACn9BVOEv5lUHV7jqJthEtNxqFTnz4PJ7KtLggMW4AMZRS2NoTP8rK5/xpVXWC0ZRia0D9qQtz4q
zXeuRiaWZ5+WSkOhVwSMJ1bDvkVFfi1kkcAvLrZVhEEiYuo0iObNQZzZna8zwmuTKPodd30zXOeQ
f4yCg5YpoBlN90ZgsQSVyECyXt1USXX9N1w15U+uUsPb/8gVbRoX2bsnNXMoXfmNd2jDg/RM7Tu9
/zqxDZOZ/t8i9KN1dQFiaB7RQ4uRkIBSu+BnXFOJRR9sD5D3A8ri2k9x4MW88Kz/6eMhZFH4ePmW
/wM/nBO+wlKa3OHZU4B+7zr4a84I25rYkyiUzOW3SeP1WtMcLof6pYhw1jb8yGHsP96V4UNOe/iN
X3YvnLMPK04IY4IpRS2FjDgdLlDbsJaEVs0AF98FSiDfLaAaw85dT06i7/7DmtP+H8L95o44+J12
XO8A+H+LMARFSfKAte02Xj4K34Xay5a8TvQsk+CeFvpCbsqh+L9704tK3d2G93vR62PYieL6c630
amSupPcOfUtkpLe3oDX9po/S/MeSlSKcecTyFAmifj3kMB64wm0659sTX6QR9c9euffjFT8Rw45I
dopBw6GCExZdO326yxQuppNUNf4+17d0zv1X1mjqLG3f0gaw8OGSevcvSreXpOOtDGuxBc9RdcUy
KQbMxI+w9bwVBCi5+va4/M7O43voMj6bm8+m84QQwXrJBWHeOI/JT2Hbj+aAvENEUaCbVc9mbqYA
ae3wZp3kSNTkL7fZ0Nd+Tzr7IWC9ExUhi62oVlqKu5F9dMbUJejU9WUEVCOM7IoGFz6Duak9Ppm2
2XhLW4AGE03TJmZ88+VoJrVJI69S5MaWxCE/pFFU36waCHsa6HJIDl32ogeuCyemgH0DPn42n4rX
/TWEyoXLjmYPGukU21fKyJsfXgCw1/EfThat2NGDvfDMUPxnTCQTaxq0kOMVmJQQSja4k/dUeRs+
7jdj/OXX3Sm7uMWkoAsa3rbTpwojvupWF3OVEzwxuU7nPcJKVYq00Emt0oqm+VHFdHiFMBM+oUFM
GIdEYAgDm8t/7Orz+WjrgMyvYq9Wp3ciXE258i0Wn7XA0HI2QXUlswsi409U141bynCRgkW3EDBC
JJeFTwNluVpJcHSsjHnStt6ylYvw6LyPFQjgnB3cmv54Tn20r2U9I7ihqd1oEWqaP6va9doVkTTS
FsNfCfTlljWk7V3kGreuCwp91rqHZW3jIFTn+bpURkCav2civVoLFqp+HyYj61bSIk77ijZnj1K5
K62w98ck8EAFi4xtxgsMZctdwyBFT9uz8e64z/DQsbKkZvf3oHmE5VTv+jiO35SygQQhAOdcfPvu
NoXzf8ltTs3tEJ0wW57/ararRncwSv2SSHmJquzsGwk4b9ihvxaGvlf4kz9MwEumy9mDS9Ky4oL/
yCIAKgN9OnrGNtp0pxo5ec8QoSxzpuboqGhn4fSu+oQ7Wvr0BN50WBHAGecXB/0EnM7xnNYS0hRM
gD/3rG3C3TCnAsWmR0csOpiG7CvtZnM03Y9rM5y0QrzUyRXqiw2TiKtE/kyzvaRjy+PfKECbaq87
MLPMqmGXv5SbSUuZH9QZNWg27gri0wNn8vr9OIC07mkrfxHNYNiz2yH15HzxV5zUC8ZwMZ46B2Fr
LoUVSRNjPM6PgI6HeLrCEchLQ7LFxst1bdwDNbzcFgYpIF8Kc4LpeEfWiMay4rTiiiz+fy2PLwNt
WGA3vhjjBZzaDUQ/IjktJmlqoSyyHeVQkI6a4IIpZbW06xJqWDPD6Lkrw6f/edetYSWO8rNStTMh
ELT382NSN/VBhaK2NqZHXQfQRzChNpIFqWprfFa3xKxi1g/jN9W0JDufGVzcQ8rvn9B9XkmcHya6
Yi0s92UROk/U24f9tM8QURHTpjMT2yaPtbgevrRuPBcWlBI7a2fL8IMhuYaY3TqnHvi/4JTmc/XM
mJbAHVuKWE9xSlEONsv5o+v7miwDN0GG3giGLzDPjrYV89e+hBoDDqEbJp026lUP8r3RA82RuBca
sFjl0WBfvnGOAqefVurgt4cEUotEYpqCj+/mt5j/LMUk1WFhApknJdxBcQOfbHiHovpgI9cZ/EeN
ERt/EnMOBCRZPbpPmDD8wsPAG4BMw5cxysbOUEpIrd7RokFUrOySNj3eV08TvecRH+fo6fPd3YYD
+pCabqb9S4I1O4+g7P8K6DhS44F9snIkaFiI6OPZWR8T8/3KRTqvrhiutMNiLGR7+nQSnAwaPL+J
J6wy4tyS1pUNEUvBsUN3FsJFNCQZ0qPoG/TIUkDBfOME//UwDtg6j/JMwAibuksZK1YSVvKh4MKC
zUcOhwoxoJRvJZxar6/jOiZ1cPcuwxB1BJ0BqHfUnvdGwTgBHdpiHxk4xUFm3U0LlsTJEuK1Cum5
4vWAl9oYiiPbZt4XA+3zB0qi54KSGtGvk5dZKki2rRjNUNRtruXCZeyfABzIzvSC8IsoZ/kvX+vT
MMIVCLj9VNvKFXQqWPJla7N2Xb2fwYPdLgRWrzx6UxmF+lUiAIcHohW73/D0V2z+8cxs+bdcxPEn
9keJ2w7waONiOJE6Uzjo5yFwqW8mJKa5RJD2W/9l9RTZER8l6QN936yvR7+5UTJiBE8DZdQMqtmK
SGBRA4kD1rsGl616TVQP4W89LkZakIhL7IzPeKRkhTHi70n7FOE50gtzGCcQdVIRZzQscZVebrt+
E8btDT6Ju40UBUdPEuVVb30kgJGuSpGGJSDgK+jNbmpY13q5WQ6WRvxayFFnOwj+rkpuFdDBfMRs
abzml1iEgHOEIOQCyVABUtyZQrhLQsogMV9Ye61LPOngUUI/hC3Tb931b1sqd9wUVpq89evPlHVu
cMPL8hNThECTBtXcUrlJoMjaOlCsDSQrr9D2q7ItNYcQqFJWeW98hZYfPlwimCag42/a4JhHnY+2
5raFsi33Aefw3XHz3OcKrPJe5EfsMNOlLxl6gRc78Q1LwRne95njhOuTg+3fQpZkTl3dgMEoQjjn
jwXLunLG1aXw9QdGVlEhkAUDn1BiFEv7eNGan079kd0wDoGSXyq6mwDR4+tA5lMpHcsaB3fzTvCr
+NeOVXky0vv5XrW4W4D7IjNO7J5QxRJ2lYX/8mcgy+kUY3YSKYgAdB1KDUh4RyAoWQ4lg+2TFlgm
To4WSvekUBXf5SvN1Sw0+WDPWkb5BIwwdzqcSd+AVcLQ+BClkkO2uJQTKejhXh2Yi6zL9GFx/k8V
BsrtBSUG1lZn/iNm8iJ1ozVijXikVmgynPvTBMWfhsRdYqAGilSKtASoIVrcEbFSaZRTbON5Gw2f
JVvZPQZcceUC+W96U1ya2k89lQBySV3mh3HUwEGajPIOgi0jkZW+BVM0VOR3kzF9H8QkWJeGP6AO
k+jmKEnonuf9h6PzxtaMDqUYICKfwbi+9EemQ3d1wiLwcui2yQvPfF+VpiLA9MNvNmfzFT/irZtQ
bH4xpwJgoLdZsmkUf7IhIbva9DwsvAVvboPaRG6dJsAX9I4arkKNeTWM9yX8SO6ghV6z9ocQGHF3
9aJr1NydxaFMucJV5sJHRy/QeYrcgNo8UP+NF1bxi0i3Ns93hDyKvj5vreN2Tlnu/EOUnLbQ3pcx
cbrapHocHYVvmR1WI1kx1gYENZzr6WxjKjCtbxll+OMwQY1plihUF1Twirvmb5XRYwOTo+FFlu5r
5Al63c9zVsxjtYXFpH4ntpAFF13UK5m5wwa2OMmYuKJhyNvF/ARDbyi9K2JWrQZvdSZf6Nc1rh17
e6oSBIB2940H2PIFYlaingorEgCIPKr3Xo+y+oJ6airbAQ0L4HpKmeS/vLkfuiVKGqUxvtrKKkgX
uToS4mHl5Rj8oocHeWIgN5yXYVQITWIRnHnoO/R2R9yvutZYGi9WEwHHpSzaEV3n8kj3Sbp/sM+Z
C/QkXiceiXgSEkx8HFUJP9awrNPkREAqGS/Mv6i7UMgKehwwd9wjVmXHoIZVHPz7CdplLN1kBZ4f
EK8CTsv1ZrxLjGiXmEGokb5J8HqSx+hMSq4+qR9NaGfXINaTLjpeHEvCDI+GOtPAvyNDg4MIM90X
9LNyai78EH23OyLqPWW+KFddWf8BJ63f+S0/QFEteB61nUoUF8T++OOY1boxixK2jdibbrm7U1rm
frRd6bM5tlXNOQnaFEuZFWEf6j8hfhI6usYmLate/PSAw/kKfVX6gicwCQ4HS3LvmsIFm8Pk0Y6n
+mKxtjrWxMMrCY8FWmkOZyGlsywZK/CERV5IDzwCPu9cXW1sQSi87NiDwp/liPlRfRMoww6/lBO/
YYPAvTy7Ra9FbPrbE3ku+8+33VpKRultQBpDyKSbUGKwcybkWb7my0LbJN97MZEB1Tl7gShxejeo
FmVmYulNoL2TeDT3JUwmifFDyxdoV62ST+Hey2QidZbERYTsENyE6WhNtjlKbozT65yCkUQDbSyt
r53KaBfdEwUZggwckM26R1hB7pnreriKbPlbfgRmtKWefDIhhwKoCNxGfyCpOCD0n7jTtppeIym5
6tvDtCXbeveU+tVcK2clLsmTPZCA00OVVrTBTVpAiJrg4vB0lvjbgERksr9NrdGIFGDoxmfTqeGs
bhnA3KpNk7RH1SpH/r+PEUJ8WFRvEfPl7fzwniQA7Sa6NTGqWBBpqnVKJWkgr0ihTFRVv5ffPr/x
A/VZvMkVHRK81xXPCS4juwhh6qNWEwGPB4o/1wZ7b7v1bt6ygNCMeC52QaaoOHaHChadiu8MjOtl
jHtJBdidkBuYNaINrXKPr5JPMa4kmsgcRK0GDgB4ieK3a1CzNSrR9kXff7M7Qxwh3blzFcqRC7Mn
5BWHDR4Uuv4mS68u4wrVojji5CoZdIDrWcatdBEdsFUjOWC0fZULzt7ivupmpEGNplmilZ7XySRo
lsErkxObTIv+W45Sao1MsjC8m5A+poswo7L7nVKqdH5NHXZzqghRGLBA1eROmBo+RROZLpDe1Lij
w82pF16mwVhO66KQNLuzzh77pA25JjiX8EZ8mIlbdVK4M2TDwLpeVCFURIZoZI4QIW1wmzD6Vc7u
ctrOn7bAz7G12DC09M2yFVuqVSZHxKx676EZ3dBjzMnVZnYbXT8Dvws6oDG40yr1PmLvDciO3TdK
aWZPrURcAKLnHF8y+PAOuor/mO/6ofub/f41RlTegujdkMqIuA5FfrONjYx6Mnf0sUUvzG7agPi1
kofxGmfCJNPvEXbeM+m22RI0M7wYjtcD7Z6LhphCwWV2HENPC/Xndqc1KTgcLcIgvvqXKyTUqpN3
u7yrKIMypvZtrWYnUb2q9BGl/HsbfCeNmNDDwt0BLj3vsbv+ILWdKbyEtUWlv3fBIVPLmhKQZgpU
XA62dIaudC2YqXUqY3XlDA8/imEycwSggJDQJ0Kn7KCSLUmFM4VZpUwVyQDfMFMDuKy+ZMyF4Ejh
owuKMdelPaId8C/r//Quji5BRpVWsoxhldJ4S/tWUKz2o59fSvGShdTTNODwwqElaiyY6YAu/7NP
STFeRGnXoVmXLe7uXGn9PiJxwzUaVBHWB4gR2X+6qqMh8pMEcWHUTT/Odh0t8EofzJjshs3Os19B
/QMLbKvWfxOEVZnqwd1XqMhwZMxU+zUh7xiju8rHRetQ0mAKQ+wHJNts3j5SeVCCnSNb9xdisNHi
BvmhlQjRO8adRaIgHUFvJQwq5RqUL1WkLuL3d8geQfvF7FZ2sJZMnBlUQ6eBgN0OErNlGh7J1HCu
CgUmNLwtQ5zUQCzPcqKJ6IaMeqiOd3yYzEcN8fqzotcPbcN/P0Ty3HCi4MAB1sdFu0Wi4ZZ5z7zD
Kyo48x9yQU3a/J8xe08d0biGVtcwKJjIoVU0OMALbdflbZCg7dbg4rWm2+lHddTcSS3LaXv2znAs
PCP5V+5Jmenr4FSaWfByCTV2lfPB3WRwQgEs+4+GZgreZfAYh7kAJWn4PgWxMjVdsNFeUYsuVcvM
MXcoVdE1UwOphnuP1WyONjSxWKq84BYIsUzpwSR4iIFZRaykqP/GEdCynnWhR/XPleTSiSq7kdKB
BSMLk1XOrjSu56gRx9jh50781YQwNCHCKPFw8SlcJ1h1yYd3FdOOzIgjT2vcaPwgDRJz7ZmL1Vux
cNn9ntC2gX5KIgjOO24FV/Tu6SUDxWttl5/CnV8L3jObFj3GwmC+03TjgO0mMCiRQSV+u95W+Sgr
meeQV5+C1I8kQZIWENYeQjeeTU5h9acYME8TG4UTSaWIVCr1YhSMAo2w9w0afXL6AaaEqzi9eon7
FLLaBeI4956PjKpIuPDz4/esZrrgNHreQ4XgBTjLHdMOX3+AMuwTXlwc22IYnsFPdWUy1JeRgmze
k8bh/GUIfI1NpqsrP+VqjmJS6jUKIYTfTUw5zj9iJv16LzyHLtzRdgSqaBtnPzjnBiYQfgWdknTO
dVWPnVjbshdaYlszCdc/t2CFhSy8ROGD1LZKhGmb5uSHHGE8GR6mRAeRE3tmeoPfhQ/AtZgcO/Je
WpJZMe7Uq4MlKarP7eQ6da0amNeoFmNNtzjzEAj2w9oQOe8WDm7H8QVB/AxVU0taW/1syzPopK1Z
jOous8MaMFXjfXD+vFxI05PfSvQNICmKtnpesWqFUhNgifI2aKdNqkuYyCs0xrx8glUnr24CJviQ
sieUPhIbBTehjyJx+CHdv0cQpYqcxu6VbNxRhdXE2TCzTsBcxgVHYzS/McnORlWQdLfnkewDUEFl
XkQW5qzLyEc49aZHXLYgLXDPc7xjxHOGAzk1aGfSixeIeHYJPLD1GMX3dY1wdYZHiGPCoC8ULNin
9HbCbF42lEnA8S7CGZtswxNbWyzM+zJqvGnfsOGM85bJP/mxSwC6UpvT6b9zwYsqrGuF7pyIJzz+
9n8wcMwtksiYAvw2DXtv4Jf25VXtT1oQvEs3vXdSTFHkSeJQObLAjVnRWEHJRD8t2rXnWmVYKWtk
7Ml0gv+d9aD4Ryj8GR9+ArLRizombypcvDnX3NV378dlvYZrksIaGM6vtV1JmQJaj/0QdaI3DB/+
szvh87dYQg8dtKhpFBwqyKL+c9HGdNu8WKaMcSMmkjStAWEaf9HZqReLw1ee+naIPp4pCKaf5i0R
3MhCyIVra3/0hK+aNNNotygpOptW/JKiJOZMsDOdBuJinALLAi7MAEbek2gXNnLi8W/reVlQvBRz
yx23OXixbSyz2ZCXIn4lvdl9hBvY/eCJs4Ho9CfwbMpUnZvkANcBYaZ2T3kHF6lGDaL0qCMAlZWR
j/STgR1bsZuq6zVUU8u0qqDu9zAKtwkv10Do3u5x0w3WLZHAPvaJWviWp1aNMinTNiHT0nrUmRSE
sIUl28Nh1fhMO7bHfRK7CBMx0ZDOBGQLHiWdXOuvD+HhEzs/fsXN1ap2ka7nRX1SF+BoR6KJaHet
WhE11mVPKN5R5FsVgd/9zk/DS281nYWpBT3Kni6tKAczropNP878eXpyu6Nrbw4kcprwcapWfNAx
1JK66+GbxNew+aX7yTLlZbhnsyrKY084P+KIuKa6tq1mH0IexERt7LNB2ep7TU+aO/hHfj6PuWwe
SzDC8KzCF/YxXeevEys02MxvtVT4ORsag9DGU4ltUnwo4t5SKZZz/Gx1twZr5sT6KX8eb8GiRRWK
Oxjdm6eO/nt5AnEQRdzdGlXJ93oIoaOLPS0mW/54d85IypEUMzRT3FVGJd8TFL+i9R6xTZUn8/ac
+U/HjxBGXoZoRtupXAtPcGQehS86C191Et2iAiW2YNu1LmlxjLwlpfTow6lxtbG5YcZlW5f83SKt
oE9Hu/22bdRhd3QXEjykNrtXZF5HjSb7kLCM4qePboFvyFH66+UGxmHzpWHC+GbmS/VEv2nuWH00
W9fJBVq4irhiCSoD69QBFoGJocB6+z4P/XNgRZpNskMUOjmmh5yOlvb3qwak4LoBJ5rracw3ZZ2l
qjHhj/oW8J/NdBqTn+2IIq0OWy/DHEiB4a1a60dyo/eI1HNxDfHmdmXxEFaBpCXlWdT/oGBgCAsz
w19orhcKA3zJo6QbP0oyz4hSiCfdlNwGMOYqIW3mx5H4/wxO0RnTprmffwo8TJuNoL24SMKIGrp/
Zlz0r9mfL8uUFewe4fWi+yKzan+TGh5eJngDs1ZMFN0MVXIpetSOw57fiIkjbc7lGnM9orKKwniZ
dTZ97e2OZFY6K/FsDFTJ57lGhLlR0qbrefE9TEqjWd2/Cfn266iTN9Rw/vnAw/o2jLnDo9MxzCyy
EECe9xIZBgWaLaaucyz1O4I6RnZUFwz3DPZS9E+QBdcDzc0BKdttDPp2dZRphdL3zKkm+n9yxdG8
Tsk/54xUNdj66OuHVYs58l7cneRIau5CUT/ZojypcbhQWUjOoOpftfMxkOWqVzLq/vqT1pb90kJP
3wwur5LB5Jmb2LNrKoR0jjsx1RZDhIUx3Z4YKX79tymB1A+IXOsBaPzzosXEhWZ/d1R5h9miOP4q
V//ctlU+ifaKzOt28ZuF2sByvfumVmAp9whS6l3gbZfLqJH4gg62QZLCg6t1Q/5uE57qozVn/tMC
xqMh7jRXyAbpGCptgsG0CZ93zrdgRWmMlrPwGsjpTy73K55epBIlEogwhFN1j2D7q25yQf0y2JEQ
D5g3PtJHPfGhV0mx4VQeLOf/DAR1p9mMug0H/0ZcLAJ2BLBlOu/2BysGUkjP9IZW8xjjf4tRuiWv
kk/2g6zL+sVeucuCUNG+0aGB9ij9OQopBjIN6NQMbO/cYJGtf2L4+uzdpxkCU/8fcx9qbGD55dLr
bjfswU9T1PJ86ObNwcfmXWQWpxS3crn+qkcOkBVPRFjAul3ak7tiCzSUgN9oUSAszb5Hkix8SGrV
VxHuU7r0ZZF3v1F2WTTOWiDi23wvww7ocwpat8jz8sWBxK5wGectrDtIWPJpZUlKRwJlcmdZhQ6A
OWYiKHkCH0rrHmIE6esb69r/28U2zjrlU+xTiJTGTfXuB9fLtTZIHYLK1I89LgH55+KXM+nH6Cvm
2ZoY/BMRboqHMKLW2Y5LZiFFnxIxOiWMEVG7VsvACP5QMh/pbue/SlX3J8rhNnBPGHbyeG2ctLVL
v2umg3UbC7g53Bt4YOjgoZxU0+tjWuCl/ktLGD3RGZaZ8wrNZjVKDsl9rOpDp4LtMxF8lmKaP3eP
GnD9HJDOP19nQJg75hIUPnQKTWPDDt2M+hX9nDiE6X+ejFqwph2abIhxU3SM9OxMyPKNKAdcebUp
tdmB1D5CJPmL6QMsiuDnK6MYmig7hS2m1Uu1r52qCdaO4EtQAKx9XU2bWHWoWsk3Vc1ZUeRwZlNs
wsOoxvpAUVYTxUW505qvvyLiP/C+d6Lx29lzKgdZOhCYzPlNKnd4rjcHF1d+iCTCQVwUPR0G+sTE
wVNWbWEvBkwBdkC5Rota7LUD+kVHOv1SA5nyOAAo0guMK6b4bmtYBKBU6A+VIzC6zMnCjUCL/rje
KktTkgXjr9n9nVgrizrpFCmuGLfiN/rbnJPCm/zH53zOKHS8mMzYyDLCrRmN9qbyrqTw8t3XhRuN
cdUOuuBamYYWwmFw2g/I0IZwT6TgcH63+rHUbHo7PMsFSR01zFdKeeesY8ip3Q6ovV8/2c7g9KZo
oKSr5pmSXRx31MMHBxZumOm4VQB1Zb+yKlTALpbEX1f9SOfUjocuisEfI7jU+fHbSVEI6uIras9y
tyvC3dieYgymNSb4bfi21QxbQ3BKlnBXsZKN9Oh1VmL9dI7GXP+atv9R+Olidc+hDKtA3eshVhqj
+J9i73nKWotYhqG8ze0/kVbk842G/B6CmtQuLA6CIiQ5tvJhROqHP5GfEbVpSVqluJk9yIDwDJUo
CJxqdGb3OLiH3iBK72oOBDO153JWy9OV21G8ZF/yxrdW+eBb6V3CwrkV1J9lRyP2ftYM1fwPmCOz
F7RUs9aAmiq03ABo1jqtEvW2FgGwAuOSp1gcq5PzByIjVmit5N/V6Ol82YNz5p20UbuxCBR1MgPi
z84HBQ/WcxvE/TnlFkMOfySPKUTOEiOWopBBDiaJGxaxUMHtAwvIfby+u3d/UpJ7MG6ePxV/Z2pW
yeMFkh1GPjjOQX1E0oDqnZDv/jw+mnewK/PHWylUnd4WoGXvA75fCIqb1bpyJ9Gw2PsiRtUOrBcI
OSqh1atGkz/omriIchvXOd9mprRJ7prT7eZ4yDtrOsouOpYPqHPtCQ+6GWsIttl88fKpTLGnsOZv
7arYuU4wrnmbH1B+6N3/eU9eMGYbHJYi59Yo4epF3Kn0L1Q9znlXeuMFVgT+ahlLOQMfA8RNMyVh
7NlK8ftmIwDcS3jhWIlEi66lG1fzGZvDc4S2sbf5HmCZJnDWHLbGHF4z8bSZ2P60nfpL5gmbF4g4
RN+LPZfSkyxFghdGgqBYu9C5I5RxUqVYm8bgC0HVgiWKaN0qnKd2994YwyP3ULn/eXWPTgVbDODm
lMgmtGvETrCmjrWvfFkg5lcNChE8oWQc1Ik23v0J4UxRHphqJ8V7glzhr13pDiv8MbaRcvxHeHlU
wcg19mVh4Xkw1mlvE990DEu33R2Ph40NZzSJHQSiFJ/hZo0NEUyPOQpPk/q0LDf+ObcXzBEAA8aP
OhvFTxoiCrD+A57/3UbbMQwSYmLvYI2IyGIk4tOdh4/1NJuxOvvIc/C18VWkDlT7HDUHTlam9+rE
5MFMvSyEjq4/bb8C4pmOTMaqBDV0XWNQzcS+Y/Pkdd7ZSctxvjq+kUkK0qomKIGCVQ6P1O+DjqCF
Y5wa94iBKpbVTr1KGNS0L7Py9O7kKGu3P/8Ais8kXx11H7pAClOE7R25Ul1YIYeUgyaqD7FObyEj
Yu315ITdTDL38Hjesd6UWIbLe8LAbrJQGOn7Smf0e+BKRCcgpn6BYWyypNOBRxCmYQ/PiVCbgzkQ
2d6G4A+BtgukxVuZUCLhMkz1gVemKPYQYW4QNjFCi6zJtqr2DRHmn28x8CiSY8+Yy5e9th1nVpPf
w8Mf8qrvVTSZd3MS39/wwLfYEgWaCQXv3PAQBkn9fn3RLz1SbowPw3MIcarojEJzuwbVeNYyiJly
rk2hxEphIRJwncF1Dmw3pID3RCFuL0f1zkvmaYTa5Mc402Pr6kKM5ajkTnSTLbabVufaI3vMS3qO
VKq6AAS7f3i4lHqCq68bf2nQ49taNOw6wLzPG2a3YDZxf5yB0kO7AKTBYjboUEH7TUt8/AfXjmO1
z60dp3hBLHlG6vflKVBtMXUCE7/0YRgFvEDxYzZe+FV+Gx6pBSm+sN8xO1whE34AlUsmcw71U0JK
nOT7kYtxHcKMpabNfh+caTIWBocEgKwpfPFm3bh/BA1ssP9kxW/9/g3+JBf5KL+LmTURZHnn5Tv3
cSMq1GMxtPkvfBK0hvO1otjz+cHpcrmNq1DFzwvIOXWt7urFlLzFXUh2KU6pu83K3KiSAXylW5c3
G2mDwjhtFW9rDX9+qtoDyjcnGOueb4+dmUts3dMlraHdx5Vh+NySbq8DL4yvSY5qso+CZ7aFxJp0
p7WhJDAh0NH0EFHWXfDI9fFYVCqrmzOM1IfBgj7ePITk/WCOVXrTeS/hHVeQqgCwMzjkPaax8VWD
OGG4oYzWap1fhjEF9JLZHC+gfmfkhawQwV0h/z6Rpt5tltm4T0G3m0wsjb2zik8xyiED/s3OeeTb
s9c3tMvoNvWID9Tq819J1oUTmIfCUJ5/zX+m2X1rGZCuQu+9LDix6tJThvdtRvK4mtkp3NjhX/PM
PuvewY9bvWahvCAieVAtpV4/VgRVMZhtKvhcOumHlDLF6s4uoVoU3DwXN7JboQXkIPIoutpPqyLM
uMwZYng0f+94wp8T/iP29CEPSTJ/yNJ0w1P5M4zu2EleL58EiQ3eU9SRydSmhtW4mnOC8I+ILl6u
EIdP62xArhzhau8Z1O5y/bG6KyTli0n/ZuZeMRMBMUYYo+oibvZ27tRmo2koAcgKS9hANXhn9zbf
23f5nmxfgoJh+RbXTQL4P6DuqJ+4xafup6UwbALtkMGNWeKYHCLAvX+xpOzND+B1s27icXYgj9J5
Sal3njqGYGHfAYAvoRR6Pip8lDK6gY2z6IlF+5s2i77h1bv385UqfzwJ4vj2euGisa9ObFhfmJDy
Tbk6NGKeghNNA7xJS3/SoTH4fmy3EyO0KLxf/9VG0nFJyAPFcGKrPExt8gNZzaD900LcU2rQsEuk
B27Blel1XPJpaE6l1SGq9lZuu5aMQy1AJSd3LVX3PPYfBeHNu08xPhy4tzt/dP0CdFVKvTbnDkgy
ZWABqa+WXUIy33q6eWKJ+SKkWFDQMsbTpa4g7k2wtPF9TbPzqHt8n5YsL+xN97g5lWoO2ZXzF0VW
O4ISOctkNMsLk3fRlSY9Y9JjGZXytL2F4I6g5oaMlTSbdyhoUi+2jQ4PNQ0K24xHZbPenO5xg23Z
NlOs2srJ6+RTfhcB58h0yFdxKq3kOeZPDsPlJ1qU9pssripbFUir8gw4viqtiODMy7P6/b2oz8Fh
Qg7bDHo99uXzzZTBd6bHCCgVJq5zFP+VNm6cXnNWl2lpEiXQINhB8tl3hXK2r32+U/72yPzUSNRP
pewm74YSeSjtXT6AZkbExk7MfY5fQjs8uVQJefgZR4srad/KVsf5ipirBE6FN/bDv8+VKgCOCEEg
m1PznAQMy1UUUW5Ela8pEe7r1NSTv04Fm3mTbaaCguiQyZgFZ+jpMn8sHKWoDGYMDVjH2VaP+nib
E0CiMTuFC0vhlCkC9dGnwPV6te/DjTYxm1/UbB34+3hlJAmZ6+SYT0oSpKFMdgdC3ZkHlD0YGbw3
2e7NGGb1muwzelulQbX838pNKZDIQip2/ZFp8rgwr17jDdzo5c+O8foZq51oL0njEj0Pv/uODFAo
PUbjmT5j1BBjKS4ZFQl2WSRXt53bnYcpP7tzLPkEhVWXz1SERKlAku2fsaaGpjbSmVBbjIZRE6K4
PdeP+cpaLBTFIo+YQvi1B+6FD0BFl+/z4k5jB9MTWpPrTsUk/SHMHpogGMsFZJSHwZYYq7vb408f
vXr94k3yFbTPTTLzmWGkQrE1eDbC73lyp24BpkvPu73TEF3EfhDYd5bmEQvAOVS2w4scr6dSWHR/
PkFiY+TKBUvFLTH6bizy40WMr/Uody1f2Rf8sRQNa9PIaV/dNQovwanyToAcF89kWm5j7PEccrW7
Jh2un8n8Qm3gGs9jvfFWRWyrXkBqflw/J0xfuQMYi9Ghidsa+FQEXF2IXPquHUlZ2stHUgSU8BAC
7yf2uo2ME21Lxi4YgJwvVJ/5DsGJui5bIZe5bwQrvG3X2htfCaDAGk8auK2xtGSonr4Gp0EWtFrU
Iq9bz+wr3lN/NR38Ei3Q9RRs4FLXDRbsUSvYDoIfpggtHBGiVRrgyj1U2Yv8TUbwfuGfiKHIYr3+
V+2PcrPnSIcaYLRUY4po+EfQOscW0/zvlao4vBTIjS4milSGbfFm4u8b5WsVq80ywQOfwsGP5517
D6Xg4l2b8KBaAOyOVXClzbY0tSwkF2klFI2kr48KaR+zmYl4cRIaE+KlWnPrw2NaPqJb65ADOsGh
vch+n5Mvt5aETDx2MTKbAB85VAdqr34+C+Xcvw7TipEpq4cHT4TjuT/rSYs/N8qe8FF97qSGmEac
5HYZGCN13lNRWQeZ+wpm8XNUzFybxl7Sq6/t0aA5C0mPA7wSNdR1e6/3uI8qeJy5B8+C00WmO/Gg
FIuIB3/BBLmdAUIiwUCelvPFJOXBctJx5mlONT01tp0ce132tkttC2zyVnaWC/jTg4vXGMdiSDz0
eOVuhPsLl/e/qFutkzX+Nymv8ZIwunLvtEtxRzANyPmu6fjdOpokPC3Aq6Uzkj7cmCeAH2vVNODr
+pUwWlxOVJNodFdLiBrNzXyBvJttJdWYqxxLCb1vJKvvqXzNUnc7v1yzbw5YhD9eAYQAlbEgPyBe
dndSBjowZ9W88Ubt/VqT9sgqlAuSey1L6c+Kj6jaY48OCBhnJlHkc8yer3CH3WERO++oZ4lGMbJ9
pmBQBMmvWQNmLFtLY4/ZN6cXBtBhcSkkLjoCs3BaWa+PyaQIeISo4LFuhnGcpcfP9BOgGQgx9vCn
/zOzVfU7H6HFVOgk1Cr7LOWZd0Iv11fVFzqZC7RHRt77f+1mMPYozcbBnVH6zKVq5Yvt39+5jgLt
hittBq+dctFvCwhxnIKnuEUjkCOmTa8cwvxhYBGofPG3KClj1548V8GJ+JCd8HZcWiBsRPLbTzXx
MVW1RN8DvK7fwywxzgxhe3bWluvOeqlxyAhh5fzyLEbFpZZRgVWUs0bhwEKNABD/lmgZ0q8GIHEn
FRBEUIcTcHtSQ3h7icP1Bk6sxujX/LJibMaFov/znWLM2DxxWTVQ8mGMtGn0aNtYDqgHnibPEXNX
axULngT0X01Qe/j+IkcH6RrEfYoX4GdqdrE/FEWyLCeWXhFetHjBtB00hqoe5Nuz0ezqO16t9Em6
MDJ8YP6I0RMXhFzO1ARkien1XWASbBJi3JEez4AiVtydP8aEMHsv8934zWwhBSWEjOAwZj11r26W
w4EXGC93Qo029IPnzgb7q6AXBeKAiZfIz8gUkABrMSSXxlPwqs8rwvRdrq5eoFQ+e8zrUrvZkrGD
56nlt0VF7KWsq5eU8/uhVIRjBR40Fl1kLpDJ4x5teH/GgZRUXqTfUf3J4M34DhLEPYdmrBYx4VYj
GNJaim56V3Bkw8V5TgZJ8xpvAX0U7Fwdtvm9AgbB3ySEFt/UPF7CEzNvLPTq0RD11nQFi8ZZ4xTX
bpPZeZT7XRrCut5i/5fXWRDlF3BMdhty7ZAS2mHR6xarDVXJXPH6q5NlSUVkP2il/fH/b8bxktQ7
y/kGZH76b1Cj0al2XiOsu2UwvRwke9b5eioTfCb/77Ou2FgUMZXkfpR6jRWU9ZAJAPC9rEFD/EDZ
E7iAFB3YZ810LMqfOQv0rEQmnet2YKwDuVlkf2esOi9MP9GVOdF7i7AiKxIdEqiPa/CuyxHOmcwm
uEtulWZTW1t4sXndC60j255OK9FnKmVOAu/xoQNRXqqDrOSoTOe7+FzVYOI4xnS4CPdS8pa5GAvb
XRRFN5kvJLv1cgofoIj0jetVQBBUZYT5xks8gcih9OrLF5dMnbnnITaO9jutbzgykyUMjhqRFTYt
Dv/7jGHziYh69aV39K9nlSreyMh9nC9uCa12AfVMWOU+fY3oAJH84snCMO6Of9bsVguY8C1ueZxK
pO17koKz+TJFPZ4MqXxZFAz3eQTueoBC/mLFIjoG/jDeYj+ch0SeKTWHVPRGfBSAzvJMVJzTN5oR
VVS4/q37SJsxSvav+4q0OiAaUGVy0YqieSdUaD/L4oBCS9R0wvScPozJo2Ypc+FMx0s1hXO604SE
CBpqnsVygwTUEweb2jNW7LqUh1Cc2JLgDdC+0JJi2Y49DRR3kcE9nG40OgQWWcUB3TrtIB65uOmV
Ff9MOo97PMYO62/GGlvmSNll4SOjdeWzBUTjMOXRRZhlHdvDcAMbn3t0RmdfIgSN0NWTk1ykgTm4
YevQXJhnEZwM+Q4wzKdEDhiULA8k2AFn/JeZvgLxpqnpLute5Pt6ky67lzjm58qVCrwqm5eparnF
JBxI/06WCjip+v/X3RAn+xMbk59oHam0nq07JKLTwNTXq8qLS46zgzkd6cCSUdrG2yoouqpB15N/
mOOrFkHxv+3RXKjx6EjYHweFg2LIgtRV1cDPR3I2DA+J2r+ydhzbX5C6UHUswDdmGDvRI1+ciTHA
B43gE323Cl2s3hgdkiWGvRmBG/4G4r+/y6m1jXX3ynlCFrcElltftbS5dXlb4ODdIH1n1195uK6d
8yxn8X/6KZSBIapmOSsolM0L7tMq9AIjjS1RLPTG+Z2Do8fCr/rgEZZUBUXNvq10fr+vUINJvtjv
VyIdN4KSDXLwt71MwL/7b4U7a+TyVeM6vJQwx1pIGZeSwQc0XOwa6kOOS64E13JBIvGQi75ywnL/
XHL0lVpbAdNUMv1rufi65ehfe13hUkJgJLAXHj8f8MjSJiyXLLYk8YUh4Ois+c9tY4YOvr7rr2lu
XbRRrLRmfshpoaVspZtHxA0knJkGJrTd3mAG8Gm/jMV1nsSzqKk3TKB5WVFRNPBYqJ2qrND5ojZf
O9CpXjf3VC+Fhn880BVslz5Z2ZZMxcGGtNsJiJE2bzy3pfrgwOw9rBGEtu/0fQifzHMA4TJ6YuLw
nK78alr12ncPm/Y7TnHZbhG8lzJEoh3uqKrxaizldCn/+AF6cBrTl8tMq9UCcoUgcfmTB34xHb+p
7ThCLROx0RwPlTePSp8MLhliJsiDQAPmYqcmPX9g7YWsY8SPj73UyuSilnQtGThqYt03MI6IXiON
uE9fPvTFCmSUaS/IxhihRwYN4qdG3K+34AT+Vn0F+TUfpTgS8Bw+50Y8Am9VhExBjz0hIKAkLbJW
2XqxW8DeI2qhbwm8cvBK2qPWwHuiS+Lq9fNcLuHfBnPMe+AJVxPan63GeG2cBo0g5TNwUwsMT2kL
dQZFtkIr6UCxOxkYpir+SVMyPXn+mZIf2551I1pkVjVegLoV1+A9XgNw4ZvqeJVsGYrWyauAnDc7
bEYUU7c1b7RGHkRpuhLj4LCHa/+Zka8qwvgXCkoA825/ZPYlJ4+lRHkdJyL2TDLAE2jdzVSpfH3l
BfgsE/35Mo8aAcJvQagK3pKbrn49foXQcLn328EcOvvZdMwj/8ZzA7yfNRMkXiObauLpSekEJznv
pRH7KH+H2cEJEMHY4JWRtg+Y9HOtKDiak1Yg0nAcutHJW9+GjYWNkNfcpESHpTDPBJ1ESqiWovKS
OUnebiwwK/SMTvvFIUH+h2i47DaRE8guM2l0aRp8TCfUZgIRZka7KuPjcxQGV45kXmO1FO97hHoS
Q9pbd6F34xPqEJHW5Pv9j/umgXBSvS0r4OEKF3tuHrKEyEBFpHqzMxGLjaGQoCsKhukhCagCT2Z0
iNBB4AUBO9iPm5VNsQQAmcUZPfGAKDMRv9I6O98CYrPYwHk6mO3F3Sbl2yXB2LoiqzUvnG8H7Ygq
Ok3VrzblBJ+ZaQ6qEUZNX/0/8S7ICM5HC8UzpnskMdxAnmME0DnmtD74+VAbecrHtwwUmjKUcs8e
Uj3aJhAayGmTkmircZy9p/zRhM0RVcGFdEBqLnkmTnO5KzfrOMPfUnwnrYfD9f/wdkJl+QofK6IL
5cTK9wP6SI7yR/2PZAyursVPHai9x4YDpCXTE2qlDJkvm81mz454Au4NNE0zX9F+NalxIJ9FK9OS
cSaSoZKEv7pz3pQF57ESEOdEv6Uhb/LM1MeLvCib3GJLJtikhLh7mwmddMb1HTm0LGnu9IWZoioQ
VD+ZwgWDw9FI/FYRwC+/JRYQF5DefFe5v8Tw4yKZYK1OmcHi8OxpEnqWAHpSaXgQ1gIIjvhuHjMQ
EHMScKrcg/3K8rVuGX0JEcwQmmhiZk1YlMftRKh3D3tVyBMfptflD8nN+vONEqtUEDe0DuNN9HOP
rHdXcy5GH2nRwWQrh/2CFKuAio2mncDKhLjm14SH5OOuwpmLPhxijNr1ns97G0zmt4MS3TvzJE3P
cSF2wCi6HtQSMLQfNFW4eCdzkIJuYchSkS6s9j7Zn8VYjyhstRuEwFBg6I0sta6Iu34vN2Uq8xf3
3wROYiC4x2WTguziAc8KVZpE63ZLuZTtQ6+mjJbDZWzJxqe5BcTqikGgR9glC14zxO77RxUXVY56
HS5NbtWrga9NWZd6tR1pS27BaVuZgKaNX94Hm4n52xuOI1x7rNYER80Euq64IVkqI21iLJSUYJZc
T/X+85+LgIVMUTWUd0iKuZLD6F/eqrX5XehbjKNtzpV+TmtByvUYMJwZ/jbRtBriODZDH18/2XVy
w3V9XNmB6bQ4QX2zFw7QTt5PMsMq4Jan3emDIj85l+tDCJVJx8vWjqA+lSnlNo6PXnZDcIZuEQrv
NMEdI0K+TAzay9tC9iWQADxiI8TiLosUy2P44aF5BNfzSOYmp23gRc4kVYRP9/sFiqctyeV1aN0r
31L20KFiN0PVqWPXFXPTVkuo5J2gQJNa8ppug+9hkE7Mht+Mqia8WSgsjboT5+nntEaXF0+u5db5
clWVQMR4O9n0k4RSYQyuRxO13mfK7azKHkiJ97Ori1zuImq8VL4qJEz6TfWZojLh7pKL55aCnQIu
eT3Qx6gonG4UgogdRxYeoaRqwgAgQ9aYWFaXDykGa8Qrydd6xVlW2aOdims5DhxkpgOdb+6KxN1E
WAG4lMUv/y9e8FfLObpYYo8xSfkBXIJqInY2qmxha9HkKAmsajT49lDejCGxIJlOqzdEt7Fr2oKe
1SumZsiy/25xbch+4ALDh4NyrIPIy6Dm0hd164k92MZbUrCXe0jBtj4gSsCP02RG2V04EfEx2+YS
Uce8lG3kcGi8qZf/Gv4/p5s2FuJ+3hr+zTlUc3+YOHgBBND2/KSH3wsqm2GwQC2uCtgHZj7P9dsT
Ch8LjK6izRuXky9UOys5FYWkHrzayxV0G8Z69bojDEF+xSiKyGwKRo3IURKyVB+KwuRBI8FshzNc
TNmkoGWDu2aDnKVmOvNRF0X4L428gdPH6VZqhq7G9dwubl8xAsqL2lmQ1dRIBuD5b2eggtBKYE8i
SpzyLvEZal41xVW6BqJxT0Z5s4DMmPx7/4O3L+b7iqGS9ghFFBxqRQ7o9E+FmiKaiKqMYDwAVQBc
A5CAWiBu2BVDhWu2I+2Al8GZWCUbzvCs89m2LPAPLNO+TpAsJhHcpxe055FFXuiMmEHxIBoOgrbh
AQOsSD1Brtb1OHW35lSZH7VINGL4hzEdnMz2kOE7Ip4ccm6tnEdj54UoVqGwi5X96KpzISkPKfHh
Oh4x3BPSHH9Ja6GKNLAQOHDxxIFjr1jCMiodPLs+Cf4F4r30kWWOBVQCIOSx0rynaTgaAhIXu5rk
QFfB9c8K29GvKisVbA0YRmx4OL8+TfQZnPexWjqzKajb4NBxPuXkLuvgljm3vDSj7MNIWzkvD+Kf
83eEAw0KAQITQS1Lssgp00uoBhrbCt1GYRF0oJZZ7FgXR5tz5yfHAe8TGW+1VHcziJoPC0NJvIqw
MnYTODpCcN/eOK7D/pcxc3Ohms9xhWlC8wd8Qrahn8tvOzqDL9zhkByd5PxCgiTTnzWkGxGydXaE
gmhyKi1J+vaZxIiNYNSzXq9Sfd29jbf5rYhiSRbcMWAUfGVgCZB+hM5JM4/a73AVTsrDJJOnTjoJ
jPpygk61ECOdyQfvmhs17lim4gg/zrQqK55sMS462dx2rCa2Z0nbUCJLxhAC09k0Wz51AOiWrq5+
yGVfJ07q46vO7cRKgtkayqFnK8grt+8WnhXcZOlPU9M7knC6BD3Dx3CGuP6NpAzIe7bPBMVf8kwV
Ax/nsdjEQmAhMs2BRezb0mhkHSJdh1ireARfq6dlBSCzW4RgM18+d+E8DNPHFtQrq9Ra77g7l2vY
VX419UlY1ifBbe2V9oVfzaOagnij7b2kKwgJg5xlZwURWaxorWwVDFh1kWK1EsnbgBluDNWhRtHZ
O7AvRc0blizOMWkXkuOgWj2/b5TAivS0/cHPkciyiwaI/1UrfGrcSND6tkueUjztonUJAOC4tZFc
/srqVXecUlnfMaLpG6uuse9NcEQhpUAF6215XZc6NIsbwVFujG0IpYQ5x1teqTEKqgEQwoGvO0Uf
90xBx94rbv8BmXrwi6VNe32mn3DcKGGc5z8p6QBBBsXM3dSyG/bPtRcMAGgDpfENceaiiE6JxNbB
8gn0y4v2Na+u7bp2pOd8GktwOkwhtF6+wesT1Q29rTaWBFN8s8XvkMGLWB78AieFOPLLLGClSNY6
jpbl8nVoarMoiT2S2beSU4p3Lqhbvcy7g0P+KnBOE4QEsI0lRnwFzea2ulPd7ut4WINQ8XyMZ9PD
kEuZ1mm4oe+TNcfxlJbw+WPbB+5h2JXZzw3gxJ1dojxuX8N6VR+JlSO4zG63H7aBpJMHldNVPzQE
rt3v7dqSl79IuNy6ymYzraaKpbRQfIthasQaIfZ67Caij5mfGvTqXLms6VedbwoUPNlHUuzb884A
VyOxkKmqSftHPgU3ZDdUyV1YuzgY595f/V7j19DyOnHmZGKYUVBdDMYJdqyHxG8bLPndljEl/wkZ
x1R3XDH4fZ5ooRxpfb3Z/Stj3j5bUznYIN+jcCxwKkagPC6UHnmGScVw19cKFmOLs25tywvE3Jqf
s58uzOTRHi8/SyVZ0zCZyBU4vr160SGr9ND2ljSeAyCKXS7dkWqOrTu11lSztbk4LMlwLXaNRLdo
QsFTC190xpJvksUzBCSV6m7eYjC29h9/fm1A/fDgIgZ8AcfgT12rXw5ZDJ1IBvUkvmXzeIdn0Ppb
arx3Q8wbusJdmL1X628nEKVQrXEesdDWC44PRhmhIl3Kd7Abtj0v7LEodkCZWh1V3llOTiW5yrZg
siXO1X8clzSOwUSrUDU/NyLWE0AXv5uzBXOvAQiGqoUsLRg574Af1ZjBjEk+M3dzow4c7XzO9S1m
4P8U/1lZzMWuO3Otaxz5dMhb5CZsD//TRtkNU0vagHbT8wx8p/Iktz/rdPRkBOePoD5UQU6R56xA
D3CxKAbQ9+3l7xqJALQJpiCoDHfGw+EIG3c4N2/3IyGFpo6FvhSZ/2/CaVh3JzjxDsCUTK/b0H2g
w8Sm9zqUcso4TfJRkmD9baab63c9VSwSm7ln35o/Cd55ETtLyysalF+4PF45Ly/uAkW8K6AfhqFg
PhVH6TQwdSLSggC8UDG2TlLCEqzdBI+wI35XH3FMnYuuEBxGkatusffolGDStlwlN8VJZmE18X5L
8WcWCWjuvunV2ukYo/uxq5JrPpPrmV1xToWqocSRWSrCWuTyT5IYHPWRDfUkaUO2N8kRaASthfE9
nHMHFU5g7tKFXlEMGViAxv9w2TD2L/F2K24g2nofrJmZpO7edJ26hn5DJLIOgxRvz9Hs+2zMAavo
Qr2q84mpCpKfq2bqKUPVosamyJUZlN9BEJi3q1kC3F6pxXeG+w/O9mPjXcw73NUaVc8TokAyck0H
26TldAIWtRxJ3pvVd0+FziWxznJCBvnR1XjUOwQJsvifhChSDVc3+hqZmoLQXk5b0duep1uE/bCo
v54Bi8K2VVyLPOmbpgB4B6EtfzlzkzG5O9rUuKmh8TUXlTlw0PmTbCfnwDv6qwO6i3GMMhCmmKX/
w4wCI+gBqtre4gHvcIi5VS8QP/Q7rOFBX+yjBTALOLpYqLckyc9K0yEiR91cOt+p2Q3YaTI1+p6k
ryGEfoHuyWjYIBlwicuEZbOc6nLv76JfDl/9zCygCdasjcuIxTJ9f91lHjm8OF/PQ8mb4GuWz8wR
w9wIFmPhyhlSl5TGJUBcOXszMflM5jkWcPdGRTiwFMJzkX6dWzB9vqeMfDvZD+HDhp3yGCHKF/Fu
aVFmopnszvnSVZw9C9UUUBLt+FwkGF352PXEex2FLUx+bUClcK1f4IBcUrIks55reu5c8mT3qHjY
tHrrVRKwlHrUD1xBSE7OE4JNR1lEQhwVsRbqkQGSSY7DIjINbCP7PQZvSfVerRnjJA+sysh5cT5G
a7mqnbMJX7XjTWgbryMpr86VtaJ5ND0YWYNTYVXJsWj0s4zfegXWnHXjsyDkAVSFaMnCZkOO412y
+l4+13LbuhTp4HeEOINWMxStzpN+EUaRq6rb+9hBbXUIyFu72fSNGWNWWGq0n1fBcOxkwWTsDEAh
MxPRQixF+xlosLB9MIt+rIdI6+DoHGn8DWJJllh3wgfDTvooL/fArcocJ90F6sdFCCY/eQgAuVnV
3swGW0I7CL6DVoseKF5mLUphaJE7M686gjV60oyso2oeqzY3ZwfUJGXkQiIdb/GyPprhBwUemHWt
3CNpVv9U8i4LIE/ff5pYKGv9dMX23UNUtL33if7YZ14p2o6mN98m9vfqY15LI5jWysSbqmElixq0
dcjF8Dr81a7C2lRErQVw5TBjvT6oucNKs9SFXRKmbbaFaXR7uGIGeTNXRiIhWs205DF9KT2qiPrG
TneCvpv6u12sajU0O7IH5aZF1xFm9X7mzIH8mvEJZ7sfBXo4zWoXEKCDbSCQyM6GRqodJUZY2Jwe
EWudPujpjtANQd78dm0uabkrVRVw1CkpMsg7LfURLFddJnMH9y+NYTrEQtVOQZhn209fqN4IOxZT
Zq3YCoIZIDUy2n0+23eaTy2RhL9I4zMKLvNq2+446GLswicjBs6+bUHA+GyGa2Lyp6yvowk+Pp4o
H7baoCj1qSiTA6DqS00XGZ4IFX4E8RgMWqxcnMKD7ksb8IbcedVmEatVlPc8OmeIh2oTZc7gDP+S
ZzMjFfMwV41ysggoid/e8KbMmLceq8LJwhKpqgZduwszw7Cz8Y8RBcksDG2ZUreogIgyimtW9/4M
XqWVHqH8Qx6QvnCKHQRwc+euj1tiJsdgg2Y+tMdO199UjRBaPyMsWXxTW+tX154gLZrOtnHn0qRV
c5bNXZKWEmRVeEQPJOtM+k7C12H1GyL8PYdpJe+TN10EAXTQc9gaiuIMxyHuasgGkc48kTtX6ZPn
MJsZ3w6sJL3oMwEt70x7syJ2ckiBcoWps52OP3Q0HIrn4lAqLqVyGycUf1Jo7mLr6GXOK3HvODPX
PFCkiw5zoeKbD+3i2Y38iYF2ZisUX0CqINe0o6JM6y5/irc04fi8I+tONlGAVjtu2X1A0o54c15d
7NGZz2ZIruNHfPMUBvxZlej98g95xsrySs+Oo7rrxEOkPzQH5VZ6iuRcIf3QzFWh4YNE9QetuAs5
bsV0cPmiBhyRuYMPpi8WThu+LVt43ISOYxW5/Fo7sqZQBS2p71kQQFl0rjrX8vBJ/80eV6tUsuIB
RMhyqndMFGMbmcCYFGD1yiNz7vbcLgJuwmtGiXzpzxh5jJoKi76yFttbNidibMcoKuX8YE9YbvVI
wVVqs3k5OQEqD9V4DPNhkuiZkUPeoxHCU5AiRPK1OiWFtfMcanxUX6VVmOSF+nte/kByP526QN+S
+FLa5x/uaCiMPXZgfE7RZ/nJGqCCzz4ChfEW/ucP1FTSWpuCRSRLHZ6Rn9voArXhXnL0KmbW+FBr
jW2Fp/ZsoODAGGmxhhiu9js0uc73wbGN0amJM++qD9BahLkja0TayorC+I7vDVNFxyR6bNvhd7ve
pxT1MK5Nr6v1XhefUSrRhXrX2LGeCcBxbGKGZ3zs0QZhi7+Ot2uxgOvTECjIVH3vpG3x5K8hQqlj
gTA6NzwCdmq4DOoVzo2GIREpLEhAQkIviCsXn3Y0GKZd4r+Tq34no61oc8LwS/FTwW05VkZe9vOf
rb5bLv4NoHHA/76nLnSS3+Hjtg1r3h+H79/hIdxxViFBz5/BGm0ypz6pNQB411nNsNBcDLHyXyoz
1pSz3Rmb9DMWWJ6Hfu6Aw+HPMeAEfdAcWgWcFmfZzQjcucTrSrPzTGYGYW2ODcQL435LEG3BjnzD
JrNN+fzyrvKiu8ZkvWDOrpyxXBl2v0mITWXpq62EPdTv4TGX+z7m/9QlXqoT2tg6S6PLgGodz3UD
pkaB3Qme4B1lw9nIBELrk1Rwn7hdHohsP233BAvKnroJJlW/lenHB6ZhjrQf6E7Jk69h6ZddojJu
GBDlSKo7o9A6P2zk59Nz0kNwy7kEZfbyDpUyk/4Fa/rT39ZPvSG9+CQwox329pzZiJNWy4NAlCKW
8fgme62UdlC6ygSbfw2Txhde75R7/IgMJlLRjGbXRtqqOoS8W2loHDzxM9txx2rwfMEUHo1MEuQ/
1zCxmBtn+0Xv6Mhmw/VbzrfIADrVmIJ6U58wwhdZNpXKUIhefuyDWF1lcO11Z+xSBjng0iBdxIZr
/6H+pv/jcLe1zAe01MSBskLfA1M4Gjq5qxiVKW9PWUE9LCc/e64uag9+lxQi8+mMsHLC1gRlzUYE
wpUOtZFMP6Kkte4VGCFworX6+frhhIBmKNzRuGILxkU1SgZvPQeFtpMPOQRhuuzxBm8lWcBe9oe4
LaNCy8c9Y+vIpqTy4IKAE2B/f4mCNaoDgSIyPYhr5Ohia6Jt/J2zVxRT9QiYoXvGG54Qkq9PMoRw
o9RzMYFNGt3PzJYOAF8Ba6y3FhlTMT1aHQtQ+7A3OiyoEX/wsJhygT8jr2QxjVPu9RD7Sj1AxLlQ
BgqJv7VV/Z5T5XLBeZPKW0KPFpjMFZNsOmgM7UBevFxQzZ5y8WvCUnraeIhovBrzSqiQY7oTMI8B
IsG7Yjm6YyzNG5K+RhOzRwlMNkOizdITFujgzhgKxz2AlqrO6qPW6j0j5/I4co6hLj5nlUtOtlcF
Hg4QNSPnzYgbi3jBRGrq5DklVfTPQZe/KfwcH7RyhnJrKR3P92Uyq+rxR/EetGkh4sRo+oH3HNnc
xbxpZK/8JlDlBGFmXJ+rBZUNPSz8RzG3X7UgXfiWTT5H9jTkt5IALg9IsQxa2wPckSev5WsgNlrG
fL63ljryQwOV/eq/pqm3Gz47a3VphTkOSq3Tdd5YiHGJgOkuJhl6XoFDKXlzYPepbL8bP+7jRKNP
BeoqcWHXVewUqztq4swJr5GL6gkCauAwAGgOL0Gn2+ZrWdji3/bDK/o8cjawomCfUXsBX6M4Gxw+
3zHQjBQzc29hGJX9vr3GXHTEPGYNWzqpYA1lOC7VFqKno6K09AqyBxODehvAUN5PIs4vd8FAGUln
crFdHUmkrcn3BXYtgelJsULG1OM0hj4G3ZdT0e/J8TeKKUcFlbWoot2Ly5nyJlvB8Edr1d+CE+qv
22lkHhdq1QZIgZkv8zvnaCob+RvcCZEtuBLIQ/pjxwbKvkcQXiuIHU+YHLH/y7Kg0KePXgx8T9jM
SC2jn8nm0ix178E/5pIXJrpEi4sze4qzW+WMnXqAUcS0qzmTByJA6rQsfKtpjjvTU4PdxjcOUAI0
sd6tVe+Kt/LI7ijhBLkC4MPZqxpQ5DPf4hdBOWexOZu3Lzj+yP45srvQWsnoHUR1cwSZP09s/TO5
iou6EezhGgzFD5Ky/u+eMclZaRKKtSDA3RQr3+h1fuGcdzleHOQJhzwxsDQKhYjc16eeI9ESOEIN
nH4pIZwIBREhavlSgZSIUQhLWC3iPmh/BA4aDwlPQ/uhA5GBinwryQXqcH7wCjeledCEzng2igxi
tjPuzaQ2u1FShiojJia/YWBz5zogMzZ9yyU/nAurz9XxzLuzjmx0u6gJC2h6T6sFN+YOhTCRheeC
c9VjPmeirTnZeRJ8Qtfy5mY1//ORrN2XTslfrZbx6B6KzT64yGjMuD9OWVfoSJ3/5H0TQvhBByAF
K/czOgP7NitY4YmZtE3X0GaMke1t5E1FgbiKkz5sFgUzjKgIn/mH/0yybVIYhOtW1Y0za1sJRm/Z
0uoHkrGJYUroI4U+NmDgqRvHaWI4q24lj5CFPDxlpYLriimtG3txm5c3oxZ6fdJvG+CJxnNo6mjx
9pwGBPPinRAMeVBmwV1v6z1Tz78WCdUu8emH5A7Fa7zTroNknbNnNhTKV9qy+ASvcJWlysAoij5C
5cxCcG/tohobVG7i9JFLD9elLltkOksu6RO0umeCGbyiVhDWHHww/B5SIH+WzxiqyZEUGljJg3mz
9EHkudySLzetGgSq1tBGWewqk81suDhUGdsB/99U5vUweWaWojVXxsqka18tBT3Z5Zh4W9WgCB0R
fMZZRg/xCpyLfF00tReJvcaubWOocxjFIa3CqCn6J4XOCYaRCgL7CdR7LFqk21lDjfpbFoxgKZeT
43twEZccQefWBI/QFg32oa6HM6f8UqPFOxHP0R2BdrT10VOzQmqxrpaObmnQVJ5eUCfMGnIg3pgo
GsbEty40e2RX1xHpZ5SF0cLDe2k51psXUlHdKWnBxyHvakCYKUm5Gws6US9Gf4ye4SgIcxXbDG9A
tVqovHQh3Jizrl0g8NAPqxd3eY8bH77o9vgE4kV4dIMTvsPb/5LsDq1t3DbWi5YgqSzsuMpML78N
9xQl3UtpOlvsP68q9a5b2w6ifW8C1TS3H8qR7LwejDMwzCEL19pNR20JumxkAxjTnkqrdpvEFilP
wCRltLVYvjmAN8C2D2pyHEI4Wml3Tg49itI2CRwVFGdOu6vH7Ogl6PCh3IZZhFGw2c3gZ3zdDVzP
51Y2HHfM9bElwWMYVxo7edilJzkBKitqNVepLjEdgQQrBucXwamsHFxh4D65uSFkvviXQDgYC6Q3
1Hh662OUzqDNZKfy0OmAgWP1spEVPMKOITHN9tUGWXW3sfej33YR3jlt3mvi7S9EUBeEBQqS1r8h
4ZEeD2M6XHF2cfgkqbMsaQrMvn+TBYWfEpt0fjdFPqsVwc8ij47s9OhzJkOHBjQb/HzNtZIcr7Yp
XxqRbq9i3b5A0vO33sDV2ghIW8gq7VXJvI3PKYKUnAXCmQYYo7Ndy+03zU69D74fFgF4hs0M65/n
XqJpFB+r5WsMm4OcSgREbm7m6Hi6t9WeuEvt9h3vVGdj3MBggixcBccpk1xQGB6mEaedgbyinI/R
UYOQ3DS3hE7EAgZBOc5mJ7hkFrDRm1mitYgyZdGbOpTvRALJtRsPC/kFe94T8/rOvtBDaW10Oo48
1iKyx5Kq4Nrk+azZ2jCPptoSPvl8X7vLw/lQaE1fUIubo7KbUWlJoZAk+9PPCvkz83LLb13MEt6l
UZI/aaBh5HZXFBNfASV4I1yX4KNWHDjs/b5NPZ2sqKH7fNfcHd33YocFVJbq8ytaxUgLyCPIw+fh
ajWwDn4MjrtSccsgH4QTt/wDvVq/n4BcNuNqwBalTlfG0fZzAfa8+Fxw9L6ScdmcC6XSiKQPRnxL
fTDIvh+kF/jugXJB5a8FKhQBfieTG9qaih6Xake3P6g+glTCYe2QQV3qMk+nqf/cMx6I2V47tLSp
U1+SL8YjjPcN/8Y6ir0kGORWiFzMgfKSR/OiDqeF8TJzozSyevsRh2nfy85HnCs5bAAYMmiJevye
iEhuVP+yOGgbU891eo48VCmCfqdwxgx3aN4qgM7QZn51YPw1l/6ULrh/3vQhqH+STc/sWF9Jqm2b
9hATQ+2CUW9TgHM/yaQqp7Pwrzn8ryhC1kgLEz5xhZ8xnNJDAKVyyTR/EDyyFBi+i8CJROo2gFSB
CEWhabPpXxpjFVmAWrgxDYJbEYfsepIhKocEsH35DtT/JEbOlS5InLDpciKi6hFA7OBiM/tStpwo
exIhhm42CceH1bXC8sf/MghsBJFJ3XI2BuJXXYuRx7N6OrQItLGWqpWcI5Zuu31tJIDGGmG/1+nm
SwJxW4fvHDv5Qb+GCdWsMlvqP+HQKVAdnOPY1n7nQKfcIGG6f8sQjZ0ORT6LJvYNqNzUMC9jjuU9
CMFZA47LvySSsoXr5JDD8chDHezjfgoYQsknZ2uTnLHShv1eQmOfYv0xWUYdb6xf060Tazk0a+9v
ppvRClORnXseVwhAkqOZYgEBx7QkGl7woIkqAPwchA4AVdK5XK8CZyijkxat7vc0lf6HGKoNBMm4
Ozgsq45/CDKc/vdTkZ+4IULutMQexj4cWgaAMPI+w5xl7sN/3c6v7YYDmelpShy+jRabg2Ncka11
PPUH7ixu9/UENnrVBg1IVqdnsm2bUt9Z/AptYXWYVrTwpk7PuBmT07BhovGo0NENAIvTAotypvxO
jmVghotTzHLfAMI2KH/XlqXTVsUV8YDQGgYRFcp05ati21XVHptKqq+r7R9FgmFA3um9WvDc2dAf
enQ8qKH/ClKkIgFBvCtfsvwPD3rLrA5J5Pq/1BROueN8tNPqKUJXDcZddtbPp7M5j/+k0Va+hpsN
RWzYUpblbQjmfOR17WMncV2i8CBjE4piFwVMqQbeCjmU94c4n7kUuR6T6/NUSVxWC0CFUf7H5ZAp
W1sNwarvbNlXodmbnjpQrArCalEZXfnCzCEd6yd+SPthMAKoP557vsewABvVd/25k+pDsA3sSRPo
w0JdN1YUN8OWw/stBz7yDxTwZCHKCgGUbcQ1V8QrVWbN+HnbsITp62PYO7es4ra+N26r8MczhBNG
XgVfIxXvU4Tpv5Bwqhu8JmBLKyh6ULVz2ru9GoebPuZ6IUs8F3LgIDMzPv042tRNnCPAcrhMJvI0
5+I+a5uMjm9g+A7/aLgbKphbLbi3iWjpivLHdlI8QKvQJoIhkP+SZS22tUSi9UzSDBp0lVbQLjFS
w+VBv/AzCxmSDOftUSiNcp7/pcs1hdlxUh/n1fkKruuQ1zb7RnsNaW40QPd1cqULrlAfXOerP0h8
P/t7QM4IHEDYcDG3oPZ0WXSmN53V7Cj3DSSQtF0raUCSOKfX+3co6Z55vMipwr/3CHa/iAXHdBpn
5FqZfZARdUPT/+j/FrraUZ0k7gEyiR727ICEAcQ1xe6cful7kXQuz0GTtO1RrMnhw0hQndu4TTps
vSnEm+WsZaG8DDk8kuP2IoxFaS6d37ka08aVm1JV0Kpy8J1fE/cJCU3jyT/+z5jKFAJlj6tPTNDc
I47TpFjE5hJXXsvhrkT6NFhtP3+bft1fCl3mxIlN3G1fOdbaElKYSahDyzuu1O4dGIZ3kn5M9EAT
9xm6ZovZIw9w0O2PaW7U2i+rOZoevFrlP1u3PD2QLvLr5QMsyWkwWFnRqisKZ4LSadDH7KDEQ6BG
zeclMc8NwuJybrY92N7qWd2YfJXgoHFtZUYR97FaKnZ+HRcQnMmTE1hoM18U2QIgyEmJqeo9ko/6
GYqbHfLCF6HQ9tjJwqs8IpgPNWq6NZ7XuP+U/dhfusUXDWaVjThPVFnlnq/aI3CT92NHGyaiZTMr
DMu3i+kys/DbJ0cQhwFvDJxXpx/bI3K1OCVuhGXHaveC6o/SyxxUJWmijc+WMZzebZc1R6o3+HcQ
HpkjBbHM1/kW/JvjuCphysI6pWUye+POE9Q9Ebv0jIjRenRKxlWjU4/5Iv369jNxgZ5NoU7M0sBw
EXUcAc4jxW5s1aK+nQ6ZOKZ784yvHe9eRDKNHU+6EnAiQKX60f28dzb7cqfo3W+8BWBWwnZ+f6q3
9BsiVifwxYiKHTfhyHlN0LTkl7UyzVyTnyscZCg1d6Tb21G1sUDLZzeJ06vbfdBolNGZLi0YibvM
aOU0ES1P/nNNo3cE+7SzO6Is63tKYCuN6SJi4DZ++25XneLeCjEbkz2mnZMELVmVAdqH80q/QEbw
WVpWucxGjcTEaF5hfaR1xxTuz2hpFwtPOTLPkxEmdBIgeN4IkVUeQgTgB+Uw5s382T8aLwfQ6hYH
pik2YpsvlXyzLc21eFxJ33bo67dlcFJd3V0KnYB9lEpEVJG8CFLqo7UYbb1wQNVJt7GBDvpCl7fz
/34duq1a8f8S9jovA07WiipqnJiG+VSQzjdUvAR4ls5NznKCrolkgwUXpY1o6JegH7Fdqm5/6hRh
WiYJQAYTET/Yug7zgWOXXZluE9x59TKCMgIqGNhLveVRTJYPm1BpiqRQ5XPFf4+5iMtleqIrTQfe
jumjaPDRpP8FoO37dbD9V+XkiEWb8vgyOUXy3OffrIriIjpyGkqZ6LGQwjIas0/z1s+N+xn9JMAY
WtgiuoBX8GTIgNHmqRc2BsO/ae73PI6MmRR/Oy01MRCWDlA0Jm+yOpXedIFLdZymK+k55Ci7RC0V
RJjXsEuqfhZwuBs+nXacUMq8CV5bbL9/sxbAcuZ6SOZGBhfSI9x8/mRf76zVOKQT2keEcEhNpx8v
Zf6pvnNkEa5hbzBEImaqbKjX084r2/UzX0S6SrFjlosjHv+L+6pknwtHOzo4vXxLMG1yL0qM5R/u
/xyQP1xMpivteP2pLhsbpfbfPjVgPwccITNdStj6zC8tCtglfQUod0Dqw848XGw8yEV3RwAYkHOt
Q8qBfQRVqEhnclTarVzq2T5qJWIYoK+V8oJWPxxfnbjgxtfwffq5R0XTH2kXlAj5Z93hHTPE0qSh
iCH7XJe6YD0xyXhXSrZSRwBU5N3NpKNUC9h0Tak2Mkq8f8acO04d1BVTAYOKTJ70jUNOorH+MXk+
yxHJ/moV/EusoodBLIH+DFlUVfasvQsFB1P7dD+ir7EPocZzgCadE0YLhGGCrf/c2IIcPS9CAlZA
4b9uqbkRfAQcG82C9qK7CVOGvn2RNrEV0Oa5m+ds7Xo9uuNmRvkK/5qlbGTvSjP4d5nvyEv/EULB
EFfQXW/zoV78KJX3oB2oS4gswLxLZv57peFTmvdvAP56AOB9GLL1nMXegGJgUs5dAPfZ5C0xF+XN
JSUIJkWn/HueNkui9FG7HHuzCyCu1l2pPgFFdEN+zMCJ3YF3KfoOKB5hG7QtGjfbF4Xj22gf1TeG
5SqwE4fEozeBPcK/y5AXA4wycXoKDRMU5wZTcVl2QL2ALz7EF/FtCAIG+YzWyRdqpWkLMVENUykL
OFoexbwlUvoVnY4FVIDlIlctbXVAaA+Tu59Xnfbpqb0OV/zBHKOX2vydc60L1IRgsrJ8E54PNYcd
s4hbBXqAzUXyVpe0uKt9uQeJZLA4zLmEQcDVvh0vTY/SNRnuaC7el8+h0W7od+f3fl6SEjHneFgy
dBpB6ERFKRcNpoEcG8Tp32CFCXJlDiSbLMFUCRevnQYeSpiwWe/6oaPE0ZYm0JGoX29BIBV0gVoL
N7buH5pCPlAU9A8o3b1gJChhUp/ksDCPcq6NFIzuDrdpleX5B9+by3PVDT6oI16Pq0nGrD0SMYaC
y9Olt9UnbcUHUgkUVPHDR72kYy66RcUT100QYTpZvLgS5cDFTY1hvEAQoUdWrZ9SyssNzF7vRF1A
fwZ7HvTDFz5fGRKgLEFHoVhOh3Q7mbY59GahMsUxoJDBg+iDoLbu4gEaHbHlFe7jmgeV1Xo1NeE1
LL/QzrO8672uko55pruQSXIHnbppkLWNEGJsXldj8cWQNqhoAnibmTElaAdynZ2p4F8NKCEJLFJg
w/jPJHC8/6pzb8spbZTqzjW6l0tQGRaA3JFxPlibRKDx3HuGKR20OS07Nmojp00MZ8QGd84r1mLA
LDu16zFmoEaF4KGmXJt2wxylu9t9EO/ksZSRYmRxSO1Un+LVoBw+Tc5hPkOKmfPbQDN5dPgE/q9T
gD1uhEMGVqXMh6kHk2lB9vHrB91LX8YDlnLn6yP4KjI1tYR2p+McnhIf+sFAfBg1f4JK8t9lNacJ
vLTY2DYssZuoCd3sAUlEdeTfT+fByOxSlVl515mc+JbO+xDbJ/NapebzyqqT78sYzOxivQVIWruT
vi4VSyJe6cjjqSO1IHU5ffBNmgJyo8FhoC7RcpjtKc7B60usCJmD/PHEc9lSFN7WmYKJtyFil2Az
W86uD+Idv4TcJdGChwpIouXZ1zoHFOJvSclOBaCHcC6xxcqOaN0j0f/r6KOUCg1q/zWPttqD7WaE
sUSZUxSnr4UoutpJOBaZ3yoTJ/6KN2yoDaCkT+8kchmkF1rGX2FVOhddUjrzDxLpMMvBZ1cUrHUy
wdH3VSmvjZdv+ZwVck4PVQ6qYYKZ+2z17nXcDtPkC+i33yCCIt+9qlXUrf6oFH0RLewCWkT0jA30
ZXjpqItcZFS9ruzOYi8v9jpxjsI7vRFsGIvEMUtkXFOQzYXDJ6g9VCsPYkn1I7GN233YH6FzMBzx
tkV78if+aUvmasEaory+GHVwuOdevL43PZDcglhODkhC+levSq5nLra5fAyuDkmJuNgO8IlBMqJD
hg8rEmWp/oWH0bOzRyyN9aJOMRraZD1CN5HIgygWdp0iiXLdSuLpStVtPMjO4TObDBitON7Ulr3Z
lwejAtfbY4rHMWey+Jwj+gouWdSHjMDKCNgvKxUeRHlUhx1HanCsVIPQKCsyjBeTzueYGPDbCHQr
AddqNq0M0s3ZNpbNJvBZ+EDLP3HquagUUt2FafRvDhaBxGY2NFGbeC7xLWvyUrwmP1fgZtVkxSKL
QpSOjfVkSdO07quDvj+65rziHyayGjMgTl1O88/ewvb63jImyNAGiujS3hKFoQGdauWzSVhQDHMf
Kbt9sbcHe09ddyQgT838TDTpiPiGmw0J/ObI7kTQOafNv+LEdpWg2V4kfPJaI8VmTSGLbRInSsrV
MuvTIoXBoPyqVSZdwoYTPgHneQIa1FVogrhmz+4q6nlipSEl+AnGu4xmgdci0VH+N5Nlrij/HCKc
/DssDIhux3exjTITgwnuTv1IUMYTCKpx3mkec29N0Kj7ywA8HTTvu9qZeZZrBFfPLdw6f3hZErUV
zKBN70qqumSFm4dpn/yFlVflk9jCUcA2OScESy86JYSWkEeIEz8bNfrNxGRjGN8I8dm1BY+YKDGi
d9zZUVeCmjgU/8YHUmPdD3mlujQ0nMmZ6axOWVI3OiVhk5IG+7YQh0wQXCheeTzn0utu8f57dNR5
3BqDjeY3hQ/FU1eRgIUKwy1vFTlrvxSCjGxZ6bYLNWtaMF5s7utwI4oxJrXYZfZ1Q7xwXFijYteW
t3c4OzD5ZJTuu5JtgnwQ1LVe9b/ZCAigX5iFn7UdPzGs/EwfG+8bQNbfJAE2HWE8r8zKxK6F6Rlw
pbDZxbBh8AXOI4BjDaNwPSiz9+QAO9frAr3/jkkVdg6EdAiZZxWwH5ezN8Kc6g/z2Ywqod7qXYvh
P+cx6LLpW2QnfZXkpr79jUs/3l8fWUj4SjkTd5DsD4liAI5xW4vXkMjN916ziWkTstwjjOihHyqs
yiudPMIVufYnp/5G4YabRi3XEs20Dw09w8xfOFm7KA0t56nwtUYqt+DILoQ8sU7LrFyiSxLR/J5z
Q0+p5GoIiV11L8ERbFOkWY4oG6AKuBIyqLh+ZmSJFzJaMYl8qG7y3IxoHja4Ruq3SZoQJM9oPQMC
fZuCOWv2aceJF5C0ZrPRecKfryndfAPEr9CuQqzo9wyP5ofM7n2L32p0ejfwtk9i7FS0OMf4uJWY
MRTJp32XGhvZQDIVHij1BiZD8esc2v1fhYVQcy5iZNYlgR/70qdeZoafBdooyqaWEJx+hn6SCttZ
pVM3V4KbQGN99FDrnXb9Etq3it3FJxU0YanWVGXsfRqvOpxNNn6FfJcn8ocbVELeYK8m9cv0l/QI
22WfnaFfqDT57ja8kdEIaswvSrpYOyCFaX26XsNj11T9RkJU13C/FNJYmN7DVV/FlijUZdS/CLi5
OIAXJGzuPwVr9+A+k8S2c1Oqvded4MAMOHm/W6UaLz3Xc+/7MYr9s8lptHZhABzin7+EmtfF/1EE
980HWy1Yq14a9ccs+74G+7h2w121R0Q58knmgqVjUUlv96kketBNykprgQIotsNGZoRltSI+Dw61
0JDsw0tmjU5XeZaVgMN60dh2sKFuyeNsPvGbUDVAGc+VZ7kL1QNOjF5SZWdq0lwxVqrUHUoZ1qjK
40qhYWdIT/5n9ai8B+KyGCtW6PhnTEQQQu8W3OIGt6M3sM5H67eqOwtziMDXkn89tH0bJeRDOn35
4oPFLUkwWAWX274zUbDow+d/0y03mCh4wZ+JidEgob88e4emyWUggh8f/oXjoF+0yUOiO4pPCrIF
tvstwjD0+p2RW6thejKbKwb+HkcRp8vRdMR0FrUTlngeVR+fdP0cP61rg3FeWOzYscTqbAqXL2cD
TRZ6xU60hnAedlrEbjch8SFCQZntdbxZFMzT8PYGZuADyxfbb2FIZhIN7W8YU9BKbmmFqake79W7
Xg0btvNxQS9zpF2M3XMnIL6ucDqI/uSHrWPEh7b5yygSqTPz/8Gcih5wizsv1krlKpctqCg0HrD5
lXmdkTsUMy25iaWhrS1oOAl77aco+jWalNJp0V3deu5EBAM8oIDbyOPs7uvNwIdpsxefu1XhvYlr
kKbwGL/zJxQyrNbfQupSab3fzCT1tTwaMmOUT+NG3jLh5j3aQ0YjOpH+mP0Ymlf+yvoSVbAMNtcl
LrAJ+5MfTh4gP3afibq8AEpro7IoK5CA0kktjnHBlfhqBKafZXYrorFoQ5uSiX5su01VnG81l/lX
Yqt1Cl5wOsy/OqgfUO3O3sf2BUXCRuevGA0l7Nms1o+d4n8F/aiqtZz7RieZNysJu/B9RWEynUaM
HfN5Xcc5RHRj4hPhl3KAF5qgcCvu8hOfoXuCDy6/oouCgoz5TPj60H18dVpPHQi+oPmZ7TtocR9A
qXUNBiiAHH5vKlyJ0AKW6E+xWNLyo1SWnXGeSX/ksQwbg9miMtdwOjjGEZ/33BcCs7NhrRktMZlj
CtKDrX6ydo+0jtwqX0Bd/WteWh/OfnVY0VLsAoq7zBsTpjNg2bHOZ1t7uwjPdv/eJRR7YRQySza5
tJdM+S9CFxTcEr4S80jlKbfbgM6sTmEcES14aaF2m6pxlE7sSwMDtOLH8PPROb5gngkYXHLiHDLy
NO1iJpkicDqD4IFBz0/UkrS6iyF47VG10qkHutV6MQu/iwBLzh5hxF7tgHZr/VGMWpl8PpHIyNCz
5N+AveteLHNOHJDLZ37J4q8tLOsU7+6zFm0OAXoQnMnysrIDdtb9aVYkbo0mLUzm4nXvQenzwY57
TFDHdEsGX23F6Y5kg5AklvQcGY9GLyj1TbWTXbjpJRQW7GBuV3+24AQRd/RpyEQi12c4egSDAJqX
N6J3li53++q899tBFb3lGl3Rq+MYwfoD/3Lp5rMxgmLQrENGBEdw2c/quveT7C+5YQWy69IajokG
O8Yfeov4PpRv4hz9MQvjHRJD2Qq7YqHW0DFtWWSIjFR1TVaThnSPIfTLJGg6pBP9tYIdSJW6YYuB
GeZTtz9EAUCndVXrfVjw5x0l+htoPr5hphGD6Av3BA7ZAXpoiVJIbTVxDYUek+GeU0pZ5JmG1CFw
FdoGb9cGerbWuVGiq1W8z/in27oNiBE9SYx4quy/wMI3SktV5hN5cJ7woPOBnZYKz2wy4qcSWEYV
15Du54Mgo+Dkx6ZluG/GvEa6TFmZeoBIYsxRDvI9jTst3IEdBSPBn1rquWzQcmkjtQ2HAYJp9crR
ch6UsPRF3e9LJCLnHYSB8Qj1/HYqGe9C7GeNVNpI/jEjWvWqvGh16euccWn3jIG/1DMyHnuRvLiw
ND7Dm4E8+/B81G6keijCEuHMl6oZu2X1vVoGUA+6Va/aha4NV1ongG2YusZmtcyftL1/l0WtJZfl
tz/tmstHvnvjn7b3hLKsz5WDK7AJIlOZXkLgiQ0JFWDvqLbYfhXGsLjDG9BSsvjyccUD4Rvha3Zy
PfblYYxjOQj+JM4IzWD/x8EQLq0wr6kOwskdh4VFPUSL7MAmzXEXckIIhXHD7xZhhyaMERUngPq0
JlnGGrG16ERRXfYdrHHLJfDb15ArxOjNM1P90EWhYXG2SetmrPO+uL09Vc4DywxEtC1NO5YyZ1oh
EOfiopdvA84taLUFllCgdd2CgRXpeMUVE0BMsdWMt2hnvMSNfcdke53ibM0ytQY0T+x7JrmuQ6RG
JCO/X6E2OpkOi2PIRnYL8T8swxG2QmUboW1kvgCE54DZ4hE6+CvQ5zHizJytNIb8KxLvAfD7eQ01
M/BtwwsyB1Bc0IH0Kk+QXNDOyhCik40zMahf+K2kYmjmm9Rykn7t5oPaB3yoE8jE5d13AMs6dndx
1n+8Dq1hB/VAFj0BqkSYQCXYq0NkkCd60UAfCZoGmGcT8rCKxrgqZUEInwB2JE/LO2w3dp7Z2kMJ
YS65WVcViVZjy6ykpfDAH+baxnk56zMViX1w9xRoEAyiPVf5i37s6MLUh7lg8+C2Nx3pY/wxG8cP
WhvOdwONEASNTscxGLCTCTgHuvBAk1eTI8JAjVhwrecqrKyxG+TfIoAsB+Cc2RjXpywtKsOUGcL7
bttvtBIIlbo4vuArr5RwEwz4gL0eg9Qndi0fE3p/W9k/nSVr/5x9+X8Gg0PbXHe3XdWQ/zsOLSWy
BnbCvbyDP7b6L0Bo9/AiE8aJTDcX30fviq4w+wq57Vm1I74o92m87qx7LEM+8JJSDpqsquvVmuMN
hn0+hRDYFDYz0WFW0IC/4R2E8feY1PND67TKTyWckldNUr6+jBuusW+WphtucoTcNOAoYCFoDqAT
UcszW0qI9ukaUvvxRm2GAZYgpOytUHPDYtOKtvQsb8TlOWl1gEXTddxV56ti1wXVnVSVbFmShaWs
ErPe642wK6Ihe1wXaaQC8wB+M4wSH/ERRxy5HI2F96EIKYCivmp4ljiOH3l07REVku8XdQlOiwas
aHZ+5LUVujORFPbxP9TRh/B6Hhei9dtICkusNukjZm630/IIoqQkahbmViUnU3P/7JllcZ+4sD0D
2O/Br4rQWm3uiOBXfoZ9d8kRUYvrQ4dna1V6l44Hi0JkNAqON7Rjwo+FIXAVQQa/sC3nol4OvR/p
/c3vxThG7fonMMiGW7QKW9ql7QXZTYIsuzIknxOSW5H7qiHoUXUyqqwefzVNhH7hlF16+V+fPOKj
KhJsAPGfEJL184GF6hiD+1YxuGAerdKPlxmg1LmnGX/zuxnD5fXT5ZwjledrHmzMTvLdEuy2Lgp4
6I7K2aAxvF6A8YwcSmJKtSWLjafesekoL59WYm+lo7yIkS/zOx+BL/SrR5fuT4oe0FIyM4Vk9ZTh
0aduTxMC1AVekoRgwo7muYklJo2Voff7GfzJJcovmdSSK2RqxKvnkHHZAQi07pCLzi/5/qgikNDC
jsDM0x10Z+AlzLXKlsWfkGE65UQdRjRzfWateryfHAqZVA7hQEyvPOe3g7Fbyiscw/vZizSDnMSp
qhrATFGWOD+O9wAjlVWK6VQIavoIDFqXXoM+cHTmSW2Sl/YB69W1qnpsjHjXYNZN7cMhYMV4bf9R
G8pYxSPBDMsWZTKhERCsdDVlVQpBwa2zdadxP4vRDngcesn6bSZrLC7hrdRUa/pZULhQf5JHP34f
ATNExOwwqieO/gy4Ywo5DkYseTwCwftN+Z9MKFjw5jwKpbQSeResi2k+atosL5XA+PUJdpngxsux
tiJ6O5rDo2A0k71+k379SSoPMZ8+6gyopQUfkCdl1JRoDqvHSrSmYec+bSSmsR4eu3r/ttyesyPQ
llKljpFZTzJy6KU/XLS0vjRoHHGsQ+cSFpxOLSCRY7C2lR4nP3dIIIJJqSI2w8AnNTiA8O7g7V+s
FM43kY8eYwkBmRCmmdlKcq4mLBSxKJvhkY2v7su7X8LsSFl9FMvtomhpx9jr9m3HZGh9xHAlBtUO
Yg07hbPn5erQztuuHsyJibuujWKCC1EmwrdAyGVDoSJjfDaTRzesUAC2yeyCcVNA9W3luhuxsvep
Zm/1dODgxaWHLKIerINs80EyWxpc+yKZCoxuATpbyLIkb+jmay7lKsN3qDkfUAPMyZw+M7PAa/jc
cSsOX4K4EnL1d/KJf0GyllUF0khKeCN9u8By42NbCm0eeqGpSevDBL9rsBxcMSAQUSJiO+4sqF7N
o30xEoJo+yb8k4Iwoh078zl9vZLsq2x8Wv4NtPDACgsUvUiXvtzk2PkPwAuNXWKByKDXe+/nJqkX
6xk6uKLJp1z+w/1xk/zaQ5rRnkC7B3jorVf/nZPHk6GoF1rASBCfvAH+RkCA7C7K2yjn1in+KhyH
pXknRLmEnCBm8c4km/NIwUbUvXGcf091jCp59WCyFOLg/mDC4gZIicIyje/V5OhS8B8CoJ0uFKqQ
c7Osu6hgXqvicwRexQPIPevfWQJwNcNl2pLjlcQacmcU7vYPiHThWQlHHZ/11yT8GBNiSdV4JB/o
+yyDRaNLvgLPeD7sH8yz/pK+Jmdi37QDn62SjJ4+bZFIn29OR6eA0PjP0uCrvQOs3UypXcwu1R3n
4Fy2d/lQIhib74dOxRnqnfCEFNkNpMvHiS5prrahV88k+X7oXv9MerEKV+oFXRnQmoi3g1Mq97eT
Nq6gARj7LU7kwQOlXkVfpIFYK8bZ9THO1R8FSz348CIsl9kJXfzKm3GCa0cPkO6e2BgGrqU+U2Cs
vmSsin2ZwlzQV9m5vAufXOhCWd5364Xb1TVyvCqIdrJg+6m5zygktfp2CQY0ppOTPlRCMsww1MkS
SbNnCE8Co3In2NpPh9oeSQq+EiTr23DkhV3lIXngULEjzOnbDD9mERIbR+xB0v+iWgig53jXartP
+b4NTo1h6O8k+hXxqicPvAw9jv1dNAoqpuBUDnhJi2R+sOsmjvxMP4Nb8XPLJy03mYOgU4WB8v02
pBXlCqCcz2fXfYBAQvmrWl8RMEOeMBgeArX++si7t7kzQj5nYhl5sWB/JUAKcjVkk8d3RrEmiBcx
eAGAtYvN7oR3ZLXMf//eIG8iOoWbSaXluaC5VTb+ofvKyz7kBI4J3HGxMw7ko+WHhbZ2ZQ22uFru
1XtC7yTpviUNqdpP9WCvhJWx5myQ/WrQUaSsbo2+ecq67hCkKMAYjbFF+SYQEdDWemN+5LJtHjB+
BIIstuqUqfXZAFkL25MT/FcXCYOAwKGJJqzkb5YOPzDspX0m88TfcWN46sJpOribPYDdH8ocq64r
RjtDYKj0EOsPbfiBCoMc9KZSmzIRx9xPIMacTCkIjBiC969qz/4GN1GhDf3JjPpVFTV6elqU0hbY
BPjUgY85lE0Rt/Dm0pq+IYNez2pbJr+CCYRAUTOMX4AMWhOVhqzwiiOp/TgXDQKqWDZJFblvdmTC
6iSaaj/IuuHqF4dHxFss2tMR9flVonhVYMf4Lp2ZM6EIOQ9Wi04em+xCcGlGF9bIId3iw07Lqsx3
DRSWbzBkl0RkLvr19dt1ObePzqipaYeoQuU3iVmok8OOTdytei5d7/ycRtC71iKqCrekh6eT4IW/
aoaDE6wMecR5fvqsZs8Iruc1JXlosq3+IV7KD6PWRTI7iLygbLLhwVKonSs1WY1IGnjZT0viiTjd
30ApkPipPqlXo3mlCSFv74B7kcplHHDkeM9EkLBJL5XAvezBDU6z4mYoTnjaVQP4kVWz16qS8B1Z
dhd0Fe4Ytp/1Np65akXybOF+kJkgVaMwQkwdyFqpCqFt94cOvF/fcXtxeOnMY592fINpQS+QI42g
oLaN3KCeuLTMTEsTCYDFhcwQ3iLs0CcEaVMV1lQUlx2YbnCok/VHm6LknWcjZqoO2yAmD30N6xiz
Zcb4415Hn1lG5W9M+0NEwGnt5Biho8s0gw3DYZsI5hbFaFFuS4NWD2ZQbaKW+MRgVsi5wWkcYGJc
TrhFbiLBm7iv8KmNG/t//1K2lFllbjOo+/wTcverU7Dax0zZpqWlj1nWknhoL6g8JoEtBgVnHGyI
h2KOCM/85OvEJjfgVAST6eGWWr+OBStqQr0SX3n4j/cZsHbUiCofJK08PLY7wzUX4FldrdDcqxrg
efkVVkO3F70MhgL4Dfr3ZRw/zA6/ooxb3xpOFzMGAfIAnq6W5Wv4dqqJMAQSzKhdgu4E9ncwHXa1
kJy+g5LYjM41VpzPyDQl9iFF2cgq30ua8r2kkVHq8OjAbrHOGcP1v+KSEVCpceeST0H++AE49Iuc
F51GPaEDBv9NUKXPcFotkHWwNr7s74ayjLwuzHQu0SKhvBpXS2ZpRcnbHNDez7a4CMJbzssiI2m4
fz0e+kVYSXff4pPd9+EXbVaHN7LL11YEIrAe8hNDWXi2WWb5U5uYztoeizivDXc6bpC029DCwm3h
9fyCxK7/znbjW80hxaV0f/Wh0Br/0F6Ps+c5iUxJ5hShrAOLBrwrgYE0Tt0hvgViDojut2222SkH
jwQ467t47fX4Bl8lp8Ipl4tTzqGbVi87/+Zkb5/KeW50syCqZYQAYZ95l4M8EdY/ETiNg6rCXQH5
ALbUfnWiLRE2d8AJMHchiyDFUIOOxeaw5PaNlNYbxtX0UU67v9Fi+rsL4tp36uU41/VLonJmvaHU
FpBDeKjkvanb+boo7Zn+PmlhXcyQxRMVnjAo1rD/hvF0wgrPl4uui2A7Y5f1cX5zc4bQ4tPTYD9b
ky+vp7mkRGx1HlqQj0YsbV3BhWK+t1QwLi13apb+T7FgvG6sXPc/caahKyfflj3+MwrOUdwo6yL8
DOCUqruXYeaDfseCNFq9Y94lX/Lqh0Ys2M3/QKPbqi1Zh50yOmnMioJdeNG4vqqZJbXyKbO6aHdf
WEyqOZ0LgYKuPOS/iANH7KydmbzZj0BsWFOVEDxX2JaBXP0R8Z63gekYWH8scSsiEUumLN5t66Uw
K66HZxbpMWHnBhUTnxM19LwJywsasplcwYAKh8txNYrlpMIxRL0Y7XfIYgmN399tYR70f1r3Xsl3
f3+UdDoK93l1P4d8+lfGtPlz6TtHVmNb/bfqMYg7o5YaD/JeNFH2PRW+8TCzM0uivOUH73NOSlIE
tSsAkZcF4TZSF3z0UZeNsc9x6FOxHlbb33kMDU2DCygeeZYlzxFrLQYCPUSGZqRZcrPP2ckIrFzT
k+23+zBUL/AGYKw3Asl8RQJxSfsVusZ1jhqnieEWt65Y8FZCV2vxqN/wy6D+34zSS0KI4XAuTwge
yt+UXRTxYagb6IpfGvs3qkNkpW3QhcOvVf4KkeUUyrepeAvJUSWl/04ZEW6iu4c3KZ7vVEpA1DgC
kIdBcx9WRQHHfKe27KVrxUdeqhsm75yRxRYm00AyvCithJ6ucoeblDUXB3mz6SbeMU++GCIbly6v
VQDRpI/4PAekp//jGBAciNzaX3rtV9hfGIZqlpzSCemeI3IBjMKFXn1bvhWZEa8Hi5CL9JdewO+7
tBdG1BdXScqaXOw/HM3iO5YUE3DfsXzx/uvsgqvQmyzxCE2ci6fF7F+6B/ABb0O09HgXKpPkDPk5
0ym6Ek8QUpDsRREtiO6ZcW9ky6jBl+T9e6XK1Yal7s7W5A022BWP6eL8O60jOy7I/5Ica2Z6cNKr
kUqv88f6kh39aHwJ6vAGReHx6Ve56xB7Z3SNZKVBxK3XXkeutdHYzu+Df9OjBiszZOv8pGlIXa2y
LVqxwsSdan77nGDB14zOmJJXv7mUi003cBp3PsLnYz7P2VsKzcGDxmOvrmdzSt6NmZDPL586pLHY
tGT0Oa8Icrlu5Z2sgFFy9QlYZ6xefV/cNXtd5VmsUi7YWbjFtTRW6cvoPiT/o/ixbfBd+MMWtQDm
o9diA+ZxKO/xK1Db3Db1hnTdc9oMwujQOPrIMFAgWlN2p3vtmKJ6+AVUoLGzAYAoQe4wNZjCO1P/
vyTdvgoO4rH7X+JTFYmw9DtFlVyH0O0Mk2ppfDOqCAOuKK+yf3kHfHhnGOrBHbF6arenJ6EqjphA
9+pSmNPNVxJqfxHr6N1Bop46/MIkAd91t9p8P0mvTWJxwgFQIy2wjuBkIjsyk7C8uhUezahtWx1S
KCE5Zy6eXdmMa4Q1o8JH/K1tgaL60DFrKhqAvvNL9ohFEH8wswPBhQ18iVbJcW+028JjGMuzkX7U
uNq9CcNTMqt0OgUhF2c28rjR4Lneo6bYelN7qdzz/ThW3cDEu0ZbI6mR744fdjydfS8Rhy3SKyN9
9abOV5Cjo1ydgDuG0/MNLdz5nGcQK30V9Xb0rRED4vayRKoo2N3pLkXfjQ3vPQrbqcGI2YJ624w1
YVgGS9/gbCv1uDNsNQ8vTS7vJclRO45QcXCCpEmqtqNK0vJmTtB+DsomYjB+uWlerLLVriDFK9IM
tup1NehijfJd7JvW8DUzT81ezKhvhgSip9BHWokbGDz4YbHTipsRbZJv+hwy6WhjNDbwDieZWTcg
KvfTZTjtRsxmG9wNU61EVMGi2SNcB+MotvddxEawDjM2+l21RJSivLs9tnHwVVW/FA4PNqr/2faq
V08rV6UK/nom0UGOEY0udyf6J+xA0S47orcW9JoX/Qz6wXzEMy0Buqh/9FDzwbWRviV0yzj/wx2B
llXF2rI0/pifTDknwx4OXKLmZuVDcjyxJwXcKkRGUoQ9xmacml+Gk+xMZj8UmaF4ySowfE8Xy8Yf
G93iRyL9FgONRM6Ich6bbS5YceKxBOVQ8F6gyJJPW/tryvA4j+IEPMPHqjYXfGKtSGUNvpIcxw8U
2arKpoUNW1lzMp+2bo/YnZAUthPMBoct7dDBn0Hm4SFvtqJx7JDZbe+REVMP1pievIoK8ZvzVRYZ
cRfx2OMixDNbsFqY2B3HrHbB1cPGz2REv55F3hHW9/xX3gxLtTsf1eOhGorfrgnHEFiGFm9MXC32
AnKiFd4HRgj4l2gLY5FggdCGp41zxpY2C8/lwIsM2tpLjYLu8CEg+E92I0VfTnGBdIKfemrtoNNJ
GusdM9przh0i8UhWwG6kzUqNNCi49/n6MNHjQU6t84AvkMbpJ0hbVidVJDUHmyW+uar81z7vPSOC
0YR/FHViXPoysGc/ONjVUdSdhhsNJPGq6MwjoktXm1HSjmoPSxPJNymxRzScm2DSn4/8N4uI+jyJ
jTsMKVSmktX+jyQAlnMJeS+hWmcb2Ka/xZysrjqcYvbhYmuCoGuqbhKYpfzMoD7F0Zh9RZSRgpUy
epKE3TXa48kJvJn1LhvZ1+KKGipMSW7aMyetvhIiD0aBHBak4RtWaWc/KYbcAvoj/0o9QfZ0SkPp
4U3WCPNZhcuD9RcDLG6o9Pp15cyYuUzhciGhB4yiVaprwMnsZ1vBEAymHC7MrDWw1A19aWegLCue
9XaBqjFQS35X1RvkzW0R9F+/Ely7qSuNEMV8lChn9IWekxOZYJ4yywVvPQqr6QitgUQ5b/v1kP5m
z0/VYi6CXToR7VEm9+QZoVy4IcKD/jw4n468RE8AnNrNLfZFa68S7wSDr1xh0cbCzVfFHOGNVfLw
byAlVOEtc+ChuODL0/pO7ICTj5J/WefUmcUni7C7JuFGbblLVgggoTsvPjED+PxfWoWVD2Zw+6xy
ArMPWWd6OfnYovGfh7mjp4qnmhQnaf7gN9bw/VlUVe4Yah19b5enoSvMOta0bwNtW7lFi2qy1zWH
ZloGf4cxckubzg3NCVJ7lU1H56nHN92bshi60On0M4apZauiVeOSwjG4/hycqbGyg3mhahtN5i4l
f7c36/YPbSR2mRaoQGUi7xkQzpi8ctef70Ew3Ef23XdwGhHQHJ74U9o3B4s9FXjbp1gf9JfJEhdD
vuAy57PtN6Q07cTat0vKq2tfrm2bT8Q8I3fw1/2xF9ZnP3rytOarU9YCSr/n9y/d9RcL/TJv8KU6
SPtPDPlL6GcPq6vI5FuzJCFJRkfyQ0MNsnxneUh5TEBNk2kBMlLpWL0sh+TjsNfVJb31BbV581+8
0lNH8yvNOh94eaU70XXwXw9Qc6rf3CAuMdzDySPsTwmMDXfQitxGNZV9M3IvrBOXhSTOv2C9Rqfo
cw3WQcDFvSX/GD2mx3wZh/0+jjgX/IDiwdrqu/UgMBMkSTxob0XgXXrQ5AGLcRamc2YqXqQ9mlpm
utt8Eg6nTVCLDgeHhwCZd6kxGv33WzkcCeoGTCADP7nlDkXfBETvmi0Jdpc+kToBL5haWVtANAlL
4gCuOU/a+0EGIm1vNU1TdUBQz2enGLjisSoO3J1oRkqrSIPeRHnDWimvkdZ2x2/yJ4vABVc0/lXy
qWMOhg04yTomXWEjCJUqvkw1iEWCFw3Ta/NKFvx6z6zfFJ+PQ8QNqiICtOHycXi9Ii/D6Rk0tC3D
h9BP0vmV06MWDPoIH+YGSWWOjZuJuUD8msCU6gj8CgV07dDHX3/r+H+F/yKHRMswJVoDUvAe1vdv
SAt7Dn56h5RwPutFlhs6GsQudto419Vnlwc3Qs5vgVoCT8uzPMcUAnIB1aP6Bhrh3rEfDqwEnOOJ
vS+RHEUscyxQjZ0JkQf4VXukltGAT+jhaXT7uv0JLwTV/aGAuRBE944bDsm7+GzTNw+YZN87HIgL
+TGDMm2oy7KC3sBn2uwa2cDAFA2DTZK66kcH1prXWuilkcQprbGoaEGr/7UJEl7WSYC3Ie++R5qW
MBTPZVARX7gZfQAugEOTzS+qgicFcPOs70FHe3VSJSpydA2K6tfZ7wv1hd2jqP6Xq1P28kZxQprR
19Sq4KPkY2dTvlIhyY0bL0pKdoXuRGVXUjtGFWpkT8GyuVdeacahrgbXxvQF3skPFwmqiA0JN7Lm
igdejXUJZUwBFBpK0cBzfse7Vj85ixcH0nNlfsF/9BBKBIx5pRaAJLtSg8KSRIuLHrbFDxYlgc2K
C4vQnDhygAn76JZcwnNBCcmW3n0/sD1q+twSOOgM85nFB8Wel8IWqdpNSFI7yg87rwSRrksBBBxH
8zK4GBp/Jq023tAt5iFwPzbTQu5jptNtifIF6p/8z7KGVrwp2eU+gYKLhyQNgmcGYdQvlcwML4W0
H4xCyoCNhiIudF4SQkgpZvJm8qrm6mlti9U+F8J5/uzwZf7Mvxk+KNCfpRF2ra7bG1FZvcMBEfEV
bE1ItbC3TbjFDam93uma0/KrC+YbXsSvASW0A6/JMUNQdnz3bIHEwt9DEes1+9x174hDs9XlcfE7
apm6nTaLo+RhXfsfo9mMYR4eRPS3qz6bHx1hVEIB3MTkx8Ml46Ve/4+B4kGfP85/1tWuWY+D5vvE
FNdV3f8onxm6eJtNyqgMsD8HaT8j7HjeBX+SBf7CKinOfM3qmwaYWBPhTqbo0+9QPXIdMB6W08ri
oQtDZArbO7qZRgU/7/rU6mNVJ2XiUYbP/3ryYzPE6NLMl3sPyqXtgZ9HGclUhT8VzIi+urfEaRRX
loCqwhKjwTPefkoTqgHigv+2e58ICkf4wbL8KngTBXgm/aamRkIDVBqud0z8MjfGqmhVWYCESF6A
u1728wbwFIqkv82I5zv8InQFk/pmzRff9P1G5XFx1lroJFcOUFAZls0TT3AOmtG7xASJIRtmHpCn
s13MrN87506QWu50BR6YW4DXlsLniw2QNXmUhMESrlEXm7Wh2qy1GUIQAOb80CpltcB3cHN0FqPc
hYEcrSc/OxNHKCoDjjT3UIAo3Jg9ro6qYEMXJIDwGPE8eNMy/ehvns+ihe2YLjlrnCjAYRurXkAj
45t+Yw1PkcvYwdXo/V79d1N1rucCCyKQ9etZlHa0E0OYQKiGigCli9l5wEI/qQH5Lntssq3P3wls
iPxUDbPXjnioUZvglEwiZiEwLvCA0axeqvu7sMEAUUvPbpOR8pd3npvdB5MLQS9N3IwFcEMtDgLP
roGJPRf7tf1JEbrj/a9CWIQFZdWVRmDjR/eHdg6CFy+qJtT9rPujEtVMQYuRV/hOo9EvLeobfqpJ
aA2F+Fa0+RDo5CY9nADE9DuPG+ZZH0wj1QtzDbAGvsk+S2EpF6vUs8bOpwGZs6DiXX5iCDe3VZkV
UHOF0rAZEXe9sGHUAeDSl0J5KsEl1M1B1bOkYbb47kdC4ltg10Pd6Uyegx56HsAPaOvmPGxhoSRh
szS3xxhmnMgOmzNfZtliYdJHsxkpRXllOGBPe5KgQdfNR5Y8HWsgafBMt5SVrwZ89VRmU5AiDBgB
7E34idmL/ZlaeOakc8TDyKZ/P0aHlPR4lFBvKso/Ir7w2SGnXTlYBvjMCY61W+96uzEOD1yNf0b8
seprpFdJcZe8e8sVVCWGrm1Fmz/1vw+i68H4t4QPKdoGbbbW/LOyMc+jfc/W4DAFRqFWcGLyYGEU
xxUNhzupYF30K7cSW2qIYQWO/8dSwwQFh5j5qpemRWcYTVoZ20o/9/BUajeMSoC7Our0jwhMO8vY
k8JHWbE9+oc0cz9L4l6NmC7fCv8JKt+e1aBqG4k20ZZ+tr2Y4D48Onx9yncPmzsnmKUXmTo5OvVI
0fg+fLqkKdl/VSr/QyHm1bZXreQLWh6W4I/E41REbVUSjnxg2jxW/qQ8sfpUh+95f7+yewZYwjvo
UPyA/9RZm504+tM7xVJgr4g3CUMSDROYQwogPIA5qsG3tHv/RSYD9B5O6V9SQkSzzHE1d8Y+fWhY
XiFRZ+UQJKzdUa87AMLrjbNb6QBnfs2yBxZ5e+Iekqtl7uzi/sdg5i4knJSSujSBdH5OoeNUaqk3
J9Ez0Qvv2TPbQ7ZZlc0B51h0n9dHa9B9mB2wnJA+mVivPmcjnNdzZYF4fbu1wi2RVLw8zpn16tx4
XWD95c6424u8IFHXsQUa7s59A8DDlv5yNVyjbM+b7P3PPZz/Ja3J6Guzjg8Cwgta2thgV+CdHOGU
u6XKpjBy1oGasFSefnaApdsnIe//SXrW8tF0FTGfZRHXXn6Kp/FF5eHLnG4GWHhD9Vnkj1ucMd7b
/WFa39JTQ0zXwJ+RRl0FBMBcb0WbmXcjhqcMFPRGYfAwM/ZWF+GVF2RiWVEraz5wv/mbVohtMCPf
2DpWrjAr61A0LWnK6c4pTLdsZin3VDoqo+JLpFqodpdfe2w/rqtchFUQpDhvQG6D0j5UfIG89zKP
vsyDibZK+sGh5jbIRf1qwq4EsPcz/DaAN4TqiuiwsL4A/m1S6pTlEN8GPcP1I4lD/y/ICJvfKNAl
Od4yomsXFFNceO+HxvrsN1kwrwcBewhpFqhswg5yn1C6+SEmK+15nvJVsMeULflv4+u/8fuNg5fx
UBOeph8invMdRU9/66z0lUSStFiBKBu5oDel6YgajzMOxqyEoz/un/A3UvITUGsNcemTahOeawTt
DIcO2ZOACo3z8CzN6CAk7IVIofjfxhxXSf0lD9IX2+AMbrOBN1ZOriukU1xzXcHd4p8TiJJXf150
QR/7CxGB4uYKYmCVbTnaJSRj4a8nZ5qOU9fqEs41ocjZc75ebVzo5pkX8GSfT0w9MOr4jW8z/n4r
2MdhSN4A772EiLnkv0BAptEIdkntTbBdoHEItXgWrZN0BdfvJOYtAjen/xVU+huuspon1M+WG9on
AA3tvBpghWLC3iWIHi1lQ+yGErBDyo4W1fkKYymfoUs23O02Gkm1ZPRD4H0VCPQ/y/I6Ihix/52f
uFl3sT8l4okNZnXYcDUu31U3jTs55WkCpmeEqfQNGgg6Eey8OgxJ3imrnM07t7+53t6BBwuXm2s5
tVrwD7wb/QlDjPVS0eqnHntb0EdRUYHsKuIZzuOo8bXaRoPc5msLiAMBr4S61WkvEp96REreUYPo
RlU+vtZg14kjovOH1YmzqrOj6rUQ0paJlBir0Xpz3QcDLchGD0cQEwLPLkGg7KzoVY55ziBA4lYi
gNHZxjL8ox50C1pnDDciN4LoFjHO3TuoBKgd6WfNfL2ngz3EsPCFscvwciXwhpYJTD+7xVXDTl2h
K0ovnussDoUakS0iIv4JUikOfOarXMpAQkNyLYPS341AKSK+WMKoQc9m72x6wWVq9JlEze8eRI+k
JY3i4+gws7HfVRAX1w8QxgB3/qPbNjtYHC9LDjOxMeAlFybtpReekQQtEnbKkwTKPtfLdVX/jekw
T0UEab3ApuD78T6T5miSvjRNyPuWQ6MKwWZbiY+GyOExpOq2gdZlz+XUD1u41KvhfEEhfWSHuRdR
5dejsR2nT2xm9+I6THKoGwIke4bomZI+AdI0+c+uIIUgLF4B9cEFxYBwNGC8ygii2LoZ772PoQIU
9WSa+5OdVGwX93Nx9Aph5WVp9jlT9eB9rC3wB7T8qTh3lxN0Bqe7Qb1zxY2/Wykn8cTiDJFv7dbC
fIppjSerIBwoW3qkE9NQw5Mr/Zxvy97Zn+OMyLRoecl2U66qzBPDbeX1nUbyfvpt/Ud5kTv2yjtF
+VzXMyBSn9tZwHEULISP9EBPOKNK57tcad36IT+iIBDI6zRN2kEL0N/3ijzkBriT+SKByMU7QlZF
078RvotjjYeU0wGf5KtJ8wAF8rkrA9tGsQ9CJ4RU+Je7PiyJ77CqFPhyH0ZgESYNCPAGBBGD0AV7
QnTxXyU/qPB3MKYSYAVAgKJ5bchy4+EvUQjX2ozRihcjTV1zAnnt9ss2lc3JewRTB+24lRJPuGP9
p5TF6MVFjpMWdiwhSfYkKtT4I68yDzjWSgYVkOba39sCN/Lv5XM5xtdK286xNLNs9lVOW0wZlVsX
NFiIm76QcKbPtXhtBjvYdDpl2XWbQbB0kdVvkZESZ9mYDxO+HXut9DCy66vX2uefi8mwaKXRfx0r
+c5smWWh5CwnCj4nSYWI+h+IO1HSygHn5hE5+ybWbkJYgB1Ie/9o6wLabeF71eG5dJsV5NSKY/hm
jYc2CRjAaW3Tzag106fy2pyUv1AolM5mzcA4muEhk2SmambcPKJzKLSxtNU+IeZ40IZTR8CKrI6Q
yYXGjwtnUcREP3Tz3gg7VeFDOCV0bB65rkwUcVMv2TshuD8DPiZr+iklbaP/se0J/pHA02ounILi
gOsI1xTA79nnxheYrN4JtOJEjlxmLL/m0KWwHSH945PS7ggEZBLtH32IPd6I2j7YD1gLqPFrGHRX
Ob3V6WalXMI/Cdy6GJeUKbqNrMZY7XPFexXy0JaGRP5/kqUEguXXv7WJoOQXl//Y1n1crqI2PBpD
K+Feo3PzsCL8O7jZJUykidOo38bHctZofvbjLh4LzdZk49w1pCMTzV0fWkVCPh9sbVYbIjT396vI
YWuZ9FynadFKFICyfCX4l1GFciLG83rLHHKsw251Q02TsnY7VTx3eosE8zKskXUek+ARe6CbUsjc
M00V46i2kwg4sjYpxdolCBOJYm4ZGHzS3J6XoxlEIHjgP5ZBJImgA/lbUeYlN5kfPEXE28G9KwHc
v3eV5OzbE0QHagpc2DPEOsO/PEN9Mh6UYwM5UQLpD542yHbirG4kciHmCo/422bA+qBFqm8YBU5V
QmzGLBmn/tR1t5X/wMvHM2tcKqcI2kvqPilFyfwcy5e65Xr1/3WRbWLMbqk9dXB0bcTveqlj7Dmy
pUz5IlM3BxY4ipyosL9BswTa0esXq/R1jQo7u0SiNYq3xhvgFvk5lzxQzCjnIiGbdOchTWntwdWh
Wk79ZV2PK4vqnoS5riiuc+sWrFPC/Bs1Cew7BULppz81u5iD/TgIeu4bZ69hdlo5vufYNhyHYzZB
2KncYfWI02aDJhlBV7PXzYYzv7xy+lSSiMwDY2PKMB8RzQO+0rotM3lY0G7y+/ZayHcJOys0YSAh
wffMImkav+oyJadU1iCvc2NRK53nU8UtYH9wqc8IKJ0VZFHi+2rbYLfQAcHvnaVA+vjHKHYxNmgW
4frWY3fz5vb7wYoDUNg5E2tT/LJT/l6rztSNCCYYaDygN83HVH450MGvTkYj5Bnnm8o+tntaapt0
hBED2aD32/QBRcppy6tsVYwlBpkwkL+Ud28aXE5aal1GGfzN6KuQXTRVRtGTutEyM5Mn11GKYiCW
gXsOtBqiGmyvx4/p/QgAgXynyOcGvnwnyIJ9BNIjNzg1ZEgWRi8A1uuIHse/TmcHDSEEy6fWkup0
d5K7H46dangiDcCLsj7tusijoo3+SMCe39kQYSoSLmncaRV57COfTvgYy5VoqkWZ9CFgLk6vXKXC
xdmNRw3mlg8qqLalUmGNdJVchNTT5NGmPJgKDWACNG+LVVTYjNyFSUb2PdzF7Efa6lcviuot4vaW
hYmBGbcU3j/rLzC4FLPNoiS2X5yABhIafLmpU3PI+zMCrxriCUklu3a3hxhwu55PCFBiR0Bb1oJi
tZ56cUr95ItgBF8hj+z6Jk4HK5EHlzbzd7LJGEDQqZyacrI33W5yfDoyvgCsE/kCIUl6CW3t4wFh
0XDzTgl+6d5BCO/ILu0leoaI2QwGIJXYnJpim6+PKoGz2zD7ptfjtbqupWj3dJjBm/00bIMqWh4P
tf6jjx9D8CBVKu4ZDEZ873p+T8Fb5p/WhLSByZDpa3CWINEP4m7WHC3OiGUAeQDv2cHNlRZg/bld
mxRy79DCHSeCxJlREFj2/etiLRbCIix41A+0N7UQx4aw2SHukSHRvZvpNqVXx2p8sL9M4Ley0MJV
cNN101qYpR4A60flFZJh23Pfr5T7TXwiEQmLwTAz0Y/DWU5gzcCrR24L8oA+piPJkYROwv1AKj8s
W3vuM0jzaOzTe9gmEbsudIwvLLGiPNTgv30Fe+4is7Zn1QG5wbNddHTgqTMjfpvgko9/EZldWh9V
K5bctrvSPuvEhcxUqGAC5q9EvWyiXG8x59MRkjzJ+K7VI1vlHZ0I9dHzc8LkeBI7rOjww8kfDwn0
dXIaq/bzopYIMb5LZo1dbMl62ZUvldJiJJqEQUIKi+0V6pxl9u/0zmPMx+kW9LoChjGtM6WkUzCy
6gLdqQraYRXzywagUIpJesBWPwpsHfmfCW8j69G5wQ7XRPKy5AUGusyk3fshaVziM0O/0s9VP1yl
Ow7Ql9WifCkfjV9VTztqaNo0RmKRLscNb0hTGY5dYW5/QMxrQXOSe+diwMcllg/R9gTO64hZXdG8
SeCbCyQIL/m+RJei8xg1/1mHkhTLlLpCSaSLOQAkF2mmeI2E+vT0sR15opEttbvSUUdsWXxLXK61
6EgGXrGe6GiEEZQ4iC8f+V+2qGIPCZQnI40XybubknbaH/prPsUkq/5e1HjtdsFvjh+ZX1dszIMq
mdyRhsEfcVDPtMWzR8o9VEGkSwTnm/VfuRPvvODsaTtyJqa/YUN5tzkFXppANoPOwjwxi0fEE+Ke
ISy7vpAuu8k2PFx2BPBHiJFQUFfEK1f0yH828wnmmF7ds2oyUw7Lji0IqumxbZCFc+i3RPgO+CcM
+EFehyYRJd+xLiK5+J5H8eM6oxO3+ogzrUEFkzzPbkVuNfzvIPDT773rihJGMFAQInpnDYFkOVgA
6i6zSCvf34Sp50PWY4mb9h4L1bwGjIpAF0y08NYShwSUPsEfn0IP/H0i891ZYYudw246Yhk7Ll2C
+em5Un38+SEmZLxFEIUmnsEGfnFRkuhq1u9EqB4vMlM3PYJSIvQ799Nm3fUAVw+m1rSNYRW79lZS
G8G70xHhPVDQ2m0KBlA9PmNQzTz8ZitiQhTuEVDxOV2OS1lfwXMJk2oizJMcMnpEEqup7vSknq4U
OYIIe3tDbHT80pS7T9Ds2pGa1Monvpz+U/YV8531c7ujVT6owbTQgw80xN4kGcyc8qCJijA3N7Wl
LiOotF1UDbH/KBBOfYr6bj0b9VRoEGPWOQYpTMIqWg6BkeWG/B4jkc9GACLCZFj+bZ9IO/nyv9wM
FvjKwVVoOwBU7/2NKc/nlUavKpfH+qIBwNC1BMRSyJK4Sf270thPG06vxyZmkcj3f29ktbShGna8
CZnT53WJp5RQB9SdSzhfho4UIJsycbFbyVEgCyMAzzEFVvqKO3Ov9em5pocwLFNPjAV6kZUM9S8V
A0b7WiqRTFwBYSpjYfCq47rG6bCusUKJiQu8Odma8/tMeRi5aDQX/83FvoSq2R4AubrRfh+Dwumi
Vsn3rQCk0P17qA9vBbVhu0fxaVHYUEKy5zwlC1bcbl816b+uBdD3JVa+BC50wbKHZGe/MKFkfdaK
abR5aoTXvXMtCgANHXtNAV36jJCyJZ+mWdJApq2tqVL4igBh5X/XV/K7N3SrgUI09JEIbda1Z0im
iGYWaS9JWniQN1vHnDNL/j7xycxJPr4FYk2A/ppGkK2N66agB+OmnDZeYXwu0nDcFff6AQAlMFor
qkWeH/JkBUfErAJeTQ+HnIlbYJHlwFFq4B1C+EDl2ltJUwLsG7N13mAWBfxgVUu41AUeTU/iajhf
gyPyanWyCkOEKN9fp7CrtGXyDMMQ14rIWK06fJXZFGO4+sjFG5HwcX4QFGJznDdzE/1OuKWhuMdb
erP2qrq+Tyx90WctvSd+zjVfqPRruVO6XDE+UGwwyhNVBDa4QKU1VY1fkVfT4SNJoj6jzYPREdgC
P7Jcr+1cCEiH99AD1yi+xoSquxuRcY+NSWHmBkSdGGAVpMQ4f08wp7ExG+nmMevYkUC/lLhzcONp
UZF0mlikK1mQdLmWkJ19xPxq4K9HFKjWpOuX0X64gealoT3DDHD2Q2qXQel7j6KeHZu/+CedIElo
CWGuMJgUCOFAUp+Zrpa3isB6nwARcdIQvOgOiejl17g/YuqspJCfAXeG4rhYoL3cL2kLrqh3ItXl
D5x2rQRovIWf3AvhwPT6aDDJmeaCChVwUs3+J6+igwYb+GQ1V4izQyGvX7zJ3ZQjjXCfkei1+MpN
KExii5UTh8WkpzspQmFjoQwDRAtHBz6mKP0ThGWQsxETGHNHllIduKDWUqIVq6dU6Z+OzECV8qA3
PD7nEWnM4Hai5nWUxyqhhkyDDZLWPAPt7E7NzYAoZ7B0LYg1xXuZHF4CgJ/FhD2VmdMmFV0STwAR
SMX7f+raHfKSiv/5lXzsLH1u9sJ5KcNQX8rsx7wifPEv4GTvIKa6/ySzZZU8QCvOQeYgMk4U8ttV
25+rMqZuoIr00/WZzCS70vgKCzDrlqI5ZFq+Am1UGz3ptsbv2m7UmKd0FIUUTXQyANb45veqpAo+
CXUXOYHX80Hyo4WwshZ4A3tRXyaw8KiCNC+l4jRSpw2EnpAsxehriwx1gZMlu146k1026k3BxGKY
EnRgUnpgbZfxyQUoQP6ewk/hgIcVwDjy9jb6xnA7hQJcWQoRDjfHvhC8yOB74wTk9zN1Z7D3zZGR
4JxxZt7rhIhSXMPuDOzgTK8I+wXEkNJThgqFqbavoqT+O3prCb/nrddeuSJ5BhU/jB/9Ol1tE49M
mbnGbQqa0+25ELxAecC7i9k2kixmWBbjIJU4X7bcKWzEb2HE09oypiFFlT+Y6MqaRQjJ87grdhxi
phICMpCZAOhOUfZrZdiZ2RRZDO162RG6unECCSFz6z8/38Yoe/kAAatherbGnUJNsxgHskNO/zro
Tio4ZM83xI6YaUQGkFiol18NUqt0UWH+a6aRjyejAxtffjAH30Njqve2rTLd44Eq0AhWlYYz4m6s
86b/LFJ+4/xalnwcCmCugJPhW4sbFShdOfllzriOjs7DxQRpb5uoHIlN2itY5yB6t+dK6ft6G1X8
Kj+H43j+fblBzat0y2i5xa+6VLMxtZS9Y18MCPKoNepFWcdXGu6OVV3Lo2HxVMYRXSpE0pp68ufd
Olg/NVAfmRhpAGZuG7ajqePWVet3Vvr/lGCGiXWZXhd+RfrJ+WEz440wi9+PnlST3YiSBls8Xlh/
KHcsVrRQVZBuDJY0e4dnPYTKMQOIUYvApeuHnUiKldaBMqgVlrAX4zaD3Gu1XE9XRFeCzgGv7EUe
+rIcRVJ/UNf5HccGx9dzeXpRd/2sa+zvfuxpQwXVb7ucOOkpjl5t57MbFqV+F0yO5KwKtfPAB8KN
OyNeetI1hMdM20P09uaurfnw7TFsSywZV2qHYaxmDqUJw2lwPWrzaCf11bSwExLcI5REXbOIhVai
NiuHJi5hLnio/0Dbq5nJXWF7jL0FeX1pIAfGBEcoSCUlosG9kZOL8NF2fB5Uyt3A7hlK+r4Wojx9
1pcxObCuqgcXUT3yhbpRti8clP61tNW4aTSVf4RxHdpJIhq46zMIUGI3VmxFfh2hhOluVbOmtbGK
baAf2wsY969SIhXRLH6BDb5vcxvFVy0iqLXivIf/tydgpY/+BZuXC4qa5zCcCrsQHgA8FoNkp/7I
l/R/l6c1PAXWmrlW4TAx47Q+6lo0GpFPhW3WtsTz8cVW08355mo2UnUW95KOyc4ik+ZR91o5LGYc
Sm6Odb61PiWFrSK+9KLjA0ARKDrBb/Po6Pb6KnndO0IN58IzODM3FSBkyRCzYHt7WHS6YyQPO8og
qWCJxHBMozbi8UL9Pfd+jHX0JZUiLk+n2vIP1y7mFK8jSOPPZBa2ExnVlaHrEg7dvHGJiTITDqVF
c7Wj4wR69TZFDNNnD1m/Y/WOoxZvbYVBNGSYJt2dD3zmOjgu1VB5BA5aWv+3nYj/QEkvqdY62cei
bhxlDdmsiYVXly70Z+QwL4aH6uMM7QuX+AKuc0pB/HJfFeHq0PuypBAM202pYWm9ifGxeBngk13y
gM6kkHrK5hEQmOTxtunz9hVGghnFm0rtczZyJL7wjdwQM2CYYK41Sd+b/Q3W3Lm2/WuEPWvTvVyr
6gzB6cVzrfz6nZwBfOIqmvbIM3UpFI1sFhWCvuWijcr61cB1JBcStaWmXEyIrHmTnlojG86hwrWg
4h9nMt48Grd1bpDXCueFIzaJUmaYvXk1z1euhyB6Hvaeiqi8nV8M9Ddpb3QZM3yBFESF9GRXM6nT
iA+ZBPlLt2wLxCkNtDo0Zmk2Th0oqhusZ9IeQda/fmwXMMxiIzwFgsPJ3E2F/+ip1SxWjb/RwRZE
a3DFYeFO87/t7U6P+71aIH198u/Zry9GRyncqVyOJDDSDZ9J/POSZVrEZraaUO1RX8+6G3R7c2FD
vnffOkSqj0vUhZ6413+QaliVptXX8PuNpDVLihj/Fk74eaBKoUxTnW563G0oWuuJy+ZpSShgPqm6
RVSIZXxJtaZagkvOan+Nq3ljRhRKAHYBA9KCWgDe67ZRYC2ahm9W2DoBNvoQe2g3FxUsBpDSCZon
mMthtQe6a8kF8ApmHiKLFd9rhzNSoAuqux6AhFUO61V7oX2lHnsUPZS4MAC08I25lyEAffF2DGzR
a2yZkXwzxW7A4XvNCko7MNEdT/Xf4N+KxN8aBePV4HNh86as1oH9knmuuafeJ4Rx7wECjC11bE44
6unrI8JmGDUzeDTcRMymej/D2TcU30zhQ2d5jhAlh2EwHOIb80r6yakBhe2MJ57Nbnxklub4dpgL
R3joHPWdb5q72J7Rhkahom216Coetf7aWx6t+vXSaXEfQxsvrFWLHlHQTv6GcLjt+kDWhMZb20GW
pUS78DvX1K5qaaWtXxVC7vDtoUp6Ipo4gMyZyVdQwEfh1VrgKJ0A9/QDatwDppyXb2JBPP2S8nlG
aG3jpS30rzv8WbRDl4IBNalFmAXhBmtcDtz1RbhHyaDJaa2ru+cr/dsfJ2IFGuWBoP0vSNo3Or+B
aUMFTz+VwKSmTVKnya0XKXc+F2ENYzYBUhqDgcobhFPIAlZprK3EYXEApus/+ha3wqdubGRUSC4u
5Gph4DmzVyGzdDKlWkuDH90E9NGeRDVZGcoxuQgNmwYDwqFJh6Eoe4z27N2zncrAZJR2bC4aIUuu
ZPKJJLsP3pJ52Tn/rC+cjkLoCxuVDsQo9Mpme7eRzhphL8GSqyBS2dZW95SmnBy/YX+NaMWWI/ZD
TDM+8oY24zqiKYFLUcQ0lLcXnq5ix0eszgi7CY8le4ImcGgxG10nDAdyvXdJzbIbZBQYs+zXmBE6
/XKDn9gDJX4v0UYaHRo0+y9xWU83cfQd0KWPuDV8YMUl2ppu6cPcZERo2uzj5aneihVvHR9uu5ZO
7dHCVb7SfMlDmzmjZCD09iGIk6qcjf1pEpqUtnNRBkv1nqLt1wYcz5T78zfyhZKeYVHAcVpcHBEc
Wt9Rvao0s5D/2zH4tVQvvPGehU2Udt3YqGM3zIG9DvFK2cCoM2KBOlHMjkJ/a7THspQW9GDwF5O1
8WBDWFzpWGPM5YYS8NA8J60fCMqkQwcWGEtaKq/wB+7kGFSS3AW9H0y5xaUq4pB+2OTcdOWu8RQ/
slNNwyh08y4A0fl3NgC5Bh0Flv14xLdc5y74XuO1UqQ35chOFnN4UIJh/tr+zhH7Jnu9xhkVuhAR
T+VwMcXKYn2lUuzcauBZiEn6KBHWTvLK4bkB402KVabSmSyF+pBUq1oOMJA0ZxtbOW+FfwMm3FAL
iYs4Qdp6qkfnQf8A3oghFK1DtAdA3jGtlqoiZ+xS8tRlVkVZoU4/spe1DC0ikbm0ufZ1GVlKQw3V
83aphlumIjOJDIRbxUbD6ZgnBP3jGqxBYYY4Akm8fsbz5qYE2LvL9WrT78Fpbixpw6vtWApfRUB5
q5hB1sObmzh9Z8koq6BpDJHg0BkH3EUQaAESk48HYXS498k3JwhrXZzvX7UEeEIg/X1hgV5iU1sx
LBGUmUjdSa+3ssxU4DflXHgPHNPk6qTPc4Khxy5J2pYUtTfs0H+VDId+OvHyqWM8ixq5gd9s7/FF
iFtCSWAyIuyIOegP7xRWw2jHeqP6oyPua736IBRKW/Ki+ahjRTmzGSWoBpfJMYwglOhPhMp4T6GS
b23KqrBM8xs03lDIq+O8YwMRizuRnN7dVosHPE+vxyTmO7JLzxZ4vYoerc8hfJIa905Tk26rf4KO
kmtGiNBvKPAb2BBzSwmS4sHIjba/0UdRF9ZJt2UEFliQzYE0XEK/vIY9yFDqXNXpqL/DX4jCnILQ
TCEjqJUKMYyBEH+OjJItUjBilbsDVy0+HAlVVTI5xMpZ2uXfHi2sdL/B6vWOGcVtn1C8NUm5WV4V
/BUEU0A6UobRhDJ/lpc9iwbCXnxgPp3ZZ5TcziAlO9LGDQhk5se9dTSgf79GbHdhtef57DWGJsVu
gTCBF3PRJ5cphN/zmaBompytDQKFjCS2xnHSiqslN9hcolScT54ubYZiLn9T8n2cyRpIH+qFvCJ3
r4296+CyGogmxmeFVZ6BEzwNfJ0FNXLndgoe5Utiq8m/kjjPqMyW+f0oQ7aH2BT/DkOoi437mpD7
06spEHS/1MXK/l7rTkMX44GnA9TLFubRLqjfwCJ2x5kldewk4iWO9BrqZ2/tVrdanM6wAJ5Jp6Gp
HX5ysNXSzciwYclE3IRL1EL4EAXlNRnviP+9acNJN41bm+p7wibaSCIdw6ftTU0B22zqoPIZrYKX
l4UqgJ581+wouPNmtjr5jTf+NpnctzStSynN70k86Bd7l2PgC146XE/4o4Apd+k4iyfvtLLZ73Zr
QnsAhfxKsaoW1hdyT6ig1yWvcSZL9wCAjlBnnEQ9p3mP2Nao3pAL/OtdH1et878IxeRIN7J+tM0v
YFF0j6gKEBMVMX3gZ3/zrDgL0Ke+Cyx+C6WG/hcVICAq1hlm37aWrmKP+Q23FX+8Booe3KAxveA5
c4dBtw+9Gdlt9FwoZP21Z6/G3vNcHd9CMpZKpZ4uUe7rrqZdvzzVfyBVclgLf+4XAgstEJJxpAFI
VAyC/bokfhdLj1a+aCGPE+I9mjk6cm5vH18oDUzOQF83ILy7lqQDfeuGmuPq8oFlF628MZLFCGJv
4Skv/5/rKIQH4tUMxJFNLcERa7la1+lhfq6EX69tjAsjrA6b0ahxB/12ZA/p7Tn+ZnKyvldBZ+Dc
l1juvqOa564ZUtNXYoAl2vrcX7js1p3NwZZiT0ocAo66IFeieu+mEqmndrV1lXKjysbmQaqkWxda
4jGOgZUq8x94CFQxa/EUPrB30EaY8A8Z2FKvjT18U1Bl3ue/eh5+M+3VGB6OLwxdHDh7EMOi5JPK
99KEn+S+scpNFAVQkVNhJ9RlY22ZRAVKg3c/TNla1GiXZFlJEwHEeENvb5Qo2lWun14K7atHKSiu
YjNjTR00anl3MRXBBd4qKQF4RT4tguSm68RwXmzyF+PxAXRYg0iQ19QGI2yuhhto5jwrn0/oY5GC
XQNtx9u+PDGqh2gl4WGLpRvmE2YWVA3YpgQ+3mYU/BuppVAdDtFIpTR2/FUPPbmNDijCe1MDG7k0
FBrmSwHC8cTr8so5VUTaiMXDpzmAYvAtZX7OgE+Rw02Oe3bRD3eyMe1AihgIej8Ovu3LpCCWG2ND
tqSvusC0apjSHUxB8E/hRFBQw6A7SM4przYmlGklbsQ6TyQje/GO1Nsr5JZTRPR5h0QgxVhQSYLs
sEsftCtqJS0lR1V0sPYs+TLg4e2ZC7IaAhL1k8L7MW2bJ3oKxRXS3kuGQL+oCE3mRvWBG3HFypkf
Ja+Wa9pU8/88NvdF1s3cVazwWMtQtDu7/oJnOL0K3QmoMGfROu8GbQZOoCHKfox2A9W2TuaDNxvq
uH3FYcQ1gf3rf4n9zjROkwk9/tstXbI7JbRe8dFyl2B+tJTclAA8v9Zl0+lPtE0WiV40Nr5eRIzw
hzOMpNtZyQUb6TSd+pbtya/2dJgvbyb1Oh+AADm1zZFis3AeYU5bduqnwJYrk5cHhB32aXrrOARq
ARxaAwFVQPS6ThpodMaINN6YgGFBmKHzdOXrP6XrNcEqWV+2aNjkGVEFXbwo1OUJGecXA0Rm+HiC
c55NmqqiXAZMXkLdCXhjf5uTgjHmazO/kfBv1ZJAICYSj1C6qo8w1JgNjpCeEqunChGrFcoBJFl+
8c/r1S9xA5DKYaKUumoRBR4exzAPhqBTI+80nL7pneGhKqBDljYWnkoZJlzsNcHfpu8s0OJGVqs2
eQcOE5+3vdH12uD9p+YisJvscYGuA+BW1llnUwvPjTFTkb+6Lthnktz/Ga5OlATZYRtcgMBWcOr0
YpYRoE8Oq1ugbm9yZx8GOCAT7fz2+ytk5pS7Zn7jW5AUL50udKO+hmJHoyg3NQcITYqnL6Kx83RU
vCVyplU/Lc32S41GtYn7M7aDVfogiAY4Ax9F7kb//54V6u0PI7VUFfsgGqClNLZG39vx0am0uQEY
UorKGyzOWYncx1hAQBag6Qj6fXP58ZFvvCbAlSQddrmeWyH5ag1QK2FBtXqffss6tRV0BTd1voxQ
lueDufznuG7JusYSxa1mVxmB1Y//JjbAjVPPnr+AW8MBLapQ/hOVcWW8Q1Fe0gcuiJb+9s4Q9TMx
/tB74zegtjcytsWX9fVfz/ckaMt9uA6oE/lH7bsjtcLDuhYbrWeN2SHWbFAuGkRf5eG/IWEFAV7q
4H1rZXpsbwbHfWqSnIytKJb5HEFFMOj9psJjUFlwkTmhhxOlIieeacxii0IFtL69hj8BvFA5Gh0O
hgg332frGk6i7UX4+J3+tXCP88RXr69U64OF4iDos1ucVU2RxXJRTsIIeOE7yIyh+gsuXTph2SGm
IcQ/Jsa77KyzF1DlNR5pSqa6AgyFknNC/NksiDP8DNBn4KVSqdmXmRPehHS/rxceNwuzrikGvvne
wwk7chpkVkOGxtv9+tnxoVTYmCOsAzVOrG0xqLMABa3SiX5Tz9brSo4o2wJpJLmvAjDTCRxoH190
xG11Yv1/eBQBQbQv8DOnV2oZnp0sMbPRbMl+MMfncGbiSjhxvHKvtbQchPYzVqDSybWC9gvEyjrS
03HiUDvUZ4J3baFBG2P0cXHzm8nrMQI2J9F4B6jo/dRvmQfGMNtbJ+UliFBcokVPeC0Y6Q4WgdNt
Z3uxeJO5iolZ06iiYilNPtMHz5Up27IuJTsRIpx/+5T1dGKzEYqnyaAg2K63pan3u3TcNG0j/Uql
IJLLrP/1LEHHgC4FBjw8lIIOZ4Gu5xC/VlqwJbOAyMJ35is94hMC+nDwmC8q171JCSoKItOLMJtY
UhGQ5W932h0gAYMsoITx7wUDY18FpgGpfQ3YRiqBdLz1Y+cF3wV5IjtikpNJKFprH4Mv83P9vDAT
rCFQOxolQ0Y48O22QKufBEVaZLo/39kpI7k64f6HfG4J+V9AtVLgKJFfwKCyRKQlV9bbDAC8cfP4
neMF103IAK1ZQFmK8L4gepxN019fvj2XF0u3Bl2Z10QXe7BF+HVIPFc3f10SUc2YmSzNUCyp9dZB
7d4GBMmAZy/EddkAx8wWgGqebr8sPtzy3UigpZvi2GlZPbNksCivxjSGYBEozMRD4otEGYn44vIX
t7N7G84eB52x1uaTHwRY8L0JjPcxrff8nRKx1PYt1AbbV+BTzpbpGBMEvuSMK8IA7LZ2dhToanKQ
rBvoM7YHiKybyFrb6GEPAeRBx7JJwJm99hAM2WXzlSHlbDEZrKo1EKU0dTfG6c8rFICNRXHjcid9
PBfVEp93/iwMZ3q/KbPk+CPBATAq9+4g1LKZeyh1aukdHXNeQeSEotnCWj+21WxQqjAIjVVUQebV
F+wJkEAe6EkqoG/Gwd8Qp5k8p4XPCoeojl1MpASaVg5HPje9h0ff6dB8qFnUOCKGYKQ0qJNuKk8e
A/vjwQsNH+o6vTgYWsOoplYnaWw4DiQwAEuIZRqRTbYxoLWRNVvXSCBk420VDof3/XdxYTLnC2/U
KZhV28p8qiqCwpYg4Wsa7yU2k+WXB/+TR7KxbzRnjga6FqfXDTHwlHvGD12HFjxBuGIQHp61XaSo
ZNzJnM9A/Eryw3uWRbbDHk//jTNPky07vCiwIfSew0ZZNhyt4zhtCI+5Owr+3WV7VM6Rc2oCOcBg
AUGlgqcAIQ2MGWy/iGS2/O1CFq5ThlO+GXwBuTB01CjUYTfvueTyJ9bsyUxcLs9Ux6F2fDJupGGE
00M/zwnY/oQbIbI7sQD0ymQ/LN+R2G+lmaVRVeMzmJBdln7lk01cRiVyef2M94Nc7sNTqVaskCDa
+p4E1g1aEfVYIpCYiK8HzkHC2qoRLHTd7Pi4G2loBjjzmJ7bi5bKHRaGJnNCZOOVdO5MA0JAZmJ+
u1+1nZN+606XfmGqbCTxeP1LBN5eyRAp9PTs+MsWZ5X8V3CWOAVGbL5koit9KgtcnXZdMrBhvJ6G
CKHPlsGEmvPKXlDbX7TiNyiHPb2jNH/jUHUMhQCcDLlkK5h5Lb2Yf7B4+33V4WERDwCQ+mQ5TIzA
Jvgs6k8aHTHRf3k306lFzfh3Bg6HGhv+zb0q9Rh0FtJAyv9z5+UTn07eAiafZp0uZGGyhFSJD9G4
CcfK1AhrjEDZvxUnpXfse0DEMKhDTnGSGiItgnIKlYEqyn7RmfzJiAXBKnBwf5tZbC3Imx+Mhxdn
KsL4s3B1EDN//e8kEKyQ2DD2bbtCurihmjAmSomx1zZDE3ijgWxFAGyp/vCQP1kVL2jbeoCiaAV1
QPDjqtLHRIN7gHBnN/WjZl/BqV44iqwNN++MIhqf21AJ37yjsoykzgGW5sQRVIeYkPbVFLMfK1tI
Y0QJzhQwrSrYf1AhFkUbMJN8OVSizYcwktRP9AXeBG4fb4wYA6P7/QX8/7arw2/OHpF8la0+OlxX
3LK9/sW+Mr9wYW76BWqo+kDMsZ0mdgd5/Db7Ziz/ywE6YMxyR+MH++kz1mIgcv8WRYKJHfu+nbBb
IEJwWtsJC+uYgEh5/8Wky35VTFpjXWqAs+y7WOXi4zJ501dRBYlIgpV5UjiR0unFPoZSAhtoQi9J
8MKWf+/5/91c+H3UX8QyLSrsnJTDdRgvm/hCxaSJA5ffmeJ2HtoZ8RxKbLqyhoplN+VEjdoBkwaf
9P55bqhEPlw7pGwOwEx+v/iYRAdlVlTX7o+KShV60DkeJ6UQ8OuLk7fN7ubc0Dl4HPdG5ZHhgM9k
jnVX1jDb0s1ibCP4ZE8tPKwyQOg8Bvjn/CS3gWUx/fgQs3zt+oFFD9LTTxCwBK7sqLYFkbwVRXZu
g3qbUnXj0HKB3oyKU7M6lUWAbL4YHhLzzjGcRqu8FSr4WZBBFJVu4zbuUXC/p541SlTqUZAlgfF0
wa/LiDb14y2ikaAFwsgC5fj9MjuFeiScFwd/kJA7lBm9NKQDK1PCi+dy4x7Ek+BUg5TmxlWuZYr4
/oEyPxF27z+4hi6YnrbmVLp4x+CPAhzYxw2CteDvaag4pgzITyW9HHtKEahJ6csHZEzhvzfj7g7Q
18tlRbT7KWTiCn0W9Amjq1YAkscurBn+Rs/rubpjMCGM3pqgldClVCaXq8WJc2YRVJa3RE+bYU4X
bMk86xNHksXNm3mdBqNOyznV87U9rzhUMVVpiv7h2voPw2qtD0GWg3XUUsd888tEBOcdmN2S55R2
0xQ51WzujbighulL6Yz2qMVRL1wmJFCyC0e3nOD7tY+JCrPMWi9FtBCgCJJ10JFPTFLwZfgunIq5
khHfOt5hJUKr5nTLRYM9sbI0OLFS90tbSqshfQZwZWc52XpRiR4rpi+Tj4gG7vIQW+1Sv/Vf0fOP
wkDUI+0PZ9JBtQGts7P2SJnNnL/E6aFjAczsfLb8REdNvzxlouEs763tdkL46GkkuKC/ZXLlUivx
vvX4ZhOAMgCcmQ5+/MWpm5NaEAIRWYhscIgTq7xc7d0Xkyxe6b9i0A7vqiVw8sPqEaMnUMAZMe6Z
z3K5Z/NsrKddt5lzmzRsQ+VpuSLfnngXJVtbKjyt6zDHQVMTGldxYXhC+KmIn80XbE61e2a3KoVs
C05kP56sDOC0mr0Wu3Aq0TfqZD7kFdTo4gtHO4pgJYbfLsJvUCizhWUL4xSbuTWsdCWCCzZxUJG9
LrEeWVYVWnG8X6MhuNuGRehX//vbRJv/Zk6fOhIB3ivBoIXH42eMdKknj7RrN9U0rpX/CH00iA5k
OetRP5KqoaFzohvi3HZrgkGafT4smflUmSbm7jNcsJXpqqTF9aasVKF5eN0SerzJ8P6uoDWcLYRy
6gkHyFdNSdgnlfyXQoDB5TychsvDrkf3IfS2dz76HtahFAZX+inWO1gmkb0OWWEfuWAzSFf0zgTN
9AetaydFbZ0v2fgG2WhEF/WJqzXReQkxQ89ZCPU5c3v0UAehAAw5t/HzTBlxfzTflAFpUBR8UmQD
tfswLQnf6xBVrXnYlEl/chZVcfZRz+zS6JHm5UrHPLGEHMQXC5BdPzg3qHvEUYpTPDRAX/0l2I9+
pVQ7jmCtuAQV81I1tXgDQMXNCfKBGdxeHs0fRAAY+EkpstHgbcxQWo755dcfmIZNxI+kVgf27ylc
mJ+ZvRjw+2HTsG+l7QZBjAylIhCqpEbxwzAn//ZLvrTr4d+aW8RnxqVV5V/efwl+IED/A2ymqz5Y
k5I9tW3c2/fCF7+tKyKUKm46hBUnM8tu6n1ksAZsZ34r6uNOvHgphCaPrjjgjIM4w8aphTLJTLe6
2itffsZVV3U7Cd7P4y/yvbYVfmgijZ3jgYyhaQJKxk15Ls9E/rGdcAhgoTI/p6vBltiliVzDNyOR
caOsPI3DJqqPkB0zqdtHpIj2ENIUY7GBy/UmrdMkmdqb/R4ou3nKpE/EV+BwormYQyOQZcOYZlPB
X4t/ZbMYanACX65HhEe3JQE24xyDGm3pZDiEqS4MJXYjfK7qZ/JN1hdH3vRJ8hM9DT8vPoPgStsG
/0DfJnnRrUiTj8s87ASZuR5hsnmUsaiS19+EpmcYeZA8LW4LkbMs7pKZKkhlO+xvn7p+YorcdqaR
VnY5DKVWQcfEOqQ5TfA1sJcqlx9rg8FB5kc4FwFPxc/If2TGw13dABDKUdq+464eenmrRofDpHFQ
OUoq+Qdk0Ndw8Hhi2og4WnV9lO7y8BbHuJKLswBPBlJSOe86PSTekn0Jd8eOYAcOMgII3BZFJtZG
eh3nvR+jFHcSBg70ryv0IXM7S/dXWmVwDHhsdbKIl5hD6XbK9GE8OWq5OLqob++20gfXVGuHCgT/
fGseXPOdVl6etubuWxcCzPPwL7uJsPsmxZTWPxvC+9JTziB9h4TH81q5A2rVZXmqg/nVIjHyuSnj
GTzTjrjTMqXy4d+B0ppWTaveA/g4a+bhiuu8Hhj8GYHzZfIVMWJWz/ub2aORlXvzVDgzfv60gPJm
y/8xmY/reR698w+LXCicE0lHiedd5Te55jKtLUBJZ+os8K78b2pwbj9bURKCot9E+7XyL4by9aax
2CSy3mrEu/xnCwCzKpVL3xAXbmIoo0fOmc12TgUn7tjkjwNo+bV1EB2/ax4ncJk4wjxx+bjHi9wR
RSbzbX79GSPKvZdVsEfxq/kjrk9j7o79eJ0kkaLzfEQwmpv+VkTt/Wuygp/UCukh/2Q7Lh8GLm0S
SaitcJp84nlvoyvx+Ds416MQCT5aNNe+H4YLKFV6AKWa4qGk85qNkibZbSlbVpu5aI+DD1bWPdp7
Fz5nEJ+CSkDl8KzZcHsvOEr1cf+Vi7K8b2HM5QFBwexB83DD4Rhk4mz3jTy7MZ78qj4hOU5nBt1J
LQw2/fLcphrjNWx1maCqRZtQSPpqeXdNwwCSxTF0ab3YpbmH6Ny7rJwyyZ24Nrqqki8jNV1QonXA
NWWazb8rbE8D28GTulxd4Au73VCFoBEIdwsVKvellDQ1qWkRJQ9KSQFjaUcDWeOELF4oOy32K9CU
DGPuaZ7KGGhQqmjoc3POQGixu5vjzy7NKua1DT0JevpKP2rBJuiLaXAfNrXAkXH8wu2ovlP87WZJ
V6wJJshB2iy5aIfiBwpKPXt+aYp9+/1605yFTXA5MsorkZE9HYwYacsKvq6Go+7MBt3jcHtnyMvI
hd+fWoPyB7ER2tFYJr0OrIkeFqU6ApSlrv/unXgyyGHToTD1HG9ZHgUCFXzPWMqSbBqDC+Q+K2yb
PT5iXepEmlwOHDYpHr68ZiioziN0zRqB62pOdxkmzonWWQtIkloxj0O2moC51p1m0G1WG1jpPZRI
XXMPSxSuk/PIEsPgCuAMVDQY2PR6n8AwMkzds+RbqUROVJfch0lE6vfnaaAXeAtfiE9E3dyenial
cm2sN2kXn6I6cUqyG7mJ8Sa5bZhazlwHolc6xYRZ/Ni5I+r9MKLktFuS44IqjMPkdUdxG7CgYhOh
gvzBJmUEEZPdXCb0H0uko9603/jOJnLe0RqdP69yBze4S1SuxUlhMZ+fIkhLJS8TVTIU5WF3bHR9
yE2C6zbJIw/7Ab9nt8RJsvE/Zvc9JU9/r4ijLY6LCfwwIpLOemD0gns8AXSjQypxhNHLo6BdV/Ng
WsKUlWSEJxcXnMFxnARJXrq1SjWztRIp6pjkJCXxIQp+uVU9f+wscmXaPXlKbJdVkAucE9wj6Nos
V3RwsemChYvIsA3pIECAs0Or5Qc1ReHrmjHZWQuUGovVG4Ad9WP9HVeBoemIXKlF1uFed3fYnzIn
MsXVQBL66EpH924H/jF1fcTsdg1kUlLOCBC/2J0W7ccV5i7CSOe+n+4RynxM4Yk05JIxd2auRPDX
1C3IWQuyU0ml1dPA2MD4stDGVWew7exWFf+V/gHuNdC/9SWIraNjtMJdkZ1FcVqDyLoqFDiva8ja
l3LxRMfwkF0o51BmIDBYDj65FTBBWAob+dq1CpOKqn+CBWMNcaDrFqdKD+++oGkwThWEsW8AG9Aw
W8f6J9ncI96505U9Fsiny5qzkzk6NLXcyznmh+cD/NBX4hX29inYVhR0ikfvwKgBQiftnLonmQFt
s3W1JOFZEgnLbBNoy9QuS2YBKFC8BowhjSoKTm0BiOuYG8pKgb7aqx7yFFHYPYm2YYh1W7Cw2C/t
/TFMtAo2UvfI5EBoab3GullcUp3eHHN2MjmSOQYsSRmu8Zg15oFHmf+zY2maU/E6NVP3P/xuZS7b
igbtbY5D1f7uWu2R3ZB+LCtoRv1afDPUPT85JTcu+Rutr4MfVlh9x2IRXFoC7gWTB6W9QQec49tY
UPQ933PdY60M1S0QDr0ZINRV+/E1POcjSxkLBosYPtASLuxihKe36NoeNxZ+tqwM7YsNlLNFseHq
nZ50NWfRVn895xr6dAjRvtDq46uYbVYBI3uD9993YcwsrNF63MMs+av3ju2KS0esZG+5wEVjXgml
uNTHAnLoohtkbXdOEfjMAO95VE4UTG+zxG/BebM8xYEb83RN8VPZ2KGdM7fLqMK1r7ZE2aVZ15dg
WIP5ZhjsRn9G8zcOh1PbdSvoPxtW1w4yWr5KcmAzvfg4eK7GtjY2Z+mRtKujdvjB6Jq6zCduI1d2
desi2coO7AQmMmhyIBEadvVu1B02CbXXS6jqSldIBhkNaM3fw9l2VyoV18A0jSMvKp2ZgRQwm9Tu
+BDK3xteZS/BcvLTKioySS7OjEiv9BP3cQAnY5257B0zYdFfGecEVUS51LkClZAabrKQykA/9HAf
4vi5/EeEI97XGwb8+62a9cubvy80PVxOszawclZy3ReaOFhM0Kd9boHt+PR2x3MIcUkvOpT6cqW1
S4mlIxuw47ey76+8P5E7L+iHIo+OH+TXTi5RTgf8Cf1nTZ/YBy4rhV9I3lQULw1Z05u9CI6HPrW5
q9Xwrzd+PJh1tNNTTtJ5rmwtr3jrgqMlXFB1LJthAYHGVqnITvD46IscZol0A0m3w8d4J+BSGOA2
xrD5YmL2dShzQhFmykOebDxNjsTn7siX+gT9TYM0xYeX7a+mzZUBErhPfQNPTCgzb2FeWu1JFtUp
1vMP5RfrbNSSsht33NwoCXFuXkbPDqChY33EZHqZ0DJfZdb6kmS8eB0EIjHHPvNlzOXMnRhwvmRV
qV/RDcGkdBpaL8DwL1xIy1sG/ubKFCOSF4fW4A06EEyz6Vf7lvbp7zjEd4Vp1/NiDem05b6l0/1+
RWmK35roOi3v1SyXdpVZuASsUd4G0mZvPCvTJA5mG7pP5r7FXzzo966S+H1ijoaP7QZsQG/ReVPQ
VlkejEmuVHObjTQUrewzJFUa6eKDIspJKCztmrIxpICi1xIop5opnjUvCM2WxIpeJcOAPggBdlHM
zLtaLI6Ajusz6qODhOX5yuYYZ7Krw/MzOLLWY17+eVMCu/rd/SR0oH5LL+2bh8/Ubi6cKG+9bNB6
2uSTGvXXOO91RH/RqXf03iIbXbJk1PJkS4/1o9SlVogfqkOeslPwpbMEaxktiEfoV0iFb4x5B4B2
36RXGeHCYAOWLSa4COe13ReN5s3RrC4q01R35OKly/Bi9yY5ZZJZg757PGN2AzRblR8zttkF1rFK
TT3KXvO7vDekkPutj1Ku6wcO9l2QY/Ar4PfjlM7QWbGbf6OKWNkaRj1xcm1hue59uY3gn+cK/YfA
kAReIdl1nTaSaL2YqyNTzbHTNHjF3WM+290TgWJEXVfZc0udCQTI7JiykMzaRss4rRNK9pHqfm6l
wwCcY0JzmsboApqoEHrzT8tPZpe5Y9MR3pz9zJde+OiNnl8MYF8u8j/jaVAygXPL7O8c3A9Qtd5O
st5Rnz4Rv0JHyWEXBSmB57WCpr5blEnpHaN+p24xmjAl1+nmUtQEk9imp4AnwFb6HDmOUyejMgDw
0oj/sIDY97BrTdVvdDQvsrUnzq1NdfASGRGqwkV/7RSlyGOTHr+S5ZegeNIxzqTapIjhIILBoR8F
Y8jktU2mdnO30UKuplpoFuk5txq/PSpoR4XVl4/QuDCtAeoGJmvJDpPpxYXZ5szV5tNHDdb8QOqT
CtO3zWEnzjYmr2rHaco+itKhQD8c7ViYrmUPa/r8MQrjAwhjcpe2MrQ1jXTbbn4MubNpuadBWyep
kFRFOIFCOL82qEBVCP9P5Ay99Lr7ne8iV6tFUnt116kRyL+YtsoKYnHM73IFph4nJYM8yZ03JK4w
k7/Ro0JYd4AHbDux6rOZWzHkok93K+sypZ87VOUO0GNP8MkISDZnV+7+YKoKd+ewJCmaP+td5ynw
JwgKEdC8tZXa3hzGMimOAnfIuYcvkjatI/AIb+iKa7h4imt7iidWk+0PMX9sbd+pq0q1ry37ddrn
L8IkPygTHRMtuvjLkpLq7Zl2rpmhf9EftZdwI5D2JvEZHpaYbyC5G4g0LfoO0fjRp7io82bfpCW3
cmmqBaEm8Wpi0BVcbjO3V3huO6an3NMQEChBXA6MPys7vB/Ip0kmc1qtC3BFhOm85+rXrJLf+jEZ
jVUcNcNHTYGu248le8sJZANV46cfjIYpOqnDHTfGlT/g0OXUAGe/0Ul0A++IxiPBlOvwl1QRUXOs
A/9OerYB10Y0tpCVNGYoWwnwtckEfPcc25Lm36grL17IOoDH1xqoLbgfg02TStLF3KRecUr85D/+
XWhDlPPaILQJ+kjgEJGMTy5/HbvNiN5yEr22upB0zQkAuPCUvI6Llpk/VeEbqdNdvFjwRwNdnLDI
+ocagIED/K7JFSgcX/87CULfBuygytanY3mnBpQpZGIBBBklluov3LjHdceCeCC67T79TBZwxXFB
b1Jtp6B6zWJliDNhdGQLHmC8gysbmmJv9tDrL+ef3hWUGyXslSB1GBJ4PG2jg5I2UCA8aIXja72p
6jcO+tEkN94WSejGD/8XeF/wjM+qZKe6O9GmuvJfhFrUY85CH2ZBQMIg56cvs9naV/1KRyaqSSuY
J+mR7Iymd/pxDZJiEGYn5845LarAfKdoebVhGc6yzCCC1He7Pz31Po3EkdzuVbSDHgTdwxiLhYo/
BWLKD2Vo6rYdQvGKuzR3+Ogq6DEFo8hx+43ioiCpjmKZ4EIiBRWBCBCfPr/en5K+oJ8kSHgMN6nB
+1Hyc1dLrj1FB7EO+/Z0d6bJbkf+zLyx+dxS9AXVFCXOffQGz+u4ZT6ZQa7azLlBnUv0oHFbexmr
kEyw6LvdQUqGgeAJaSKX1QpU7oTA2DcCUhtn7JjeLwrqob0QYyjrshRB9wsY4VNF6GuNiCjBF+0f
QCyWK1OAZ4a5EK5dmYzoeGBk2LPiQgy3Xk3g0olUvgfe+c5Z+jtb8eBUvxSLzaTm83hs/tOX3kc6
Gkd5DQak/OZiSUh93CgKvWFdHFCDXdEDaXE8faHM915AFwZitOlQsyLndLJ5ytJBAV+URIPEEpAd
D/qAZHPT8aswGoNBUNr0S7jlgtZgJ2FHxpZno81Xe1e9zmt133aSkP7i8wlnQselk+g2le+kewC6
mHFN++aX4NwZEIj4rx0XdnoZRDUjFjGM12hacXobqQ8UqTMduqYiILJf62KKsA6ECiZJFHEOPnjF
ywFv9nppTRtNJfA2KGYBYxqX2eQidNvDt/vHuGs+RT83GNihDDt6JlP6a0cMNpyNai2EGStPEwg5
lUMUyZ38BUqTfEcun4KIpbI3w8SR1SPxIvpRcT5Nmp7IDo/cJfIOvW/1diLurZHQQx5w5aUAgMWB
dJLKM8bFLHyAL+4L5yfC0eCg4G0HJrV3G1N14tGF5kPpdgtM/wFvvczDG9rfmsYx9TrYf4xLEBwP
nV7pWCQHzlZo9JT4TiTEZJ5Pc902WZlYBlzZgQ8igzWDZmutNRJ80/Am8rT29Ey8jfaMw5Rm8L8q
4+QX8rrSpPjCL5chBrwtHkXQSbQ6myg9wML8JjqTtY8+iG5AgN+pdLiQoP7Qcrwe1kNioDwJofit
VRa/s6yACokoDOdgfaGImpLKolYylTuebDu3Xb3ZB9RFoGwoVoT74ZJ/iaEa3dR5zIFF0Kg5bd7R
kL0IixtaPVSeayr/k1MKIP8YXtPXnzpBC00A7SF2P8J+HgO/YNqnGu8KXm33ENYgFxuVv4eRixbf
zhvbyqDvXMV3fTupBSUwzwj85f0UXHnERJ8VZnA88orL3MCjXsIlgx5O6+p7Oxb+Cl0sGgjxJMjE
s3mQmeOC3mS+hufZAudG+TIltdyEeGqWzCZ9S0wX5oP3/VrrWyxdFu5srj/xQ9HK/gMRYy3OP+8a
0tnct+O0/OKuxox/pg6QKpASmZxrQnVfGmv91B1tiirv/oceeV/9rPLxTbRVTProoxSVClK3aJ+c
Qv56CiZUd+h4avS4rTB7hP2x9QWE8ipCwUycsTZ4FvJqMXGOuaX7CENDPMTBH/OLIXlgmvEOzEHE
idxHVLfdLLjwelcfXzRPNNhd/oBEYm/49K6L6tiUa52n2ZkDX98dTq3meEWWTB3YqtaTZBWNSu4G
paWr5bI46P1NdoFCC+Bz/Yi+/tjVjxnZIDOpWHDBovQh1aTXLaFCsyRikj0gNdKywHB4A19FMeQx
H4EA3ENUmQMC1UWmGNfdtW4pNElkc78FqTtJKS/ltwwc4ddv3zceyyhQv22vQTMRJAnd7/xoKAQM
mMf2iwTd5fjK5ifBW5lLeemXTd3/XsIwwChtYAJV4llhTiJZN9qDOECu0FEgCYYTvPtZETTOeoUS
Od6ZgCKeP/+JjkIiA5f7BomqKOMScxtCN2kk7lFCXlbHTmqemw1X+LhmlhEk4hd7JgpSs9NCYDF2
6gu6+5J5O6LRu1l4iSZcRVYP9S1u8Hkzhl/y5fMjECBByTTg8uO7po4Rc1v0na6O6gGVuT8R6AOu
Hhsw+sUL3z+gYoQC2gtERYxI6+CRZq1x87rAfl3G0xQO6QKCHUAFAbyHoyo0iTXhzdJNxkrUwF5k
QYNId5hszEM2zdD69fpvlHfuwh681z41f+7Tz8/OLX/ggfHg2r0VyXuGiUTZ2jso4BBFpW8ChNp/
sc8zcYP4XYSrhgRgbmkxnLbGhl7UDi5aNu5YbJ4Q3qzLsBmDGKazplkFzmUngBSa4yrFTmPB+GCg
wPCOcgqb58fnJJd/AjlTE+gxJPHVwufwxdJcYjO97wp53xKSEdpT/rbG6BP1bj1XAfOkuTqz/O0X
JYLsxHxFX6BZzjHs063VBF73odaFdRAUZuo8WiEqqArRB+/OJKdPba16Mu5hKaZTtTLeDMPJNepH
HnI1JvZJoDTCQznsvaGrI6elDH2YZxbgwPnzpwxZhHs7XMvWLZ8rCh10bc4tCrKBRh+nXaCh4+ri
L49Sdwjt39wGLDtjjTriz5bMY+G8NKInxQN2cVvnbyFlEBs+uhrD3wpsMALYGw93wCbkKufcs9vZ
+7mlc13hoP9AciiT/6cB6a+vk7Uw1onOFYI38CF86IsHmwI+RUvYPd2jWoRBACvH6g3u9I+gjM72
D1uEHzj3TJn7f/B/TqlnnTIb8YKifznBHu/6fcAk/vQhL45P25YkZt//Q7F18lKm/O52Me10XTp6
hdct6sD8rQusnCSjwpKIYj++fZg6UgObUY8VtG8CoERaBXny80Pvy132f6B9Sa5TQRej52Rj5F4C
74c9j+Rd2BBfIWJzXHLYcjdXLZiwzrmLsTEoY+s711e6aYOuwW6kM8lDmgqEcvogifVdTyChrG8N
unMF4iTV5yZAsTYtTmSfQJB3xEpe0p0TodQipp3XJYE/sLQRpaGW1cSfJBRv7ykc2OeaqCnCZa/3
kT3Pc+1a5FwHzW5XQHWq4WTAMlqtEhIr/vEdP2P4VyVzp+6LEtMp71S1pNOb/3Hg/xlu+GYLR/X6
rRks36ME5Q3VBaAvCy1z/HlFn2XGoH/bki3ytstnwMPSM1hjyM5CjfpcdmIZ3l6Muuq8Q0xO4Ciz
2csd9JaUzdbaczu3d7D2BfA3tSfh6q4+EUSpT/vN+4XPkGMX55xA5cmsIwVwulKDwhduzrKdknmh
7jOZzWNQLICUL0KHH4W7wFtE+NFmI93zUBzWUuB//9qTWdkdlpYChJQWiMEYjgZxKvF7y6fHw2Ae
ESA+JouMLLs6D8q4I3X1RIkcuiXsCv4VEwHvMTFx9U1yNAvldwDfW4WXy00nXWCtvIayQmZpAX8c
KFNBcd5Y2JzJu8MJ+rqT6iQcV9goCLj7yHPLfbXayyGVV59T8rlqHwX77yc2VtZuly75+kNw+ckX
Q2RUG7Y47ciJYUvo2PO3/LyhcGvSGA9nuOsf0hhrHTcc2PvOVTctqB0JMqnhAUqbKjz7RGApiYyi
FrHbw373n5OqZ+zm30/km7AMNdRkkMyJoTvSqucpi2Xh6UrzNdXswRwOTg4NSMQZbv/q0bDRTGP/
wTk/pWAhWDMPHUPEih3j5A8XRP5kCbi9T2dKhNDBG8XgNuPUFplPSR1cP0ClZww3JQFWa3bqb//8
eATCpoHv2LmCtcjrugVJ2ZmotB6TPZHtD0W1IkBvwbpkbEHqQWNxg1SNkRKNuWXwX38MtkMw6VBc
MQaaecj3VyBgYFn0nhyxUMSWBBEPZNH4mfLTOYCkDeR5+3644Mel5eUuu9VppkO50EHggwGMiExM
2EZSFpKkSv6sVc0O0GgH5E0I7/NbQGZzGimnsOmeigX7DskySwGgkJTmNjKDR0dsMvXvTrcRREXF
fX8Ihbk8D0pxLNl/fCmYxjOukpei9SAGOpkYBwoyzQ2oXnUb3XtnljK2BUReUDA/UDdZyd3DQr1T
OvstrMos8X0EfrpnWh7QZ7vK07zVhOUr3f8mwJDXHJtSLT2Jq68hNU8j6v4BIaURwPWfEsFxMD6n
QY0n7CdVG+zSUltrtn1O4yHm441VQWSWfPe9IAbGqyfBnY+vUEAdsp4AeeFIEZSbbzeDFt779FKX
085fgXQr9YdPWOvbMNxM6wfbBukCt5UqWSquYr8+Io9yTHCZHrlcjj+ZIeiolO+ptdVcJDDjOBxW
djPHey7zY9F9q64N347a4WQzw+knGCUkY09h/PCOFYpK1nDboKW5EuKtte1q0zf35I9KpcszjKpL
ms8kDb6uBTRdI55Hb5hpEUEtk7tJ1hqgO5Dr39mMqOkzRHEZmoBDtb+vxaml9gYcVLl+D6Ca9Bjh
aYK7m78+RjAtE1uUgcN44lzLpGpbFAJBElDisrLYYlZUXUzO8TPonzegKnh/S4n4wQVlHDOAiF30
2SFDegxEFFevkghH1iK/Ow4Q/Qp3INxuxtbU34O311h2HwJmBMOF8f78u9yl6JDU5yX6w/h1+BWI
jj9+vh0sdiPl+AwvONhhnCsgcQZvpUs3/ISBWXjt3/94xRS8bcGOPPKrJBUHWbcneknBzTfTSFvQ
Mn9ua3r/dflFTfJPeHLb/hJWe0KDQ/XeQhyAoxxUCSuI8cgnoe9LtgVe7cklR0D6VXcA2fAMs1yn
ML7yBGgwkwMoGqqfeko0QF7vRhSifvSj4aZkPFG65bvVw5ZtpQH+xmerMHYZxWG3uEiOPLQpIJbS
Qcit5rKcePO69e6LDwMD1k8Ls9v9hqmQBIwiqO+DSutyNyMlj/8EGGcFmFKTo6HslbHwS0nKBkgO
1era1SAOrdKBsD5B0cJi9mZl12eIkbwdHzFipH/npmmO9gwaKQJO0cJ0flKHVDjHg3/fmf8y6bZZ
X8pGRFREfxvAbQ+K5t2zC80MszftonhzO6W6IjTmPNCszc2jkhWhPhFJgMv75JO3+EpjaUFPOWDm
esfC7gwDobgE1LHfvrrJm9ghMOZM8wORizqIc1V9nPSsf43q5wDUckvbovU4tt86uW9622khjp0W
nXhXYbk7k2NvAFm/FeWXlObx7CfzV05HvrCA4Q0/nZfXBsvORkUaqsti/nF2xIqBBhWoUYklJIyl
TPmRWuZ4VkZYsQSkOf//TB6Wu1x3waGeXaJhav9kJ+HIv0Zt5kCPadfR5osIS6lshktDUOQ7bQs9
h+2nrfIjIA+ke3PzY2UO3rnM6wVtQbyI9oGwFwMtCXkg9C7zHh4aZzwcPfqka/uI37pMF9y8yG7o
zbkL6eQAb5nAR5s3JOyRd9a+6wlLG9+wtgy7GHTkRFtWUjU8RCtfzTPiWKPFLz8QubgkDN01rAZ1
Lfwb9ix+k8Jkggzcc0w2Xd+8/DxOuO15VhnSRUoWVWtOPqLdakfCyVAty7IZ4eKS7S1XDsoHZvps
6Y50Ksp/c5s7kZFkMtVKyyqvsEH2OQ7tU1ucwu+QEo7N2N+sfobWpfP2d/ic7qlAc4iouSX5i4w6
EoteNSOd2GUphfLXZkxvH+7Q7Tth1z0jxlDJxZVu/9mVs7oZjMrBPh7v1ba6E1eoW3kYLmYTQMVr
bCYaYbbzYsnEHQENQG2WkBdrwdevbJb7A55B4s5dhT7NULz4PGbHFHtO5H3PU/ukPowItaoz7Ixb
LjjeKTghGt5ESdsZzuqefSEYWTeFcobA4X6d6qWkWzpoAI8LtTxWrdIRpEozwA+h4sGO/KLe/+Bd
/QNci9Dl/cs6f+WAREPFmtcJZbreIlmRrDexvgGqjp8ecXpp9YhTk9l5ueyUPFZRPWdHq8cPcZXI
eNuW1Lue8lI0sLBCq/t0C3E/PrEUIUcRzraWK70XlKwFSFrFCAsCLPCYQnHTU0NR2et+XPznN/rh
uEPA6Vj9enB0a74LlK1IBYMVTfXISYdScOYITr7RDHI5CiLSENv6Cj0NaiBDHUQdcsJWaNAMcR0d
+zTfUBNMV2K+OmjSUwyID4g5B0H70Evg8Y1j3EA9ZZ3Y9TrdXWWjG1jwNFBweFXWiRXGubNMLGtH
Smyvh3O8FP5CZmD+d/LroNusv7aYol1SIMn90uo852BhBcbFhlcJoDG6p+jRFHBglx5W6OjnOp16
1TThQL7HrHTKuWlGFRfYObUZnoM604IbfNCMNbq1jzPV8yrLQtCu6EKAlR5qOVpQfaN/0sMi/tqC
ds58P1Olhf3JP7RFS9E3BQRF8FGgGa1c9HYrD0UaiZ6Iui9F+AcORLD/awZAzgcBPywTHCk7fYRG
Bs2ih6n8cYivejJeoEcyOtbsHUpvPewHzOt5sFyWRrTDmQXTrjheJCx+CbnvAKsb6qLR33wB1bFN
fHZMGAIIkxhKtxos8lr7tomreFvevvDvjNjr5rIbyYwiv9549I8v4BaAsRaJf0JK5jYME1YZ8+PX
Nbu00raSaEuCbokPAuRh93cDId5HWXrMkdGb7URgU3cRgGvPQUj7ae4GgTLUbk9INN4usvVbFdeu
OU5XTVmuyCKn/6yHxtmDfT3zIrRC2NF1XDBDQ4oU3J8zmdNmjmpmW7dk8EiP2QvHW85Pp31nNymv
1u9LON3ubPIevXHlXqGyt+rg9s8e9teka0IfM6c+Pr+gTxurgtFVVeNYfDzFhW81RT+HWmWhn5L/
mHR/wATQoj0YwFBnl/xPSTIMGYAQW91qMpxYnuOUuwrdth5gpA4W8O5YRSS8tV2WNofT+bYu8mCt
SwqzAw/C6OaoI/xOoKr31Bs4J67QIEAZ7Zzmde5A5aTGYN4Hk4jmdtDvO2BxN8kYvvH9cRBvZzsl
w5UpzlChb9HdSMRv+wRDo/fW5BkWa3cu4yQFd2g3GLfTNCMHbUdLqA1HOGBZueN96tUQbAhoYQtF
dq80hmUUYo1fr17XbKDoWk1l0FbAfKQ5V7VMk6R+DuQH4id7UdYftGPs7SgGvV0bk9zz8Nf21a4m
Xj0IN5rrhBjIkcB7aa8z9zgEuEOSGwJg3z/KR6YQwkNBCPLOEtP5Xj++YUlA2H8sIG1yViJuODCY
Xny3hCEeyNyGB7Bo/BJt2zMabVkbzMg0lM37mCTRDUOQxK64Psz3nXqXRufAd+nplwMl1jnQy15V
fOGB6X8lOGRLLnYs3iU7JjHRfqkHp5ZgiQU42pJR8PRu2aayDvkMgL17XUqiVd3eRvlcYad3Y/tB
MuvAJFBh8uS1RlazPlCEd3yjO7YGiIeSGs/xhVhplb370ou05i8s8peveRCun3dF4l3Jd/X+D2k5
6N4jsJP53j7AMUx1mhUhifI5n3nTC2kGppRENhc4d3OBAuPN3WGwQP+sYM93up7fyAnD84z9HPXU
vsFtK9SfT1xgMLtayGvXh5iXVfezfa30o8roIxZ5PYeHFnGH/Vc4qU8LA2HEyi1zruWW5DAl0YsM
/w6brTpe4+uM/zASboEg6+ey4cddqiDUMhS8BNmLS44ot9AcwePEKgvQN8NJ+SGWAbnnfz39s5Cz
LLoM4rYnmhwAEEKDrNk9J6t906qnPlW2tHXnOFnAlbfaXs1a1YNczDgKKCpj7yK5W9RLkAVUjYma
bjxv3ol3XhIReX6vT3tpqWnNKlr5YqJh+TagiMK0oaUApbYU3SB06ahXGhMUnf/Gdm4d8vE+sRmg
hl0qHo+LK86xLxYMdttiCn3hWv2ZIl8S/JTXd+aB/wAb0KiTJ55wpvs4wlPIePgNB6Bu2oN+xoWs
hytV4DEQObbkHEYu1/ohwqPUX0sar2xPtYcGjdzhBVIDz4kABx/k1lBDmcqdbi1VpeJSJU21xS0P
qzsKUzPBMxvGxotCm78KcsjX/bQY5lHGiEsphhVNdDjJj1dmDeP2DA18x+t432O0i/Car+IE6qx+
aHtfh5G728rgHRFzJB2GXKlzI65aUolvGNv549fEXepI7Ayu8WOh/wgVS1IUwnFVlFFCMy5UtFP8
xSV1qmS0tLStUiC/py38xqLlbh34JEZj1zFpRWSqD2v0ySBT1z7C2yU8vDlxmavIg4rwuzFUVDYe
eWuXe7AniRjfTkinu0XY1PLqB6KLT16Fn3t5gY1kK9lFzzAHBeVR+8oSKt9Du4lrMEkZoZ9vTjcp
mAM/WCABB4ZjQf+7AW9vk1Z6xP3HAKK0LOJPmCa94KqVYTarENG3lolbj10YxspCx3s2Y9W96dVS
j7nRRe5LY+dfCBSd38k/icqs/NQOXVjRRcTSuNNM631ULY7R2ww4HAEwjTHIJvBlC+orYGkv5bBS
x0jypr9C12Og2E86DYMz3puLh76/eAZCu9w/8TxJHmrwyq3SXydTqXnhUak+p6wwPnulmnEKXkB+
5ZYLUR+8f2tcb3YviU000FucpzEJYnHoOYRIFisgZtHurFYa0hnz1W4D/FYMstiaLM5Nf+1q1kw0
SDG5lEi1iDWy96/1HABSRntFlqyLOOh7CPmYI63rNxDtnZkg0VR/CmBNdkXrCXhBmzL/tWBt2qYa
BVSCHAM3pE0QkFlYXvRK+J3eGF+ZvbKefoN+XPx/IpL5jhCj6FlSPEr5cloV4srKhw54oqHNc2s6
ZtoRTVkbEmSlWOVfKVHOVs3MmZ85ige/+1G1U5WLmPS7XsZhW66jjnGsJZ1JD3JgysyQITjEdKNz
twcfjFrLYLgAmmJ7umNK2u3320f9iAgKn0X++1TMLNhG6BzipOkdEkR7uTyqVj9IV+0wu0FbJv4d
9g8QIPtzrIcPZdWkde2nG6c6UqeNOLNprx4JrSc4xytStjsJeTofe0CyW8B6SB66Bhlz+M1YalaC
1698E3pfn3Ajy7DdSHDhVu59twd0HQN25XfpC6Z04/l+KuTjSN3hBmenyIDwKGSRnGIfFqD0x9cA
urMrhF4Jxus+3pCWrO/YTPWXUE9CsXRi5yRSCidmgj/jf+krNbtXQjWOHCsvimPOwLJWCwBA39HO
sTDNwqUzW1KSJYcO4ynjMg3JnEdazzcsq/1q9V6n5ywH9gAKRphigfswoW3iG4iCrcR19R9FP4K0
kk5q8mUILMc02tS8RBwPNB/NgH0F6jTbv2CmGLiMhTsskfE99j4BbtwUW39XgMRQY5LexFyAVa21
zPA4PuHJCjBOrgSO9OqmYUkFYKIujmTVVhhorFvisH8IKl8w4NBWEDBKdH9MCNPda2GmvYIGErSg
yOluSJMvLYbd4Ey6TkAOORvLCqvTBb5pqSlXa0FZ9wlYMJjhQ0jG17cxdJmbm0cBsTcnlmnh6HcI
kUFwpv2BS6b0btf/rNx0RSbpAfBNwLpMyjAbwb5NiOf2dZ8cHvsrxPYaHnbN7ndWCviJyYdvP+0/
W1X74svdprhqp3pUsBjc51+78DOFJ4x34RdTGTdFzfyPe436Ld3FKuMI6EeM6SvzE/u/KSE3eQRZ
V+kdaV5be2of4vHICYPkx17GXi4s704UXJMrRTHRpsazeMbnnUK6LI9koWZBbL6IFFVaQi49VDdB
noabgOaW8Fxk4JjtcLjBW6lmhNH+45i1xQUHSM45hxCTG+k1UvMwsAs4rUZUwUopUDjV57B1E9qS
XjV7ca1BbUsrUzNPb9IbIG6/SYwsPIffgDJfXvznF2fLLvuGjp+uJAw3ZFY+vBW6DsnzEhbPq433
N1tLhqbjCEn3UbN14J9v+XDxqtQVzoEtK37p6jZjCPXnFKmQmZ8Zg0xgnvznGUR73W4dCUOnVs9+
HKS5j61Q4Av5mGUez6o/YtjLN1pLoTU5QNJRGi2d6YNuOBEd4+TqsCSbOK2RWYHab1H/aIWy8aSW
2pOKd0NO+T55SmW47lgh8YITWuP8vb/sod25N9Fh8j0XtxFmRJ1B8il7KsC9mPj+pEBCreSVt+ie
7G9kJ1VLf4A4IWlbl77Cj4dUhDD6+B3WBnfvAyxH+V1OMAgCQy9JU24obp444nC9NZhEvS49MdiQ
HQHMDR8v6kQ9slfcK/S6UA4pwPPyjNptH1o5Fsrvh1tTJKhdECH5MuTODKX/INb+AOSmiQGW+FEY
Ya8ZhnciXv+iJJCHEFNa2FvpJ/mkFKp6Zvhyh/jBF1sp+LsWxTdz1vL0HNzqRocqBnLGPmFma03k
q/5mGBHI0921BCKlwTC/KSPhlz1hCl35MuXt7km55lc3KMd+/souzDKxgrHpZJN9tDw1SQwCZ6pt
fc1V/8fWsq5BdoJVCCpe1mbTnNolY2WA52kubvvMu6ar86E2GNj8eDWupdb7JMkRCXfPQkuAAeUf
LiSJ0UXLr+qQ/FAcTmzFqChqnLSAuCpIHDsagnxPMvqL2hEOHNEcbrA9/LYt4f2Xxznwvb9j08jm
3Hfz2I+For9kOK2DPpxfZ1YNC002fiJP+R6V9GZ/aYGIQeQ9G50LzOOZYuWJoBskIBhene+/H86Q
WVKrNQcz3vsWrB2d8uRA+xQ/wGw/DxWpgpR0zy6JYX4XzLXo7u3l92uWTCQmdtrwmcYqsl5Q6L90
95wU9GAZDf79h0kOFAYzOVc0vsEGSlI6MGZIVilYMBvEAmblzMbiHmWodX8a1GRFGO+ofWBxFFHl
o9WfuBmN/PS34HPf8VpW0kUwWvWLSaO7Wvwysv6sKuRWkx9j9UdF4+V95GxSqD0X39R9b/ae/vL2
0TobQttmorp2nRui3fHRke9SI++5LF9hh2rKEbcFciuaTeGuYSYZFnKpJW83XnTaoD/vNmJFC+/6
dIz6KpXsdjO3+zcceJfMmvkKyBwD/gzx3NS9lPp+fMFnfemDXw2bmMdstsvG9BEsGAYOVX/yjQfr
arc2Gk4z4WZ5UJQ2t+X4hhFa24wRhKCl7pnRw3NZPk/Kg3fAkRodEusoH6aTE8sEiIZZJfiTvjfY
bXMM867qrDP0iVbKhrdc7yX/30RPFCyxe9DVQVg9BpJhltbWOwMCd8t+wdGzw5tXpAj0lYJdkXoo
tE3ZGgV/2Yl10Jj9/+ZMQ+50Ont8ebfUgS/uSmRO4Vd+x++658yGegzGA8HkmqB9mmDuO8nrjoBt
mYcMVJtD0zXCsEjZTUTT7kwqgBZlSTgucAp0GdODRaIlJwphEHBbWC/RwJb4Z2Bk7hYeil/yr5FP
Dj9Yy+GBjOwSUFus/97KyEhohpYig5X88gLZdhUKONZIp4UGhv6GeoRmrWjJNtYFg2tIfLS/sG8g
1BATRc7gs4s4uN4XiqW0CmAPXdXKf6wKAh5hBaeH0XkXKcYwhKbiz/lpY1IQdxnsmXNvqAeEwAci
9ljxcIkw1b9OIsGvhR+VMYPVDrBh7dAygQnyd8W12nEyWmiMCyBV4cQYYYaKxxdcUJ33+BCRyZqO
5EWey5PsjVwThkljYihw3t/i7MCkPjdilQn5ALYqTLoje3JN3S7i6RxKwRNOZnCQQ4rYTDToHjGH
zrhYqgBI+pxa2aad+CwyGcVKPKv7YLo3/aom7ZJQcv24D/4+QIcvXwfr/U89VJNDgnPATyEpG33L
NZLvS+548X3xYiDohMoE6OTS1zjw1fALjOdS9mJ/ITD/nSJ5bNsD1AZLgVmmbz4xaw5ApZXilpir
tRoaRUZ0ATZ9w92ncV4Z+uj7rxgQCTJdrZQNSlnQMiZlyapK8NbBrToKZE31iDzKSb5g3Z8uuSc6
ZkN8q6NG3cExN4LX+S3VBF5V7Ox21Obo65Rgh+CxR+Vk/wwXGlIzCCLTAI56tFqGVK9LqMYDu4lX
FwBNX0KSyKhs04A1DMXvFN9c/zhuJRnoJsWjMrRKJVDIVmjU2NkeyMLtWlCJ2echunbIsOBIwjGk
cfMECHqGmGMoA6g79de95Gl9e3uI59CppFeA2Con8ICXnqlwZJlAJjPCrsvHCkvvZnkvLgpy7+zP
5BMd2X4ZlYoiU1EZ1ttADn6bMWCiekwjgkj/bX0rmNCRshD6yNW5QVmbebHWgO6OLFWkLouKi4jt
6eBnedPTryz5q59AZ9CbS5neSziSzxwMAj0FWZjthOrapU4UlGtnGCUDCyfJY+En7NqQDwtPiPio
qiIlX98BLDyGWvU7Ge4Vf/1M49uH344a8TVkR2Ld4tayZwwolrHWy5iaJX2+989NpoohD2CeojhG
0zalaalEKHzsI6doIR3RA0SPg7nkXsxZrxcwMToKK52WR5FkBlfB9uCALHYfY3WlJnJx59aFkb1n
C/5+c2uKo2Smt19R4wB76vlg++2betGnMYlb5DDy4u5TotdH5DxBmBXsUdEqsquHXdFYnInwTLUi
DOURDU70AtmlFIjC1aPIkQ/uIirS7KDKAWuNVDsWJs39SDbuMuyQ466ZdcS6K+bTq0XB1HHclBPk
ijWbL4ZdwDekMMZCryXpZ25mutcjCFV3/Upoy7ncGOprRrF5TnEvklDklm6nNcGUoaQ3TfD56Jnn
BNJpB4OMmDEUHnq9WHHAAHRRKMaRz93pCmDdGsw45ko91t1Wxl1D8gaD0jEkynVG2e6l/xEaDlRP
mZPK+blla04V4Dl+IYlPF4tq+AZHBNE28dp8hqPC7bPykCNc9JLsDcxutpIY7C0PVlD+BGN5yFoE
VQiQFqZSttk2LMekGTIl/4VKCm42eC7OYGoTeAhi4Os6JVFWtKE6J59ymqcj4LOTAPlQJJk7QuIq
EiiNi2hFooISG3pdxXntEAN9zSDjsyf6cmRysV+BjVZVjRj0WRuFI1RHhSjKVgHZKWhEESPuH6x3
OeyUPrlIebEr/NVprMrqHrtzgRdGS+468GnoqEd5h7A5000VdxYXWV9ve1m0w4aM2EbYbxIwNJ1N
kEinqK/C4ka/c926FBjFPoWlfcQNophmtzNPqZwXovMb/y5FPf2BPYhl2SUDlqG6OVRPGuMEweMs
TzK1Zeb86CH79UJjx4meRQ2bbFE+otEVnJXZPVDAy0faWOPBEtTklcnVpM4Dwnb2lUS+sBMIr1yu
jsz093RtibsKL6uRbXYra8vSXn0MzKEbvmimwjnpAcxEj7d5iZfy1Noi4nvAe8YlLl0bVEsd4d80
bn6dnt1bOlR1w67Bl7GpbVu7y8Y4z0OfCGMKHAJGwLLv3rl5HmBChquLk9DN1qvbIeig5v0kEQDE
EZYz4Iw8m9oFspjt8ftYDx31yIjrffmhg3yjJMNbi4fWlFrKb9O42z3Tni9xrnXvuYiz/Q51hoKe
fnVn5yP2wbpgP7V5lgA/3Dhgt3Hvmei+VSanjHicu54pS2osEn22s8YP2c0KTJD21BfQ5c1mFidY
6QgCWxbrQNlamP9NaK4ltNxJanRjuIxOLB9Aou+zsH6F9CBuCsMm2Gnw8Vz5C3G49aPiVO2Bn6fY
i0iay881fv2C/Zx1MJxADrxJfDJa/aSqgU1w/obRFWUJ2A+WqrR5IIIoihZa8AXDLH59PBAEx3Wn
oyd68TO/m1WIrGQX2lOx1CPkt5dZAVWDs6pgm1iIf3ssl8T2rhZ4joOiNMdWPiyuel/+CaacYUJi
FvsFjl2xGPk6Kth8ewAuWEE7LMPoHjztMfrQV4HUQpNAApwUsNopfmvqoPf6bsvjU9cBKKIXe4Na
0+U0Gs2fb3tTjmSbejD4noDnjamesFGXkRNi7XvZlQUyJL5zSZDnl+A/g3MrAIzzY9lIdEvkw4Hn
peDuEkfcV/PhzPwpn15DksIgtAswLuAcDFmCX9HDiwc0xqQj6ZE9cYuHsRAfhsSRZCtA+j6JL5Mi
NAeCAoW3awJ9vtAHt6iXhJLhKkPU3VdkWYipPNbrY9gGKZ1kNvQyRHkhq8SCsIKaDmLm4846P/EL
+litlDmi4ZQhVCNWQdF/pQtZQ2dJVX+rGUj+IGz9TnHR16Sz73kppBFWCOUld4WASnvi2GI3HsAm
xCGOqByXowt1zSYQDjub4LCectCVGNVxzakb49V7In32FliLXpvMyc0sVdJf9gv6LQSjIcKPMD42
H3s3bMe7Cgl5xQa+C+RKo8yBxV3/2gUH9PkDTLmO0CHgdy4bpQTQv059gSAhOFhoALE+/52c5ISv
gSblQ2MZIJiWRN2BTJ/ReMiJ4VKxMTbD6zkyXBqf1RbGJtfqbZKFTvYKRl3416KiUSwfsySryZ2+
hzpNt1nGr7YFD2PRRrtyhRebaFQDaqhzWy+tOXqp3lLfRl8EsRgksVDZZuKFeFT1TgWR78kUAhUP
dyebKu/cYo1asvwlPKaIrhrXdaZTKJHZb4jZih658ZxbRg+Ls9kGZ34b3qYrtMDK6+KAIXMIpzE/
2Ss4Ju4jr65PME3u4lEMJpQT0XnfIY9bFyTx8P7neAiWFYM0GyuBj8EZarzZ9S5dCXYC6WAEritj
20Z01A2kz8T5lQQ5JqBLCj6PrYan7Nel3gyXv9Xub/rfynkPPs63/3xnP4Xej5aBRFw9AphMjUDO
jEBL9R7lgnAbC3BwPr1C6C4Zb4uOUnq7LgTz+cSAAQ1O7mqahpz521u4mNzDqMra7cTInePOnPnx
jQEZGk7BwAbRrkA+yVR22+J49WdLcVhxeWKf3waRnhonGbp0KDKFfZAIW4qyMP9fmU2/fE3W6y/5
I7FWp+EhyT7ZOdH420dpxeheKX7dOZ4XzTw73l0WCCOdMabuw4K2iHQ2t/a24pH2XBtMw/zbLQj4
7Ykq2ceXHWDYYcfYCkge1iIjafzB7ZDSujc7r4vfubtKx+SFLBT+S6eGA65J5j1z3j7e2n4mKhT6
X7ilAp4sAjL/FXJSE/VSpvdGiIvaUsPzxxYL1rzffKfeH4fFnLsILRaUzsA5tHpSLRFjDifmii+T
7j5Fh0N+znlm+oXyndt3Jyk9S51I4POsU+e+Lvnml9pfvfZq83rmDJay6vtxuHpxX+gbQFwLGPHP
sceTQ6+dzYd+T8V3YwHTCpLdS6ghfP0zBpGYSf5H5v1R+uQyuFw9/zqkRSneJ8sttcqtmg8rVg8Q
eRfTRY1tgwGnmYYqpuVeAE24bCk0HepPQXNfKfEnAlw7NK4BTY6q3VpGQbFHKs732lTEVUefTKty
aS2+6gin9Kc5kdsD9zV2DUJXAJIrXQu93AXlFWSbiBXJCRDsCpioDdplFVWWmxJ70g9c6bSwZkWV
gneOkDEh+Tu7mnkyFs+99gWXhsdkqRGZEP2mhREGqk2eeAS7bcELc1AhT5qixCXMSiQS0wmp1y5j
ZYM7PdFtgaZ++Eln76boYFZH2kHewK+mTmzUHOAmDz2H75gJIm1O5z35KbG26S4xngqKGT1yxYDO
yqK1zPlbHOdLJbAwZcvQadItwej+9z6Dxlpfhc1wpPN4UhyatA6eofXbgzJN8cguA2ovByS0edaq
+VgdIw2YRtR33jQFTlp/YZ2YdHMXUqd0sx7Rj1rJo520MiRvCkJv8iN49nxzuVmlDXnxwSqEck3z
E/zgB9yMjap6rjb0+3KNbWY3rhqkTIUeVj56ssfN48sX60mLSWSIKvBbck2w70uBQKxgPHtzQCdz
xMGg0LwjN4JNPOKJdaVsbJtnMY/RJMYR6n0c9/wW5lmnq9yBpist19Wmu/MaQIGI74JoPKdnnwjA
+slUEOelSw3bqpgk6jQyrzTEDYATtA07ngkEYjgqA0GkH9cW5ruhXJ+SFd5sj+C3to7KR1U6Tonw
UjucqsRjInNpSjTBNnmTzc0nQ4uoVP3IPNX57/kWhN4Q3masGV08c9zufEz/l/BTrjuSP/Wldd3I
rZg+uiaj0qU9hJIHs3g4jF44FKJuqVOSO9VECSQO79ZS1uOW0zGkYx4rUrVSFpo7HBcX6SIPVqr3
ijHPhIGFId2KaJaJ/V+neiZwNomoXe+k9KRLwxSW5DNeiRRmblKbLMlXaK7eDmlTO9ZrKT5PbNui
4GCU9JOpQ2t8N/0kEYfMoazUChy1UlHgOO1CEDH9WQ+RiX3xHeqlzEmKOEB4XxvNfqUXf1EuvuZA
AEYP34+71xPtsmLXMh6KIbuJtQ4iMIBQ+rfMcHMHx9YetiZ9F2JSZoQ31a92lgf0g/md0/PGnLWk
g9hjvU8Naro1iilTM4J008T/Nz/n0GXKG0eN7ceVcs3wqYpTN8Da8iWvENsxZbBeAyYSM4OkCxJ8
VhOOIP/AjNoU2sFU+CQcX4hb2Yoq0Zm3TStSAiIbhD8hWboBY00Hvd8OYOE9RnpzjHGYV4FzXXQw
qnNrw/0KCD8tBLzs9vikbHqebWpFsMzNHJuA92X3ZYHBKz+ajYgBNfn3PsNFFIg+n94xcSLIU985
+oyEJtqSD6NsatfQSkY/p/JpoehJ4LPSMwW9DOhh7497znaWAhF/zcfbY/eHINb4IXzyklzv8hgX
uV/bGYWf43wAnsqCGlKbXekUGHDPJY5WY8zVicEGm/TpOMYlbTOgY9jBt93i3BRCRFggXTmNXY52
zRMaUG1X8H1rk4tL+5uTvqg7vtARlecbcTKgJNIMqZI13Gfz7sTUjZv6lQvEXCaG7dpL/OGYPDP7
G+h86Tt9GSrCM9gF1afnfnNR9R2GlXPgYqOM+OGVbIFLNHEgo+AqZ6jPa4mhxew6I4xR4VIIGDrZ
qSP71vxEUR2v/6mGLCXgbu0Mqu/ihgLnXFdpiRNbqUV91NvwVgdAuyFMYyb4qAflTlQks7xB//us
JuxE8x9nB9/6O6EvkyRqlNj3OQJOxS9VVppaY/UpLyDH/0xgOgEsM4mqCS/NTJJ1hEv7gbsIuzUy
kkg9CpFJNumRiyaKFTIEBOxtZq4T5/Pj9d7eI2IaA4yJCxKb6T7RfjyDEmhgm5SGouLnuB8LlLCp
ZS4sddVUkMiFNMI/DSUXbH8VgIl2mtcsDEsGfzaCJ3yVsgg8MZ2uYHTuxyyiFtwlCHljx/z9/EuG
o7LLzjzMDWZthfwajqpkbxxJAIb7N459OtrC68qm6GLlc+tgBh2hbvhIiB/PXNQfCQVRCpPZcYq8
2WO/G1zNVRYLKfcxBjxhHP6u+dvYESrdr+vxN8WBME91RfCCOZqTVmadEHUEoUDLcGW5cQS2gshn
SwMUBsUZfOQ0wkEky0kylg5qzjHURn5geYAVry1w5ABjoF3Ui4nReG7LAY7P93c8evMRoUs8dEcT
nsZjJvUGkikcGuaJS0xz3iv57IWvUVLq414HMsdj7JN3YIAQJedKfn9eWrI44gDXph2sFvvaWC6D
2oRSZKwPgJZlJVexHFKJft5vr6IVvsm/m7KzJobCgEb2cMw6pEg9TN2aO+XL+f7CO1lJcWFOEs20
UPuNzhuKDC8EioG7oMrPNy+4frCnrjTchzj4+cLS4QeK6VoL0F4tSNwkq3Pkged0aaFTrv03DhrB
DSbg5bWqKnyUQNLNd4SgDv3ITO9gEU0z7/tefhyIs+PTHLHZELYvji3zJxH5zBONeSesYhVffZnd
Li8HWZ6RNE4WmodZIayakWa4HaUmi/EZ7uu3AkWjsehDQzyyGGAhjxpEzRf1hUiWj4EFpaoKYGaM
r5TqBfQxdYkBAeJUjbXShN0A8O46/AzqBfp2RfPt5m0t7X0cT7SNm6VplyKv/LHHNbd49gMjh5Fd
3o6mSC7hjjw6VkQY9gaZqI0GsPosgguYxujKB2jF8vqRpo47C+Es6dI+IfCXWuFng4pXg56uHep1
8jI0ZJZPdlnWwKUCP6U1HQegkK1e8ykcJ7whd3Ov0jpd2caUVquguHnpB8CbALBLI5E18fivTvif
lfN+fgFBuUdoxC/Bi3Zo/ShwwDtRvaRwgkX5zk2X5pum9zdsdRE8kBtWpfBngaE3CxFynSN3qVP3
YN3mlAhy/Xk93prFFeb1LBcvqvLK8AGkMoSKvCB7eWj7fkjI4Dz2GWCijjIH4mbOi5nDWSJKHtRk
LASzjGWjJ+v0By+Ke7TAO2lMqFR2E1moFU/RBE6YfJgmFrc35dqLqSNtt2QbkXllBpDF9eiXxsAk
YkSIXR8Abcg7nmDGto/JukXETGIZTU4L6qSSVbd2G1Da94QtzwQb+Qe/yUeEGGx3/2YINaB2BgUY
NDvVnY/VzkPqGFgk2A/iNkBl7qwEG6TkWxqCrb+vs7nN+DmuSauuZCfwjY0w3kmZZ4Q5tOD9uFwq
ahpsQNS6lIfbJG0KzDzEwr4StpDCg8WHKXpTfR2YfYbpCaEbcD8MDD3mDXZo0t+oxJ8SDFS/qyKM
D6uRTIDlRdAFK3U7KS7tzHzpWij+fRHjoDQo+gNocgCuQRB5FRQ6hKq79yXTn4iI14SXMFjZHcm/
7wI6E5Mn212bFTR1SqfrtFtpD4jXJ9V9nnzs/wIj7hU3NYz8oZdp3gxjsQQXrj8jDuVbcVTZQm8a
ntFRwV8rHlruclT1zSmC9VjEJ4KtrhIexOtVqseb8bonPT+unrR+UfI//c9B2ltsRB2COgW+3OpX
e/LUDyLDL6t7990c8GqYIcdXZj44OjWX6mIELPJiZ7eQEW5vxJTX7LLIwpM8dfC+WebfZvpGX9hp
Hbq4w8rS9BFtpAaCjLxq7gw4VftaBn2R23bHqXRyoxOfJvLq8e5xzWjMnFn8XckoatfvLQlYEjTj
pwkPSslIkogt3RN2KUVmhQ8jXD45UhpctmFSViZEsuuu2+aLtMn7dEXJs/A6+NtfeUzRGv2Hx0bw
cIAgpFQ01SKLGAFBrmaL0tkxa/qQR5FFgLOmYgY0dR7L7KpWq6C+34zXgyv3lV+kclBLNhjl5ueH
SjDz8MeT7Yc8nCtn8E10L3/pcUKxOmRFaKb7V299HmXc3LdDpv4FMK9blViW8OJPDVZCEB83F5X+
e069cMnvOtiN/NHgjf9ZmKqZDFRBsEHrr0Q1bunYZcdRLEm27Svbbqpa4JHW31Fm6tZCKsgN0Yy0
3SBwUMV/TL3deJ4Rfu/qeHDatq0BYE/FkZYHZAiZcqEdiXYFMcHM+SD9s7u47dDu07jgfWNa5saQ
tWoTpFi//6D4uVWWdzWkj8h9WTeD9M/sBkypUzUSQaAxX+fqJjdQ4HXg4gQPGIRyUMyakH2BgWG3
McCRjiImGNedYsY9Gy4fLBfxDxTbmgHT7HthxuXzdLhFCY1Dwye9ULQ2hcHH35c56nUl1Q3iEH3+
ZMxoHLmorBuHkYlSyWNCMq05ikFlNIcXHv4CEVopmFoLEq3ae+KgcwLAYTrRd3LU596O8/tqDfpr
Z2H1sTRamofL6HuV4kSzW4rLhOMB8WS2H/z8p88jw4dvmquSBzkWFTOlSodsBEpoTuQjAuk3ve77
VYSrUQeaMCPwBc2TaKQ6nE65PCIWLiscWS6QPyFZjxWJfmUi+Qlv0X4T68WRSWPr6y9ClGSQeZ6K
/MaIXlKdaVNhwPK6TwQRn9ylfLInKySgwobnWze8BAOpjQ+SuyW9i3s4ozC9KInr25xdCZUep8yi
XbvalwFjVt3cqovCkMfrctkzmQrzhtIPkjDyeJ7ONEyKkWay+gLfV3d0ia0GGUd7BWyuPiX8KpAp
nyHcfLxr4TuOKcBcLSN71XofsvFk72aEJLeNVzpvgq/Zl+txxzbsxkgWWaTC8M4doNsbDj+MAdgY
qva1FwsUF3Mb7zvuFAFBF+So8JSvFLs87BHvsjv16yOAIOHC+14lmpP7rnghG4B+5GAGFeWw5L40
6wFybpzF9sfnT7wTXQTl3H+6KBNj9HjmVF4Z9S8gZJSD9msGhrwGdNoVVvbe37C/lv4OOBX65J5r
XkYFjR8rBWdmc9OGtVoqif+2D+DDIG4OGi7YXf0rOwuXb3oqxGWhrmlBUt/VwYUZ42k6/4M2LFSU
NozvdGO+KWO4t8z+ZR4XWs5vX+K0uz9KoqmQDd9o8nD22Zl4Iu1phfLC7IIiDF8n6GedKIFhIoqd
g0BpHg3nYyFbLmvGL7XzHOpjAOB0/c8LtsunoinnwfA/KO2ncAjzhQdbSlgHiL44taWq8u/SBTeU
y+FVJnL39Z71HniKE7wM8mqDoz/8O5Nqdmv1fQRnlt7jEOAPIC8XPsYPbjD6EnFWkKOgEx1Hrcig
9B7sadSQsugfHbKIpDTFMU51zcEcGvtPy2aLJfMZKDFbr+rjJo0vdlxea7JKWF7vex2g39LfirQi
FasUrkjiqo2w0dCwDoKvernYU7C8Wxhn+jDjMiVeHh75xNdbaGgb0g7eaEXiZKp9/86zxd+XN/OM
EDwRJ6dwZnTOpNXURxIRjW0zwI2/soOuBqFb2ztgm7JEYRfgmIdy3max4wajYyIA0ET+kZd7mfFY
CwDeL7cToh/8fbPDoT+lxCz1z2nZuHREj/F9wMb8i51H4veUgtd7xWAqMeFnjIk8CduKcc9Oz1iO
1Tu4pInxHzHNb/bRgTG88Sadly3Xv9y9rOPtYYWz0EJRXh5lokaFCyaIpf+CcNKHRslrCvQgavd9
ml7UpIjTXupRGAj19xfFtTsemi9mL2z6GYnWY818dSVmnpkNfzwoHT4L93L7qCn/wRyeAnZzKdCk
aIqZ586EnB/9Qc0nzrLYxhHpiyVwfD4iA31r4TQLGstGQ3stLuFS1W9Z7hb7CzgKqyiFPBOGKeSj
HKt09Qu9ud6rJnv2dqzFz2uvT5mQ+i7QmCRuB2gKO1zstJlcxHZ4rW0H5xqqlUzYiZP8lf9iOztu
fyaFcGW2JB8Jn3wCktHIYUrm5faPDjBN7S4EV1OnppVS1BBBX8JeOYbLNVwl4HMo7QvLNxGPwtxU
tHrxzHb7BrlMzxZdt0A3vmR7nFOGcsjyfcLD30cadrNeam3v7UkrUrjUzHyUmyzmh354JSq+yUUp
jeEGxSGyNqmPUgmRpne+kuM3A2TUhXNcF2ws65JeHDCkxW67NvgFYIU+bS6o2aRZU20T8J/9iI/R
fIFgQ2V/FgJZ4jpKZh7DhGy83rzQTE/A0Y2JIL8pBSmvO5Y6PG6OTf8a+/hmnb0Itzi+C/6yJK9n
T2LxdYutA+U8g0iyScrkGsPFnMlM9DssbLAEb+IwLzJnoR3SgS77R8UAbFnbnxUE/fgZ4DlfFHMV
R1KFy5VLUkLqVlz36xJkvh5Oi609BfSFQBsNgkA2c5jSr8wJHxlJisC7mh4Pjv2emMkaiWAYdtUB
7ZOkWPWWz3PU8ApD/kzq8QsjqpoVq4nk4R/Ka6RTZXuFqmFogSiFyFmzBnSbKesTRCZFujnO9xnS
SCu3HVW9Jaxh0pVwxwN5/DxN2/WDoXNcQSKljErfBcu+ufH5HOzrQ9F/Z8/lQFEiDo9Md8f7OKCW
slZS3QXLdclN28p1S7avYx5LysDUjNLl5ICC71xZJznGwX/Vb0wwjZjYo9uOxOETmWMf8N+0Qh4B
wo2fdC4AFLAItKv4kbjCNrSZ44jb3/t+LhgWljttJLaNUGdkwcnvZJDvle8qilGXqI/EcBdBncV9
yFgFIXbckwOvNNoEF1WTB23lBmCB+VOPi0abD6ijQhcA/SefKUhy00vDn5PA0yC5XKLIU7LyH+cs
VZgvGNgzHsjBuck2HPEeyFGfR01/y7qTq3+D0flUbJlGPEaNJxrQLJPV5MwemwMfDLJZ9lmO+UFl
k/FkYEv7Qj5q+e/I2gBcK3xqi5gRbye/1FoEM1lErrIHXr2MgHqB4eqk8D5suc7YxTqfXxJVRT4g
KsoFACBRgm1VEqJESUHbT/ZYsLVgstzCR1k1MhsOhXe9ud1lkp8F+Z+HtdNzTuzhms3RTv27Vqij
1bJOYQBXI987IKx46tgNGQf8HglyxIEBkmcDX5wKLampmJ5niNQWx4GIt9pQe7c51LOmqBrX+VFZ
KJKgAcwJM60WsEhV3zNOOOZ4+cEDzQmyIsUWr0NUr5BAGLC9blzdOaIDsl1AhlrJ4ll2KK5VBWS8
2trYVRocgsj8LwSAmNdNFo9n8jsIwdL9q02vK6ahSaXWsHAr3IdJayg+OI4lLpgA3pRh3UB+KjiN
QXVB7Huy/ihFFR3mbF+LGVl0Yfgx+N+pwICDdpZUZzMmdXgmpfnQ8Yl8l2YVJY6hTtPeDBuAZmPL
TVUmRfaOZS4Vea168mdpGdGMI2RnxbaWPeZHLGkeQ46pZaSL2gs7PbSq+vsRjHVpGe4yGoP8MohU
hd7BoDUEC+6BI444AH31MxP/AAVZcN8/PqT1ZL8a+c1/79F7EDVg678t8TPoQrqxszTzyy1mxFKO
TjwD5zx3BgA2xrUF2K+aR41huYRlgRAH9KlQ/l9IFUqwgxx9K4jjCYFyp4A2c0iiybV8XiIrSttI
d0Hesxwl1NffBj+Okzof+3YvpNch6xqlNrZwJZd5AEVLGwaOTTl6s92TlTktqjZORI8NPxN+B+Wq
UimaV/MFePBmyHxX3T8+z9r47uk6egiATTM63aNzIkBysP3d+brKjHIWcw9FLuQxR2GlS9uqBn78
kVm/G6+yMH/ghacOKWq6R6PtuelbvkNMfcjs19gkLK5qavI2fuTbGHWklyVcNsY9TFAbUM+6qaSM
dXopPRVw2MiYE+bD9w9NAb0bLoOOs0X5fmIOyIVlC+pcpFZL5DMXcURsf2k/bIK+6BhxCZ62IzAI
p88hr1YdPaVp5OQfh4bpE7f3VY6AJMTUHZ8hUgL/d5CuXKqBdVIJINRIJRaZJdHhTS2MVqcZDxb8
e5MfY/9oi3tw9+kF6JrkmzY1fql49mbDB/fmU1b2nf3R6cgG1jZovvOiEfykaYk9xj9g9AvZFck5
pixBo3X79aYHTGRB37EgOHD6AGJq/Mx9tUQfcdYttrM80I2jgYkze+gzTxckVP0feQPqqSbdYLY0
ofuEzvPE3E2T16ye/DIwHc+XU2CTCpN7LKBygJdp4O+/QeBiLY9Kwahn7RC+l5LC/pgE4NWEFyxy
+k7Hkg4sx8iz8fkiwRYyBvJCA8j7PdW3yqtSJO1I/nNJvvAoBrP7qObb+YCCD0oHP8M2WSFkkoIW
AmB8oIufQ3k57nWqWBiN0faLIUyuZE2qgvEcIZ0cXrUELLnJeb4xjVUbbztVRrPqXpiPuj7++Em1
CvuFU+x8I4T+hNS8ugGcH7y3ofoDX1unXr3LksOBQOefGoYepELdmbluRjJ9YX0eSKma1ykinX5I
7mILbtuImfPYgFctaI9pSsbU5B1VaFCKN/8aVbCpxgAI9kZjkkKCqm+B5qa/8QaAjGkxCs6TB1qa
I4lmM2rB5usbApZWKwOTcfcegDHvlJ9r/0klMuP1BiZ+MF2BDdpjkhmAX8+/TFqM07bbOwQt+YA7
6qngFYhRh8GKoqE9PYeYg158JqOqaaKPCr17gvl71DxjrjsA1pRAaNJwP7zY4ch6YMzHYENNXg0M
ERNQQYqBS7onrkyj3zWucAftZcbXP6Z3vOUQEup7/Y9lJtB13Jq9VbWULRUn2JeCdwWddqCTyovX
88SA81deK2gCKDOkVIPcsK68aDmG8uXoZgQeirZnzDbOBeAfUF94zxIgQpxczNANzpq7RnI7C9R4
y/Xr0NnEhpYauNyhxoNL+uCJWEyqEeK/jeLS6f9PQZKnFO+hEeRwyamoGnzj+JVlm1zEh+WGgFE/
0RLMmfvOY7l3eJOCoCU2cFyzt6xjrcMRDXqjdpGz4M2xuQg/IjBwmZmHjF0hLFvwG3Ts8ZP/JCSo
zjEfcZT9TWnyNeEKevSMRUALAJTKgMuaweOETsivTSGnfP4OFkVGD1NFq4rN3HxbjtUzSkKPYbcE
do0GE1bXVpqw8bQYl7vFjvQ5luPvPcH1pkCq3TSiP55YoWFv5baTv8y1KtIChXikkIGJdnKErrPN
dwgk1Z+7Qi60J1Co9dR8GMHQSBY0zF8MU/6/lbAh83Lilw/oTndwk3NV0n8XjgvTABVWs2iwDnQd
BKLmF1LSrbeuUBOtZubVaHX+5s2UXGLIkR5Twe8/FqTBuJ5DcVXPANlru0gN6bQuhMobivmw00l9
GAnLmcVYkkGoN5uc4ZP9k0KoCOYJLg8d/pGOG+Q/WHtwWX6Yqb/kvoK4qu1/+i4pwl6zVYdsR5vn
xR7wjPCcCK9uXCgbpDPrhFTtjzuDJWOqravPlVsfuodf7uoRXl27fa+i/G/C5owBhhEWqTrwwvVk
niWkKvUo2s/SI2ZhxnUEptLuZ3pYFTOfWegZJYENwE3nVOIyjYB+FZ3BtWSbCr5Z+xzIb+Yf3nDD
L/pMi8T8TYqFIF+q3oKTl71nczrNf0HthW+q7CFdP45vMc0AEeZw0hyKncQh5XnbdqRUNTMOscYQ
0/O9qNuLKUoybyCbipe6PPChzLhkn1PYrfVW/DWPcf+6yRhwnOQVdJtUYPQWI8IT9UcUjsZ6IJYQ
bXyAxvEkdP+i1Wo+nYJCWhI7PVrJv1CkHMM0fbvphxZmTFp1XPFH37dMPWPjQY32TrSV9aeNjt+o
WTM1QcPRIhXQ/0lEEak7X0Yw+hlMf7OQuqYreclL6BDUZPcONicjrhbVlAeHyi+8d3AHY2OKGJ41
8bEJ5gQO3PvLIQPlxjLu583jzKdmnjWcwXkq5/oE0M+/evtmB1UVyifSusLo31EV5hwr7OoM8/t2
hwLp1E2zIz+mAr7krSftokTrMB31h8Cesq67iKqS8dR8WPSmx5DUcxTlGaqPDJtUR6xU2pBTEahB
HZqPop7I/RUgYB33To70bPtZnuvAYbSzhBAKpwCeWVhebe2MKm6wRXRs3Lnh960XvjRn/MAM0A4f
CL3sz8kaCTuQk8Ifxo9hLRYb7F2Qz1VVWel2tRt8UDBTD5ZAXmPuWGon0OcHQ+1iv72ryko4A4mW
frtDMMZTbVCJAzO3C+ohQMHD/pSJIublnSmhQ+FFAfa39GPB4W1B5uwMUI+1eFT9YgujjoLa1v/p
rsfyIN1IEm0iK9gddGTGoYGR4/wLZfIxaqKU+b5zEiRwnokLUMKRA0vzMx3SdKH+N5UObDWqO5Ha
ucBn2tJ6A1yXNb9sOLUdRirtmNWHwBXucMELJWuABKk+r6lgz2qR4yZNXlTrgn2iGbq5Kh3c/BuE
Dn3nz14Dzp8hvGCw6D0AcPQwGjCUnDdcjqc8JE0ry8f9n6txNuMJBCjwuRjevBHZAqOgQB4otizv
noHim3eqKaA6MhaG7C39avf2arJGlfU/27yTCyMsOQKgI+cRlMXx0VBEx8kLWTCeMB2q7xepNHAm
on3q0NyocGxydVJe3Z83TXkNO8M++UymUAEF1gRz3YfLiBD+Z+XHmDAP7USG0acy0Sj6kGqFE1dx
tc+zGPzsCxtJs6On5tBxAKFAFa7D57aKv/9/qh6p2R7O6SwH1Wt+J6wOEtHPGRyTiEE00pHfGhQA
w3tsdDpUTyFkSzNM8QyFK/trxORym2rnqAi2oFFod/mdkpgOLgiQoPSZp/P+LE5mfGlgQtCpNHZA
iAY8kLkSKcBXQBFZNoM3rMJo79cJNbqOe4GSpb6V0y5+NjH899bCT4ECXy3q3PEeHYrMSLoHLB7O
0Jz57mbdvz8w6y/8r9f73vfc6Nnf+7zHPDR2p/Tf7SeZbzF+DYUDrNc4/+adNlLV8YweD3LWd0LS
onbQZWMgGnod9Ktig3f/PQGHxL+jGajVkjTaD6eUleKmgU2h3jtEnTkpY7x9xKNf15YlQhLdwCg8
KaGO4ysh+kr+WIMMh3jOUSBQVnpozOde/5GgfKc8joTGUhhWnDMMHqIxD3gZXJlGYiacATCASb5W
vBtZr6Gmyu1LdIyZXYloMqeasZL4Gi6r1oxzTcmSXieJ0UEtFkzyADJ31bqZIajgcqJa2+Bu0Xi1
QjfAHWwAI1lc/rakC7sFWnsWu8lq3H2WRmYEIhHay53c0HqQQkx/MSJMAbzbbZ5m3e7nGdVvj62w
iSIZLdEX9XdFUNmOYwnHHdRQinpeIcCnr3RR5Uf1Qty8PAPj1wxWGGdNheWcGXAPyzS9R0qXXmJh
acvu3H4w1Lw05Mh2ffKWDRpQviKt8An9TmWNF8uJB3zxVDLFa7ANu32W9JGmCAAisLQ83tpliqys
Y2TVTyfJwAqRDLhghcY6had9fu3shDTk9eQL6JF6ROhH7g73JziLrOwR11J2Hkd15tS3JnLrbOpi
jlFvVvqMXTXynuG/A7dbKplGK3cLBoywQVlpfDknKV9gT8IcEk2rJBQ8bYSOXgrecBEbRjHWBaA8
GAVftJTlkiy9b+rD2+fuKp325CGoKfLnU2Bk5+F6IOHv/EENCq56OPwfd7TLkBXQDc8SkUl0AMaU
cb3r50gde1WWQPPRYnYE7RieBdGzzOFnz92QM9fyx85UFuibwUtaEcVbkQkpI6xu7PBlKon99Ak9
JC/7uMXCS3hvCnD5zu7iHmSzFkQkmmtsziW1UuqhhTbJt1H+Leo5EFhlq+XNWmu7zszLK0xxihpD
EiwAzhNDq4Ko4z40RMs4nRoHY/+gSONaqk03ano4ExGyCFj/o8b+/ijifJeSq9I+nnBgCAw3Wuzy
7rOXyrjj1k86kNrXS5EHbCxq+MfacB9/lIgHnWesjDqbb7NngMsip2ievzWcb/p1w0f+P/afHEqU
B9rNi5O9BOcJ810/Qeef1+khh8m9wWaixMhTd8OP5AZaUS3hGJAvxlG/N9pBgi7tt06k96UIAnL4
VtdLyw0f2Au6bdtkcWUav82G5pdAbRiSnNWTjZ9ZF6x06+6iDULKLbl5rtT98Jfrt56aprZr60K1
wPJ5j2G4bX2e5Abm7gS/s2wgumbLzZcGSJdTUJpzxfr1aHe9HIkSQ3JfRrgfZevVVSdlcK4NxTEZ
pHoi2dVFL6Xh4fPQy4sCxxvZnS4OuCKETxSUs5KRa3hdXOXseDvoXc+RY1/j7SVhq+iLm9mBVbri
UU1sp3ETerbLHqbNOe5vx1Nj3wbC2lAyMyzVdgPeos80sNQtuL+XCNHozeITlThgHyM8F21PEN4D
Uv+90NBvraNDCCwxUzp46JRhYpnNobf9zA1jpgRVAwvPwB7hBDYsicB2mCucrOITL2NoAq3EVQ+R
9cVeMGk0lxfLvkJvLE8bxM9//Z4TdtiT9Cb142gbHFJ9giRh1oaBgQ2OohcE2MP2fT5+GT7rj7Uy
q4EZeoJcdUnbNb/5Hsce3B3tiEwpILbqhIRRHo2xuTjpqStaUir/1t6D8r4Z370YaHwstVvC1/g8
nWDjowoCdWbaDe9FdA9LQKuWdWQ7CYMGbTBEyKnGjnhAU1vrVF0Gq6s5mHk9vqN4x+PcReZ+n1dA
O1o1rTf5uHqgj1xxVQ5HkBesVEc/xgn2FCirW/SiqK+/+OXO1ES6YE/DH37hgQ2a3fmamBTfudG2
jOy0fVEpF8GlMRTG6nqj6SNzLVRZRYD35ILxOk3N66idUuuB5J14iQXjg/AG6FWkATRN8IjdpEk+
84fCqS7IhKVOhHTIHRLxK2tny8g66iO2xE1y5/G1BuCrfX7R849BRy5bYVbAZ4uIIeDdmPopQHHY
cAZqUGjwFdca8E95/DRP2zT2Hn9yv0ru5yblAHMyFo3l3Q9aEoG3r4ns3mOHZuhuRn/ZGypE84WI
MRX6hq5bpnV0cPvzQNMUXXK90UWJM2jFhY2fpV/9RFlQ/knmg+YFuQGZQ0Y1s773vphZ2VObFZnI
EiNZBWn8shrOYWa5R5RhoW5F67nQ0JQp25//h+8X5cAMRWOfL/gdJnQv2TltzhusUpGlE7S1s/rd
uRdO414m/rNQ6HD6E/2eXyXl77U0yZPk22jCuAxOOudw4eKE/LKTfCagqKIPiCBK1+d+bMV/GesY
XX3p+maSn8AJsmIJntjggE7jgx7GO47F6OrDlDwbdXe1Ib5QUEJ2p/5h1iZ7R2RKcZImFubdD9lQ
tuJFQjkd/FKiSkUpozbxKod+3SSOq9rVZjCow/++Y6HxJgFGYfqOYNxW5+ztvvtzJ11WHQSA3obx
BPUxhXlLXIBIyT1Ku5ogoguN94UEIG+XPccSZBGQCB+BrnYMwvpvXrleGDsJheVV6oMuCTscWV4B
Pm5XQlw04GV0StyUN4Tvd7WFKejYq+iR0/js8RTzSM6pMiFwe7LyccRixgh/ea5qoSgqn1U7jE12
jmd4ZwgjK+H7kOsA2jDt0TOCz/pf5smNwFA7ieLAXcXNQ25WhIGhYmUPbXO3O121Hi0Rex+4Jgx1
7rIwoqpNwrMehDupBWrgTjo9RC0VEVt1Vdy6VW2LuURfow9DzUHGIpbQN88/3eBqaaezkjMrdFQK
45eulFqVu5W8C0CGnNRnwOTH9RvrWYVb2FCwdYItn1QnKjtOJdYRtEIAfHOHqJu0rqXYyLCwZcJV
gvDkDFErbpStSQgLe9ElbC0f/Uchk8F/YpEMN//xNABl+5kMNUZfQFh1tVcO6cx7+jGw5uKLZLkO
Bp7I9QzebWc/R2ieDOGNAiOwUja/ymUEQhcDzNEvOWcTqm0YnXw2K4nQAgZN60y/JnNp0cD5eroY
adsyHetkARq/eJI1vsIm+Dh4g20Sb0laEvvQ78IjfCoZjmpdAhe6Hxmr67zNqBCkEJ/wdV59yfk1
p1cj7PgXnCbRgcx8QmtLl7GAfq0brbhAGuyTLsJJTWMw3Pp9A0q2XEYANgbhEmSvuArAgiicSCFV
84O9pnYyGf81Gj428ELsLP+uEVqu4aJFFAe7Pz5xsyCDnbnSObVDrrCBhi3aWIxh/wMH/DNVsE8l
qGFqY4BSxneFJaM8Hzbe7W2CLLKjGJrdSKEtNxAY3HeYikfTJeaOcW4O79HLRf7Wyd/WQP1ojxSo
ZIfftyjwhx6zAoIDmM0gl7qqb8ZdfRLP2piE3sAz+oHNnoKb6411iOhhfSvqs54w63IQ8R0xw66p
kprE/3IrakjAJQNSwohF7ehgiUP8OjjneFg+gMO/uRRgvBkNyJiZs1+C+5yCBPMQm2Fs9I5L/ZCA
LNCmqd8ctvgVyuf5TX1k9+Q8gxemjPrymhgE7qTV5LAKz4Rio1xp/61RaIGdaOYkTlhPTaYBYc8e
6DgaHVYeQaan+dyffp43Jc6sV0lcsVj9o8XZxthpDltusJkGqTTVJTODMKCeMSo3kUE2AQ15iw+n
cJxlZNsijNSi84i6v2Uzn30VjaBdvPD9Oop/J7xT4W5sw9qV4G7NuOV2YihxmZ0X59s3obNrs2hz
9TbSaIZcLbSnjyGkkc/OZcJBc5dcEt/nO4ONBPTBehzw5jmv89zLGj04/efHWNqOCObYhow/RgfC
fN3KjqzlQT0568++Og/TMVELSKRXwmJNDgPiLZBBuDe09MU6ibQspgiQSesqKVSwoV01tNJWXWqC
Yp1amyI0mhGLaB5xFalOZtFSC5nUc7PFh9EVBjVRxUrI/+Mx/IGNiijE2lAiRb1/xHU+dvVWbHy2
FfrltOdW1zzF5cC8PCoFWWKwYXmKEAuiqtdXh4X5Xe/IcnSbeYh/GSZSbX2O+tn3WDyC5Ek6szDx
4rWThgwUl6hSrAdPUL1jT6FCEZ85/7C8s6A2vrBelncQ2v5JIFOqRGyyIF/nHS2XkWA4M4UixhnU
QW4/r+eBdkRwNC5Mw3LuLBVKYmqvPT+qqImyF5xPKfv9Ycz/4yapf/3QtV4KnDU9Ft6yyLK8FAkm
1/ydXuY1Y6q2UkxbQuNGEhk35bh+nVCopHp8xmN/KAgFZrpF07UlPwOz4h4vhAX0UMhkWVob0vZ7
airYVmCyHYz0axD5Y5kz+kJUf2JFPQ212nKdm6rM1uuCwWUsLLTEzrkuf0IiRZDwuBD7W7acClYG
HoFzhTdSII7Ky5Z6ily9sFAM3lqSHAVwEbSv/al7maNKwL6muXIzhKsidNRzYROO2Uh7IJN3v0yF
YWifbUqUbRaHQ3PCQfp4zvJbOJCs1VygyijWFXqqCSaPj1ys0/J3vOoQl21LLH/Uqbnq/SwwEB8N
TqzXYVhmigHpPuf33zrIuN6Q99Vr1RARKu/WkMbZPFbGXL8txM4W6u9LNFvDYaIhvSaTm77Cl7oN
jQcdOasyRnBLeXAUCn1qfloET7KoKA4B5wIYCAFtkoqlhqgxEo+BJcai4SUrJjYIoJVP2wmHTGU/
sZ3H7LywPe4dDHK79VUf38DDTyiQTmRCI98kxN0PM6G05UGiL3EMDF6Aw/RSXg7tFmYLg9vcZS/4
K+8T4lYplsD1Ala3vDmkbmjZLdPqOlmSxaqXpY/OyDy3ptKEulPPhDHXCkAYrJ2EhAMNe9h+q69d
jrVRyPy8B6GeWU1gZsPOQYOjwaidDabee2Z8vucSRdSa8F33ZKbv1i7NaQG+Y8SlIa3I4frM61vq
YWTT6Xd5y82JE6PKiaNdFNLDaoSKXpd/7Yo/WaPUyzvh6e8zHZgeArnK81P9+9k2ibVEe/7lK0QI
6rA5hGykG3zQco+dtcIbPw/Xas5o2S+bnZjuWCQ4/Q2POGHnMHApmX+YFogt2T0xogqWsfCStcSh
tzUfH2vMFxdbX/fx8OuTP7uyaoT8D8Ki62Pj1PpCJguw9dV/1WUryG0U15XkObwq3MfvQOcvfoSZ
z304+TJmsO2RP5tx5wpnSKT31U3oKF/fdFGHwRkyebyYRuFSBDMQFydhV4RXg1ikTP/uukb7WNtM
3tpfeowRwm3m8j9CQG8EKcyQiYYDNZ3Te/1rgHHloVCWOtge/+xPLRz8ZF2QqXnPnI6SPf71n3FA
dFKW/2WAaTToQyvBY4m9gTWNr4mP5b83XPUF8g49vLE85SLk46KIXdn/9IsQ5PFs1fQoFK65S1KI
anor1czDq2VLvwi/JG+8ohvuM2OYYaeHnxiR0/66y/Siq957gln7FQQ2n1vNTxN6c1W817NE75hV
KCtRY0ZfKClf0mk6KN7TGCyGng4WWzKg6NAafnjs1VzeiSb6xQCN60zSe8qEsRHldfdYoww6+pcg
pUk5O2nByzMOKvq8ndVhnuxRtfOKPMMfKDFZH8e2lxXxrucLsEnspEwabtaWN7P1yhlTYP5iK+gm
EJIghPDQqwm8NQQ78xxRRl9yCoK6wzIYhLsWSum7ljeiu6qIRBtuFzKMsn/Der/4ANVPhS1Ujy46
BqAKAbXD+IYBX0O2Q9ZV7BjuYXUyJwtoaNXq3M4ikj0ToxUIC2CeESzGI/8V8IorH3m6vtq2oQ1k
6DABVysi3FekZ5H46FOb3WbYQlsY6EEdwZlemHcHAZ9+7R5oil92lDF8gVGjZpVCTUZ3VpyG3BSR
ARlz7TMh1rLcOtNP91Utze1z5wu86teRKhL2RxiQYwiNgv4pn82qWwy54EqyKuhe6tLQg1TCAq4V
dYhktv0NjmFHyBrOW6xcEQ7UnP6jnnKXimj9zDTpvv8qZkwReNy4wHhUIsTapOxuZMB4BKdoPWrZ
Ew/O+opkj+zyh96LvEKbnLXINGWLyhs7n7Gdk6pL67GxgvzdXHBgJZAKuut4E8QILPeDNpc27nyP
JCFZUw1eARIt0pBzdygxvulqSQGAL20xmuN93w9kGTz18jnIMlLDfWVM+McyoHHzplzHZfWo9PcH
IiOZvpJ/We5bNGotMwRHFViqhCRxYe7sfboHZsGDfINEWf5ByX7LwtG80NuAHx1uKww/4XKvRwW6
U2YNigG4LzL5T7NQpxT0HPpMKsDhc/PTjA0Y6Nj6ywdMghurxyoNCD6RHZ56MARZk6FYSafkYVXa
bUNFzFiTcuRid9sx52hdZpORRpgqkUHeQ2oQ3GHW6UvhK91C2M8AqFzskmCWSypQTqpBr4NuwsI0
SIDkPhT+Q2Kw7qr+AMkO5tR+irpGXp5f1rmuBSpph4eAQv0BD8SuI9imlrgVc+8MCbq103uZaQ59
Cr1Ty0aX42SdNsgF8CES4aYwUsWn5Q+VcVoOZSo+oOzITBfaD/ExwXsfrawWlwkhn1LqgKyDYf62
9CmefJQMbQotcox0v00r9o6i0pXCC+CO6Sl9tEYzp/H1X6malYBFoPeTZkhFAPduvq51j3KRGq5j
QO4CMGRSZRJZCCYEhgMBcrSwJkvNKvAusCcD0wlo/TE9y17g2ALiLSBXV4GLEmFdAwj1CyuLI/hD
8QKQOMjAv0OxAM0U8QY9xMB8ruB0o2JB11+08E2zpv65oMcio/UnoKnl0tchPPZJv9qMUzbiLUHt
/yExuzBVTMCuQC4JiPuiRc2hqlhn+Prw2LQqDmyv6ZH63ePyvIgF8IoqTAV8BqHBGwj2a22H8VNr
ZRZTDwVBG64ssVHNDnktY+xW+eWAuSB4E7IcJq3sn5qdQsMeY5AHsVuDzT3/OYlegCxQC72938Ry
2p0vmZDVdFZpwU6gAo1vKX6/8Pnovs/NtRsdqSm80UHA3PYaAm7ZAapi5rnW9r4H9LRvlepN6sM5
NrTuom2uJ8FzrmX4aB0imaFn7ozRTrXPEdy7RIsVjuXLZdsyinytdEU0Cb4T7EDkuv78XYqqAb3m
KN809GZ/9vQo1ACdXW+UgRR0F0yBDyRDjmi/1LFAXj48L6QR3PQNmsC1pofa1wj8BQ1SM2tTO0CW
4D1IBOZImj8y+/r9w5aJpb/LAT/fGZT9ZSygiwITo7KePJhAcKM6TPAt6WgsKizJSvBOs05HnhZe
//6NtYqf+wK2aO+xJEN11U6mNeNi9muryEWLFDSpbgmBo8qGZX0cSVorUM0ccEXN7BXvKFx3UQlO
28r8GPrpYa9Csk7UyVDyMrsAIUQZF9Xncc/mqBeRG9HZnxtwYhtsp0OJmxzUf8KwFWlMmRDQ8WNT
ET9mVRLxYd0SVLfnzcS1izkUEp1IAOKlG6nWhbUdmH6rfK4DnSRKLHT7XjSm09YCrQbtCX3WvKv5
1lZT6i0Vz6pAyiIKD4DyqxshJSb7EhkR6zX4WKQAHCmGmuLKNOsY01IECyRyuZGoXYIrdkueV8Dh
GOyiQwUCsswo2FrBKE3bf+OL4IQa1iOhCvcAVWHvRYe8Dz5p0Az6DTJg729tFeIOIrpHPZKmj985
4QlFJleMsyFU/fdW5YSJpsrh2onp7pD3iH6OF0x0HLjf13Fp9IrzSnJD8CDzYZ30N5Iqz8MYksaU
CgkiDC+91jCRvJwtDgi8jBN44nYoHtRucNhOGmxdqPd5Nhvfi/V9wu8t6ek7IgiG8LC+5KJSz9cH
OiETS5HxE/f7LzA2AV4ddiCq8XjyWa1Mlh/s8gZS4H7czkgijZvCUurFTqj//rAnn9xmGlEQAUxJ
yYuq8PEIhEOXjQoZrihngm9FJbTPMYTjxPWpYekJe3WwcL7qBS0M/uvQyzGOUo0/e2MSFXv1NWUM
QQrWFwtcQv0mNNBpS5IFf9bEGfPNsKs7KORzP76AQVA47n5TGRznxs9UR1464KLyR5RQtt7C/585
oi4lq8WA4ZcBlmaxGV1rAHusSlcvwwlDV3g8qsAI2PI2Xbx/cdJnSCLysENjnm9SRVC6vzyn3hAM
jMEkSCHKhETGJsy8z9FAHO2YYoWdZjakrVznMKdS+ii4uvf8wh/Tfsaca87R4KSCq7wEG6ByXwmS
ZXfWt8WeIgZk3Qx13scwGvx86zPQm9vYlGCax/iwfxMSgKEqpB638vn0Z7IpFaVuiniHuY+pLNZv
Uu+bfFycKVrTF/N8MkVA1Yta670n98BQfIQ1uNdgzkayLh1Ff6+xADgMKyhMRUfk/PxW1KMj+6fw
Ui1ta83RK+VZxDhC4jW5wthgk/TaSf5XRI3vhpVG1Ijn3fHXLj/gRKSZDY2MnBE/wKF9tDZlKk/h
M+omIkLE5GuRs1r8aM70zQLRB+/PNqeIGN/Ogpy1AEyj3HG4/pltou4nG96k0aS4EdMhTo4BJmvo
xRZlfM1AnJleB3aU4xWOf032sbU6dlrTfhqy8HPJGD4vtuEpV0ejfuAzP2BcRUVh5QFJ2lTo2XiC
p+4sv3LL5hoUf+2ioE/fUjpWECZx0IgEuA/5IC80pzoG8WfsclUZiuXjKRmdntQgYCNhUTTnMOSI
pkjsNx0pC1/fFIs6ANf/xC91Ur+FmxYuFnoC2UT3sWoG+GRWA+O6r1ckiOaZuOJjp8sodu7cQgNk
gokmOamBMpmLyn7BYcCuVUZ1Od6aFa72WN5M1ptBt2ThWgLBIRa+Z9+nhc20RFfTELYyaib25VPc
Z+korWCgZN1kKEBPC+h6UwyFIT1AyBdjlJu3Gtz7Z6AQJq34EKIJpUuRsjo++MHkbSqO6VF4dtZE
RqAVyX4YRE6B9pIz4f75ddVgzP9luaodjcO+EYcyg6Gwu1B/DlMEKCZHUIQyqppz2JZGWhrSj6j3
dgoVX6qpk6+a09K+bOeat84T8FcI14iFQUSj4At08fDgtbziQFNQVvYPIWIF+Ogikz5uw9sLa6bL
+bXpn/QtC36HL9aWBbGtrrhtDsXyB/6up5Q5znroky/IljOiAlcffalOqOd0Swl5W5yj72ZA36rw
mWSwa8XdtH7pUpONnmWiC/YWCiElUp17gia+cQD+zqLqXftPiLoUahOGVR6wdu+tBlZ8QmSuYzRV
AnC0h7YHbJGR0AHQmb3Qyzf7QSYZJ9MpcH1vCa9q0p/j9S7mDtRuEYRDPOTKZ9utcXjnMlYjD/vT
OOyInRkpnxGoTxNTmFX9DPGRsVXQyOg47UrwpZuC0obQ3sa2iysDMjlhSqTLYco/hLBDSsMxckZ/
bMXNj7TTmMCxM/lCOx34wUwUlmypaMl/zz5XiozQB92MRX7OMddCHbJNc4Q1DMc+g5rRKf288XHu
hIk0HsYGefEE6IF+zzTZ61EchJo+YbDeYgaix9HIHxBS8KONKeSYw9ZVPl28+bEf1l+BQnr0Bao2
NSp+1l/Jeqhn/DnVg1zo7PvwVY0m3Jx+/jss2uOj/TkJLsr8blF3QbkDTsyWtCz7QHXAe43iFR+m
u96hcLbskP33xB8PIUl8t8bTMHP9OV+PTPRgXFksyFCTWyK9X3YaL/oXjudC/0WQasjMEVuFc8Cz
exqYQL+TIfQI68OPFih8DA3VmPb02B/IY6/c08ZFp2u9ECXeTp10rPbeFdjZ505VHlU8fBXfmQA6
/h3stkAVQSL4rlgVOxAZQcWAP4oY08WmSKnJk4+NTb63hOoHhEGU1Zgjhdfmu+YslGzAAMbQzCOR
Xg1VHERpzZPHjLZrQSbsZDRzH3WH0nehURsXyr++sfr8tpl837o/HqKyPMDi+R8JL458s5ky28YB
Z+d5fWXEVcUnyArEsUK9ofrB36nKehmpcbuKoPvFsoExuyMbOjYA65EuLOQUci7qJR8KS2VKpwqU
GqvmxrdBsjieaHAIyk+ejYI781+QB0AW4kFtqsY18+yQedwzPZLvf9BS6uuc59XgzCRP+bhhVIrp
dbcJVOH4qj2ivFtAK+SIk9zLuDGn84VvZgrLWFNh1iwjIdzBekalatGkgQE/H3DIFe2lS80lcGdR
PIRTvu0DHc0FdIHORCKnQx/8Tqwn3jcn1eajtDkUgy1oF0J99VLliVF3OEDGUK9ADqq8bBBZo9Up
nupbKDD7D5FIRp4HODAqlvGZtdFpkudsWsoKHar71YbauIbtHLc4Ignv++VP1dP3AdzMsK8XpXxR
HZaUdCc50Gi2RVWtDTSioTtGYnd6U464mRLN1Ya+prbdQlD6lEJiW+nuLM11QG+k6dFlEuPUtwiU
6PKGqZGbAONcueaCJ0sMZEyvbPOev5PT21DlR/IoUgh/JBHVMhq3ljsVA870nk4aOe2ndFO2DVWq
mFvyTAvnvJueMKMwo9FjVVLLqdzsUJsD0cyLnR4+MTJJ164iEEuN4YLbmtQcLBpkh1mgL0t99QTt
BguQOFyVxZUJHm4qiubvWZtsmYqmqbdRWH7As89lghhNlQRoQeHqB4EOYPxar3Rx5EsTh9ofB080
KQvP2mnAthEQ+OI/NJyc6Jqm0bTjgVBhQBpOImK7bnsIA2xF7vRKEFFaDXIDEEkOHlef+PbmQz7q
KQ1y2IhFxgPQQhSf6/meIljSaPh05zA3JgD5Sq2f2z+Taj1ttKNQgIXg/GkYaWcq2fKlczIj5Z1j
yYIUAgAzbiJ7q/uqk8BEzJX9qVjpVsGYREbB0aQQLfEm2y5uMshuxK/cxnG5IktUPNRNyUXBUTFx
g4BCFfTRVjcHq7z4weguEqRWsTip8s5Sx8n7monXdNZgecbyUSy5LaoQj7uP4/nyldsH68aySX9L
ymHW1xqnygTkWCI4m46Pj6SPzWfSiEEi413W313QZ9pazX/lREKfMqcQ0Uc9kASORjp5GnRQrFoT
ygBYEJbjSl8ZsM+El4/xAaT6B8u8eJFIDu90G3ovIkEjQ7rFcFuIiP5E7bolZTxHi48lkLjjzRSc
94bIjPuYmUx93FjP5rJvkE+NthRJdtEVVh8+4aALdloqOIYRASr6Ze07lh3CRX07a/E1zSaa1KvT
srr5dxIGfcP/Ugq7Ac+Up2YUroiEAd0Ns7ERtcJ1WcARrOyzpYFDYmAIOXKExj9UXk6zw65jTNYq
8Hz+hhT1Uhz0fc4pALdZyEbalIUKfBVJFYsA74g7tfhxH5hFZDIbxvASxY/bCfzLCvxBsgbpfT2g
/X145UtKyfekxT0LZFepiqQXCNz1BTNZtRu+cT8yxX0JRzIfwyo+z0W452DCqfq5losxyJw87Lro
3hV6I43YtBpYzgbdiN+PhimV7ZnSJbq1DUxbeP+xb+aa9uhG7aJhH+9bDvZCzL4gL7dokFdlr9qb
YM7V3K6DZFh9YoRhSPbUgDpiFqo8rqvTF5B/P3mUabFfCgN+KyslBxr0OLRMj2A+k5eIgSFr4Diy
NCUn1yq4sdOjmm4sT9QZbczUoNCJ+JpfjeWU2vnqxfhiLpUnXtiU7XXXXC0DMxlblOHpJmDdgsju
qj/8T2yFD6aNallvY4K6KNGc2l57SG0cJOiEok94MB1cpU2mtaIWYrh0TVlF2X4A/RS2SR2MtvU9
hOmXgyavtZvrAydZAcO3AVEl0SvxOjNCkukniHJ6cPyXqjwvi2jzXjtRrCyIn45SgO3nd5kftPrp
7U9bAMYF+KGE6PsNVnfMxyihCHcHrwVx2zh6mBOcipBnFQkGy3JJOQDNHJCEAANzdkDja2jFP3AV
RejB3dR8ycZz5AKUoNW1o9wEMsCseK7x0lPRu2OZvFxWZ2R7IM1QwsbWOCoX6me4MVnqYRIMpSVl
4L+O6c3YLRvLczGEof0V0ujR5KYXsDC9ebBqOHgej9bxTZcHTTusFrGff4hH7Ilex8VhEk4rt8Sw
iB24qVOONjkdvOYsB2QCgZMlYQ7LBACfwpAImaVxUotFkHyrp48BxqDwH9OG5TxwKNoMkvU7w7bm
3P1u/dIHqzKo9FBlv0gZtSnrC6gmi5xLyb7ABhYuzH8VxD7wiA9Sr/hWNBCVtlne1fIx4reSqRS/
GDGdqUBLvr84C2n6abRCCnOLH/PAY+U9hx0gJadirlxQCr+Qgjf4ms1STCm/14fNp1WOz0Qcv3dB
CAxcwHzkn/HwjGloaUI+9/sKEmw+pg3B3e5G+XBWzVx7bsCBXa9p7aM/GsAGq7oCgZ03vlVfuUin
JCKPOXzYnbuPHHmBlY9qGV096czaEfC40F3rDhai+hkduUZOQYqajbwaANVp1hTMCU0vbY1uqd/a
nfQBMT0LgDE+oVdjjDDUIffDgUaQ72dynlZMDKXNIPgLSG+xdqKHIryybFuiGI5l/VGyeHXVdcf2
kOEvNEcYLxu5qm6FXF25Van7GKF8MIN2MMi1N8COnoMKMQmsCCRx4JiuH1S3wYan9g+V2J7b94qR
1muvCVjhulffv/w+AFhRfCs68goOA2gebj0jQ3m+3ZcF1CGUkoE0SgQzxdkcJylb+MR+BcA2W7Wz
jTRtGFVwkSjZLkql5sjET/DvGHC0IEKhX2o13TFW8wwJQjMkO+EAGMB6K/z1zKWU3qiWGAtFOoGl
axaLiIs1Y0TrQZDkQmuIsLgIjty6kmZDiM9Ng3T7CHQpTOhvlZ3at3B+ghgNTQYFxTCxXanKeXvT
lgZci9z5GkZD19Pagr4hRJjJTvNwFVBhaTW5HTWPqeBsgbEL/59aBFc2gy9ld4xg4BQL9u+7giyR
bE1GhuadShPlSiD2iZt6/PSV9QsbCb8KxIRDkxoVWQ+pzSOpNj8V4IACF+Oz6JvCnLo1RtoBwype
zUqPK530sRUIV8uxryyYTLm6kDN39NNt7MZS8ODx+j+u5dYUiYfvYjOJAM5OYMT1WNmzMn+SHsxN
OcgR8yJSQ0IrG0XY8gUf1MYUXZD+jAjIgL6bvy1ikoXOM+lZdw8CPIWJhJ8nF+NpTOdJKH73AA3G
KJ4McgkkQhLy7/yH6bQzf35DI+kYoajZ/bqt8OsmAulUtaFW4EVapT0a839LLjXATrSFjcy7K7az
7LcoM6/mRgC42Dc2rJi8RQ+HH6+OuASZ4JJLWrub0vcxWm4DW3lyhuQ/Fa6lPH5jZU4HUzwPLJ1f
UwJ8wjtvxqm8BpX4Oyii5HUWRYQ+av6+A/FS4oLoeqjcKbldAXSwvr7Qw50EJLQ7i+N071ltxkEy
pTXFTFq4SVtvyDYbibUQDo2aRQqGYMeflc4M2oIW1Y5Yno4S/HV/gx/L7NOECUDwgONIOJHtJLdw
/vdySQk4PwQLXxm7W9qgizWuXMQaktW8q7WzT+EF2XlbNUA4cheacAKnj7wzlMS4PhXYByniCqd2
15XyjTPV9EkgoC8Q5CUPfjRZWIXQKSOZSShgD5N89NgjL6g35TuPCSKYcGUKWsg21ufKMwXLVnpy
JQ6380LwjtKJ4pTovCk37tHR1/4yQFhBQ0fdQSoJt2ZGT8H6joem2wWxSEfCNwO0ZXZoxXTEf1vJ
3EqtHDPtb9OPRfeZvk2PXoXIsH3EnYmUaI2jLCx+RNDBUKtcF/t3sN3dLk9ohml8059j3UMngV3C
gaBEIz71OjEQkIAPAcWEs8RHTQl2hRP7MUat879YO6tXQwxVZWmm8nlLSnFVIHTfDOltqpYqmOyN
JY8uPqUf2KKy+6tWcOnk4HPy7I5jOggvZZoBK9UNXuAJCCADdOmewc1VS0VrLRRuItvdGWpuH9/J
X4g5tWxoRG4GOlls+dpfTciCmUlLyLo9G3jR0BzKmj02u5GUEb2qMjeFzyuBhNOhPZ+NZuGktDHb
URvDdMU7+XLybBYkRtjrCj/WLMK5GqB6CCgDSqAMGi2/lVgZDyPpGlW0Tl4nFM7X2Jhmm04LyQ7S
Tl42hF1UEHHbcZG2NioojJQ74TNNUC5MJmajXJpVEJc76J7LbdAP7T4i8/6oIRdN84DByFKKoW4F
gUdkXmYAbP/pc0AUn9/ecmLtFmyYfvol+pO8LPdL9bouoti+9woYrk6gpvj/aNCnxKLAKRrttFTP
rVYtE2Y4d8mGHrVwrFOEX93MiA01lh5c+c+JqGrDAtLIkSy7OxvwLH9EryTaeQKQ97gIwD5O8YC3
Xm7G+7zCDLFbRnOICVERvR3XghLSVp8su9pmxbXUuP3mK4tgJKDVmX4Jzs1SCkML8sHQ0Yp6rEWG
sb3b30VxU3bgK7iXAc+usrIU0SjerYomIEyicCfNZpLtfyadTCfQuX1GBJktmpeUH8F7VUItkDOj
ATIPeEs+htVTaNA2ZOUNu/iWRplTDQDI/0eDiN64/YCKUXy/6ahviS0lAklSjajKZ3Id6EvYBUxS
ksW3JmETWwBw2c9ftIgALlEpMAebIBmaDuMZee6wBncpNA+ftCxTdQblifnYeMViIh35Lq23IG91
mvd/Rw5LMOLvdKkOG1nB0AFt+NjQjQcUc823L0DmBHu2vGMIJMd5xtHNH4qxzdlQRUzPJRVnjCum
+qgcQ0rqC+DdmF4Ad2TWA8xeBORLxGWdXyX8YvUsqdWIY4hgyohgU3HPQHgywCf3zrAmXcMiD7GJ
WIAhJ07FBTlufWGcqkoLNYQL5VKc8e/qkAQTW730Ue7ZfV4WHBQONg4DssVNypt2BM/T4mpHlHnX
B75focpu9AwHc+EE/JNCQtY5HiGITwWCH+0RscxYJphoQ1NRNXBrHya0xQMBNCkLo/xJ2Jkts21O
m+btutHSCP6Wza1cz3srr7YXhDc3qe1xCLMpz1unL3W3tXT2ajDFHBYsGmF+LVCCy9zcRvJFluT6
dPYMjzKLJqxnb75L5YEb09AZvW3GPUQY6H9V86JC40xQpD6K0Lhv+FJ7dQ52fthe0ifPLwEQ7pPh
b0xz2ebJb7g9ODVDgdtgwFWJIAYH6mwmDBmM9Sql5ddYgzef95UxwT08pahgTe9pTmpOvfg0Wur8
fFrftBE1//YjS11KOENFtNJv6SrjxYRa4vJ6zNCxfJis5stKcT+iyNAwspxH3Rfcs7cNCNPafVjM
SsqiH5zG8M8pEIXpxi8appyd5D5jTvUlzkELi/tm0MrMSvW/dd+x6DmL3I6hPTrfzd+O6geZSOQY
PwBly3e8yIISrzFS70ci45lCgfj977TmRUL6/2eD8lc2kEi03+nytdLNPrbbwvoxv2ZtTZsigUt5
+H3hFTk8adcjVVJKNcxL8ID4KllI7QLqk3VxoUiqtxzd/qrKVFnASPnq2aIVXwuK2yodBiL+xYok
S8ViYG8ATHKlOf3u5G3gWp7HuH5b7AlelccJ6ggqZl7IiG4/o8Ew2GbasX9sqZe4WSRMKur/SkIb
N3+Z9ax9+mi/Wff+huO4SwLPWTohKyYHlqoaAxHTiVz9wcoj2ncRWShmH4A9wdiV0t5Vx0JgyeE9
e8wQ0sTaIDl+5lD6zdOqM5Zv8i784T/ESwdCvZ3iHCdxPXVkY5oZ73QFnS74luYh8NldHbnTpQcr
BGHlwTeWGOl/7Oh21k8L5NJsfc6FY4+OWN5LDKCeJ9Uj++XbPxynZyohmuvARKV5rWjAas93Eo91
0zVobBe5qOLxR7yacXDfyhcCIs6elRFOqGMlYAOY8SzyAsMV43Fvr/SnK/ydF9hu4nnzroqx3z8c
71zMVCPpifIfj0ZgL/nIF0231HPRf2/EACq3Dker8kHL4nCrH3YmBdvPKeZ8C9Gwrq+pW2ztYekk
4maib3PiHssvmAdKAHvUz+wHMOcZE8cSGy4wyt1NtEdIv3Ax/z6y4S8jWAQ+JhWMNTv2HazoTi2t
xBFX2BSTevWgOTYR+xVeKpm+orXoLj6n9v3rHPfBnvWtLTWdByVl+cLVK+8o2OJMt1T74ScA/GWF
MpEHdZ+UcdP+eLmWeRQL438tSqdWDUIlRab1MkIZz2SqvDewcmnc7K0BKM42CwGCJzcySt78fy7U
K+OqJB0MCzo8sNJNuA+WLFl8Lsf3I1rhQQF8mWxPkx2wJ02Mjvf4o+SPdYJKXwENZIKSa7R9EiNr
4SdTA6yjt5XkP+XBK1j3wRS+QEpAJLGfpGtjgPXXrh++xdE7A4+l2idNqp4dpmGeccyQIjGXE/zw
bk9VwgUXVMHCNPrq5q73jjoEdq9daRern7ZBbwWxQ0563OqIUNuwxGLOKGIWmlzpuHLOIKACLaIO
JLqEQP89xe0W3B3zXk9sCqkumbx3/fCWXkJwuSWoqLco8I7R85mkC6L/3koI9QYIDxwD6zmsFiPi
8Z412eymGX2MfHfNACtglJPMA08jOJdQFvV5QW6QRP1PPTghDssRtD3o5QFxiFemhOjwxj4BT0er
2MWF1t/10fWmvKK/VqiDCZC5vboqrqTciQBJ3tMPqg20aneyZ/xGXW/Xm8s1hvTVKbxaPedi453c
YUG9oxi4ufRCMlLA2BS8JzbiqT9LOOkMwtxxfTcK6YE7yh1IYJzBJZCbqXCt4OpAVfhGC54+gdzc
HXNTzrem/6lLxKqpeSTMeHJIIFwVhGtIfBFMdQJPcMkUgNMn+cTTFhNaIWzzqgSURrlE7mjYhBDF
JCqoPgaR+CMYvX0/dvs0BgKg7aBps1A12yx1VdP1pbFrxZoONJX/3oL4XWgoRKFV9ntbgsigfOHS
heV8Ennqdrzgp7TO+nvOM9mH1KHSXNRVoVGiAVIxLDx6H69ItvIwLhaG23bC33KaJ73k2Gm7El9i
HGRpOgCJuHD6T6YgFVXA4W+V5WBuOWcTzIuh15zl/VvLJFTUUxGKH6t6pFC7mBE/bDMOio+BsI29
PsFD8COI8Jm4+1IUNglQNrT4zy3MrVJSESgw+IYe7oLuUbB3e+H0ic3bllj3xt1DZ8fMEsH/9VEc
1hMbXhkgWxgnVHArg0biY+ZwvmgsMP6fFHU+vWJsFLbmzmJi4R+2YJ3H3IsBtSjmb8nKpg9RQTDY
+sA0TjGAajQVD00StjXPgO0nsfcMGx5t8767gp5Ny4Yi7ar0zKthXjs2di4vfRm/UzTkAmPVIdC+
3kNAauKL68qiIfrGEwdVoPQpIS9aB5b9h7r0U13pWzJaem6KNAp0Ot4jN6jhiyLGf0QfWRYU0O/C
B4iFE+z0Q5Ijz7U2wtoZBZE67ZKo51GfPLLaQv94nBDvya7c6T6gcsrHiRxKSeu9A57jd9ZAAwNz
jF/PNXCamOKRohbSUbgxiOIOQyNLnzRyJToeXL0sfKM3MpE9kgMCuF4dQL5xQrUfkKHl2XLd+5qZ
eGsV1nJ1tqcZ3iXHSum1WCiXSpy3QqnDGuOw0jgYerInwGawLrhcv4zl8kV5Haplt3upm/pLmLQb
lsKAEdbaExmHwnARPCDAN25LS4TWcix+VaRfw+bJ8wJQhqC2NbpsEzsooD5TM1W8Szj5BpJZ1kXI
XoMmbs3kU6X6NADnmvOH8wahpoUwPfqlQIo2jC50GCRo/2LzqzGjvjEzaEH8HOwRLiMxkHO5KpOX
u15foISgmf0i4q7N7zDeJboF9kLRzqUSQCAop4gUrROx4K4wwtaC6QFzuA42ENNnFr+FQ2j7jCsU
fsLwNTDMozwlVLBj4wA/Hc7ucY5VQdKS3qZg3YCNOtzwIjpizPRnCxdCMuPZ7QRd3knp2sepootR
ecijgOLETAhIZsk9cvoUTrPs7i6N45vsKP+Zs/GIMn6xR4UURSU6VZQvE1qCQKZVWPV59BMeW70L
Ic5vrtesC8UgCO/SjnFmWlCYvZI6Snhq7/Df87469ZhL2q25GE8sVIs9M40FqxvLHULx5LDzh2PG
fugqXcR5sdRZAr7FSZZ6fm5VhqI0ecXZ2dLCT7r1pLFBN68e5NIN7y4e6bj0jIWAmC4XydkSmR0X
XP5woWKIknWboBKJ/g87O4c2p/2sapTXKW8wW1CoPx8g6SNQXfIDhEhrLmoN26o8OkLS8jegcSyr
2uEJXE1d/czsCdIu4+z8C24RqNQN6Eod47LmkPSDBlq6TvvlNVVaugzyaGf5gvyKfGJoIs19+IKN
7ajZiejrHTAEDHudvELoU+4O7HBt7nrztK2ZUmG3yFpY8qjWw3/b0+B3Rv1VQoHwA68m0gF5kRk3
ORYARToR2c2JSrH7CUAHhWH35z3e6UTqkAaUtcvGdu3VoYkZn21CAfSv8rQ3orEkdSDU4m+FwLiC
wWhYb0Zo9SKl0MvTFnz04PhdfU6GJerV65TI5BQsJY4QiyOfmBDiNIDFEfdMSFv+/hQyjt9UmaQY
mPoeNyapf471tnoUYl9zCep66emqnMM8wsSsCfC0LqD3M6dZvRpptbuhqLS8FiLCXgpC5FyprxPq
dzLk54u+Z5tBfyJPA94pUg31Nhe6XPtnNWx2qn5SOErFrulQ5cloErgfsOHl4cV3OlpGghSDXosZ
aMUmOQSK1cd24HO34XDcF4r/Avfxl+EJQxsHZa03E+4w184XZ9uw8SaKvgd54kqEc5xR+r4ith/Y
e/1kBj8qir8i8z1+BSzG4KLJyQQxckQUL9F72asSFEy3j8YXo4xq/Wry+yuQJMPzRt1IcWvUqdkH
STQCZEaZffQArNzx98RlDTRtNYg4VAHM5WUDRDnYVoaq3uWPY27rER/utplic6Hj9Pa5BOolTjVo
DepU3DqN7Nb5gdn5tLt5RyGczofLToKIka+GHoq7MgrBQ6GnjkI7dZRRL+tgsFDpXjLgZHKFkTtZ
3dYWkOP1EQyuAmHy2P70azbkTw08DMLC43ckIwVrYklTbPj/audthKgr0515mYLESHS6oS0pjtld
myrooN1UKF50YGXgiLJbfMcvVcgPSlgUh0u+X3Nna4Myp+TJPM1o+o02jvkE6+6UixMpvXqV+tWW
Ds9kMY8pfSQN278d0FbzggBonNFEMTPL1dyZjY8IKxqLW+C6KjwOaoN6qocYsdOhhmRSix+1ZLHq
c/5X/xLncErHy8QF3hTw3tYe+MB8pw6Zkr8TU7mst1Iw/oYq6oNijhlz0rIYYYDYgjUo0/Og+5z0
6oWwoqcVCvAVCrOpIqosZPNRCO4sf8Z+r2C1WzLV5BsZJPwWqAwb4IOkOlyPv9aOWla4VNIy3Rh+
5O/L80XVp7+k8yMt6CMJwCnuP2dZPkX1lqIo3Ray8rtEjvjq3cNkW4xrXmEhyj+2TGCdXgm1pEcE
t0aEIwCQkL0LIWwvI65yKJtVBpde0/L052OAhSPPx4O0s4/HsYHV/CJi+xhpRns6QR+5kU8R6zlW
cMoYRir0g8JPHpt9Iy8LKR8i5Kho+OOlUsoRZ34u4a3RMg5NySsdF6XszJ47Edh9nRb6e43LbiLu
08Vse/zrD7Rj4gtYVaRvzRvIpSxmUYrPy55PvEPQUjeMAH+I5Ui6xZL8kR0mHGzjNFTUllcQjjSO
wylvQjvU4tWLeto5lbJXEPuLfRe3ao1QYw757lRSxLLstwOpdx9uM/E/69UHXe/kbjLCsMIBRwKz
xcqNN2McsrhQp5UKfHUn5tfTUNQWlwGzmEcvwxmXxdwQJf65+uFE3WfWuthEDBEUSudGG0gGI+a0
kChXKLx5x9xR7eAkM21su+8OtduktDCAfR+yI4OnNmcPtI69fTNuq9cSueokSt3SHfI2o5qnlK+h
79wx1e/JK+tXdclQaJS0wCy6Ies/UVVilnJByavIbsJEb1NK7j30B9tMnTbi3BJi+azDGRms64aF
u0xPEMyzxyR47UmgmsmApMxVL2K9Ux5VifJho2ZT1N/z8HybDEuo5C0GPSeg9R3Gh5nMFwsSfwKB
ch1SFRSPA1lHaWUEneQg/9y4+Pc19TU2ff59/AlbQmVoWGJtVuGUSNx4sq7PE/oH5sQ92mZrIsv/
CuMSsBsxRpcH5cXkhhdcYRbmtLMJhK7ybB8AqbSnUXFxsy0PFfJcfLukeUbA53y6vn0m7e7s2ylx
QUzb57qRu2RcIopfKG6EEhyDtmwDmcPWMxOGCrUkR6RBOa83+fZdgKoXCduoZRdRvGu3yHZ78Gq6
KoZFg0pb8xfiaDUAzUhRIn/hFbF80gK3iDv0RFwisrkV9oBFfsWOSbsoENnAZ4UjYM+c7oxx2ZRF
1HrHhOK5K18bud+35rdmPuc34ZXMXUUny6q+y5yhnsJpaavRsI4Fau28snHsOD95BbDK57SH8Ovd
PpwDpxXYkZI8xG+GhMW/eJVeFkvE3fQSk1tybWk9stNsvEd8BBAQTG3fBkAyEwsgdOTdmRZPK9QS
9ghKUYPl+Q973wjyzz4gbMHdYPvEu7rLUZMaovijdybrSP+2MRBfDA58HyjnEFgOys8sVpXEzdrN
dAGrQ4T9sSPkfbgCX4UOMOX0P/u4C7DQUte3TmEexSzJpxV9Q5kdRni8HMFbrf0gdm2Krk3xyVWu
NkceSYvUku1LFbwR4rIFWFtdHP57kdhHJh7GcxGxPcca4esv4L+qLMHdZgRMVi603xXL72jaUmIH
IuBGeyUmEw0y80ITg0ITCk3oGAbohOB49NKR6Kkw/1jp7NHbs5V9Ht6YnF6sSCSpnuwx1gydxQFv
CKjp77oCPumgSM7OHkgZK5OqLzjP7n/TffEgUT+6NxUhvGCD7vN9y76pGFVgG5KHeIv4KCwtKihn
A9Ye1Le5i8POkInVTP9OM57Lnh0UEckCAif/4dKayym3lDwdPvFvQFObhAO1zujQ8t/C5RAbkyRW
sRuB9Lp8NHoVvZwGE7FbhF04t18/aSA1vNG9zS7p+AHhoS3C1S94TtCr1Ng7HMDLjJH9/ImKfD6z
o/3AzNXIb16rqSluzkOpd4N02QVImb6lYgp0mD0axU4eCuaCFvZrVgGL5ZYcXgdvuPgJeCG2eE8z
3r1j4EhpW1IU4fhQaMh759c++/NPAY5tuNhBshg0/a03gQauwIiOe+Yb/tGL/Ki5aFof5NpOB4qq
OtsXMXnfqoMWyy28GLs0JySzfvSNRroG/Bugf7So9uzpPNppQZTQ9nnOMN5COPEuogSju+Ijju40
jhFE5kQzq0tjO7owHXdQ4E4QRC9P6NWoY8mMB1Xu2tTK5inyFO7Bb2HPMjd1uzw5t6BT64Bsixn0
dKB8hW7uAaxV/eA7+bsIewmRuGw4nxQ9R+VYvHloPuLO3JMsoNQnoXLuPrr2yuW4DJC7zSUroI/P
ebKiMuUTCal+qxK6HokUYDPtSNsTN4elNFapQrzm90bpLMEDw5T/TxMIikTuhkM41W6eeYQpoNKU
62cSVidtKaK4JbLIbXZ9/Y1fpmdUmNB1GZFFZLD5pbuLgxbAgs5YzU8NE91Vo0jky6j7fo0DwCeU
bDfsD6Frs7jFYN9GX/oEEENp9QJRQaIta63Gosrt4rGyEqMR1jgGBX/ChOizovguZFpNEMMPjEY+
YZ6nk0AS32z2+s+/qxx/7WWQLZgTBgqrlVTQx+LhAa/6g/PAbKOVfClPdHAAQR4YZ/30qV0uHVyh
82ko/0rtT3L77xPL8hQvB7U7ntjOBW7y9VHPvsisGMSBI+RsXnMx0dcTpgHuIzgjcH6e2qjTVbmD
egtt8D53Uw4PPqQ9oK6bYDGnIJi/5iDZqjX4HE8md6RztLYiBu0gSjzFO/+wJkMViHWtX4st27FV
Jo5K+MeqLmfhYoPDr0NFAsEb7gVC9Tq0EtiiaybAfpEVMRIne1qyVpaBSPIOpB/k3vlW15pyVP2Z
SsGubQZuNtHmU64V+itxzPn3HsG1H8BdyC/4wv2cV4YKxN6m8hyIGW6BZPsyEDoSeqlgXXUNtGpz
PSIlaov2Vgf4c22Tl1d4DdTl6H3XTqLZ4nwXAtjMR1oFWFwlskg2u5d+Ji3yPB6bUrb44tjFwp3a
8kWUUgnn6LmE20Uxg87OunZPR2/7dRiRXVQEMxiWCmMF84Rcj9bDSvz86Ck4RknoqqIUO+jRax9U
3BmjAx0He59/+87fxX1k+HM4J2wkpwuZHVxTA9gvx8ZZ0lt3wd4aPVoW1bQB3FOgY7OpJ3d7o9Pg
ebOCvfrxs/3T782N5c1fheUF1DisKwfauqxyZyIFXFPo+osTbY5Ct7KS02F/UCTB6kNqZoo8yxQK
+SuCUX1rU0jyONCSv6NCd/N4CDxCOKSc4wCobLGEfXnCIvbhfOF3sdd2F85jfGnkWtkNfTbGfFuY
xbzxXjQrtTagAr3G/XhJ0cW7ysZ15nhunJCS3hioPABUkbsxkSOGmZII0tybkfMDGRJYHu9k46Ji
GnowiBhMSd7bmHhrNdylakR7eEbjqrAX5zE6TdGDzylESJuapI1HUYzixdp8sEeRzoQ3ofaw4djP
sek99DWXLjguTEeCw89/J6GUv5FzboWS86Qfv2p0/oSzx1eg6tl4yG3GwCUjwhg9P+9+YfcHnC3a
qBdti1mN7w9jwUFk6QZQ6Kbn8DGbUd4muYboUvb7pPJaVsFskY0yYqDaWOVyiN+qfbCteMdl2rUA
yF71B/8EGBMxJ36GUc/ZlFGBOQreVSt+bBcxqb+2eqk8t31ccsTVbP+rTKJ6gI5uZtSsELGxwmZi
bdwDi+96OvLarQXzPCvpMSfoE/5Q0W0tVxzNEftPdC9hKF7GsEQ0PiRUtjF4ph/anZ76j1LPIy9C
pfh27m8YEXQrvvxWqpMvjA+9aHw7wDDIkI0n6giLNgZ532aaVy80AXL7bhVu7OX+9+RCbg7d+kzx
fCPU7VTsY804Bie5K1eLzPEc0EVpFKQzW6As77u1H5339dvyM3Wj+Pqah0vjGaHCFVqwuYPaoHZG
yeBlwlMolCMJYDCL8jLwfF7WsUbDp37XH1LdB/g8jrJM7x6BDt9jdnh8nZ6hCae3dshsopWgsdrW
uCTPf2quCzKniIxaQfHoVeFsx4w6jDhSTRd2Od747T0yOy27nP3W6XWwNpR+REIYsmyjpffS4Alg
iy+YDeEJHBmtBHAH/Ynw9QPfq8rI4i8TFgogBZnA8EuMbLXxwe/azetjT/TcirtJjU5LmCm/PWtF
FKt/cvG7nmc1XblxNCLrv2ifWy+5myLyK8/fWRkr4ETXstvvCLCJhwnCkh2t1a2GbspSwSKKD1fK
VE3ZX/8bdwyQv81vMKyKxNgAuyum3TKPMCnjSiTu+k49HUm+MD6Y4O/MNFgBA+Sx8k5upxnAJNHm
2QaNdut4Ea63kbIeQ6WWNXHkGP47NNINRrD2B7nGF/WvclKIz45muLmo/G4ckO1USnnkI3WOsL3U
PJWDWWH/09rJ8IlZYKK6Uul4rDVW0Un5OyRCXcZQcpFCIV5QfPZE1b4uyyaVUqk3VUggUzXHUbn8
Hs52Esp8QnjQ/OrfPRekYgfhwzv585vK6tVN8i0TssfrdhqIkt+QRFjyRy8A9gUug4rPLcKGtjjO
LzNgStWwLGPebCbNMa3efJ+CC9HvSh0aFVicaJCGeZzx9+lRypqieJ3PNMmvLKLfv9j6bunYJwyz
DvG4shkmsGMChIYQ2KmwwBLEyI3eU92GYfRL9CfN5XHtpd/SBtkuY/obqjwRqgSjOy9g8zw/CnH7
1KWyGdz+EU3IY/iSUYV8gjEj3SJH8VkM9gGg9gHXF90nOLTOjXu12czlMu8zyfByt90d+3R1f2bw
ClxRBQ8zCVbVuhemW/pdkch63tAgmfUG5c6vRNEyyzTGKePWN+cZb52kdkJ+9NNcdLmQl8TKQWyp
ucRx6HK+z62m6rxdRs6IXSm8NmhLrJUnM7dMUreJLP1/mwtijQnMJNFIRjCyVCSXRke0ZRIHTucM
6We24yNoNqotsJAynJ4XRWK+OLusBo8b3xR6tqR6filTgb3XJ7gjwdOQZHgSfDPZWPHELbRRy3g8
jkOgBYvqDfb0VpFiDQoYiKECnU2DqV8/hPwjWqwcybE0lSbnM5gJ4ucKf21NfNhBvZYHlFMp+v8C
MkBT+pYYs9LgSRvoYB4ykmhEQ35YagIPnmYGAjZz1Kne1YaXtXv1OBEvnbAcadnQxqtqv7Ee73E5
jcu+EZkvVRmmmctWRoq/naKIN2BjIH2u6JqsRyFlvMqA2lTB7dUGNUewwZWzvFzm6CoLxxOpbFfG
g50mIO5V0syCEvD710gqor7jPjze/rpmOPI72bKXQn/ZdJFnSd0TNaOU3XHzR8BWxwYCEdqEExb4
qZBtvNZzNl5+DmQ6ii00ibRI07M2MjMwcLTVTH8FQw6wNoB7wWTnuMGUJ1H5N8QZHEblHiKcHvT8
HZ7fJ5Xnb8HJBAJl2qX6aSNDNz3V2yvCrbUU1oFtIItivCM1b6s3kITiqI53L0svKWYKabzQjWlj
swI6LNczTZiAoVt9JxlSYvZ1f6Knf05IOFXIRWV+LAY3ugn/0rd6sxpIRgjwxSO5I8GiSUkJjKJ3
mieQZ849mR1YDLnrOX2fo5Zv4QTisTjhETzcKCcLHcwCFjVL3BQfMrdS/rgxSr0Yi2E3bifWUHc+
UPVU1M1AIJaZqDSKTy7Tcfz8QZvVz1ol6MX1/7tpSQ4P2dvOgNog1l8ciGexR4S7LsY2iBSl8it2
T0zQwwOTz5UgkyB3WIY5MDtKrSobxGnx8gsmMy8qV4piKn08bFzFl36qyCbNGgQ7sD6v3m1oBzVD
61+yDRan1PDqHpqXARPj3FhEWdySlpwIzb6v7IO8qT9xcJM0Umfqteq1sMM94j9c8Eb5n0b7AGPl
vJBVb7E4hwVVvgqgab9SxbjoLmdbA0SsqWalmtESaIUytxisn6BsLSDnKqRbIkFkD5GkoNuTRvGy
rK3zWAMghxVS7uC4zViYBDSVXXUvx8n2ts7ToUecOql4WrHm/5pO4oNqwkE+F2/LZaRvr8iLWbks
YBZ8p56GGnWk244pN30KUeiNk0+Mbl2GYpL+RzgIfs5iupL5mCVK6Uj1HNzhGhgwkoHUDBQRu3ks
YodlxCwI3e/QUirO1vcL6Ku17D7JKreitutxal0n3YFlveG+4E4ywsDw+YVbtUpUuNgGRAPukPAe
+8FEJn+lOJCj/fXu4Injb5jH87Skf/fst2XE6qqFQQYKFumET1sHXOBCyFkuhiV1HyCx7in6naNl
//b4/uiKzu7kt5U8rJdCvbpWm5KLdsVU8kGSH8sxHo+5XksH/O47PSxOFn/LMbYB1D3DsJgtvcTv
EV2lrD4wSB42P/4QgXi+u6ssS5L4/j3c9aBWVY8o5CTua0ZN1Lm/dr9W6kaNMM9BNT9dfzKBixdI
bZQ2r5inoW1DmkplQXS726IN2J5t4OdvnM1I2/kC+WniQSflevcJYCsyO7fCkcPolICPMhOh3snd
lSI5s0gCUW4GB7kln47+IFJgSrXuxeQYO65F0+GekCpGKeNcwrS9qib5cVRecu1SV/6pmIZ3aWnv
icmQj1Sy3Y1veArUsD0MIzaq2ZqepuBIUVo9yXYcfiy8BHd8PINM92s17UvzjMNEVLLJfBkw3gXK
sAQVITAbapVVBreZ0IlnZKUR6COU4t/Ct3UOfhgoHPmGvx49BXYAZu8DljD5gWU5caw9vfgpobq1
esiGD29Km1P+JecJuh5rzkCqnX59QXA0eBXrTOM54EB/1nTzQo/36NvzMA5R3H06K5AVqREyDz5Y
KcE7w5ESkd3UhJvmelL2Ps7bmRLowo8FEIF4kZh0MxSw+jjxmEAhDq736htQH65Sv+r9sq5tq0HR
868odan++WTtJdlkbz7UCreYviiZXEqalFiEwZFOjZ3kXQLlbYGDbGyF6eV2BM43ZL+nM4THBGI3
vkxSBKlw3tGW6tXz7Q75axBw751WXVsMieZdjTWD2ghN2NtB+8ImiJ+eZhc8sbctHR2alj3jVpwS
2aohreCsspPZNsgVRfdqmxisCVC5DERh8Z9Sbf4KeRoSN0SkWglCH8hBXnBj9aRbBFCCMQvUwPKb
5t0XkAovc4kzN5+A7bcD4dbCJQw3JZnd8vVtcraKla+9tenCKO58k1fKSJEFyY3yP/XFTjtw7ajM
2w9gBZZ4Q9OhYhisjlNg1APFU46t1HAnZBzB/nJyXt2kvDXVRp2uZR84ESVS0Lq5ImcmFX8AG0LD
HT+d9214FOXGFpVPGq8S9pdZ5BJxBpN5P+HiGVKYNrMN7MS4r/7GhNlzabOIWibkDs96DfZC6WNY
u2HPMRDgVNStlJH+7tLWyVG5tZjxYCtsJfeo1dq/PrEILReaMr/sPhXGLdu+eOEwUO/EUSG/fqYr
IlXPmHW+qPHKloa7TkPFyiQ3bJPGAtzdPmqypWpcH0FAa06FOtz30YRBH1Uw9zbhlBbz8meypETe
zamaaG1WBsVIJUHv5+RDb8JDShPTayFUCRW7ZOtPe8CiqGML48vND6kIHGpUM1YfSb2ojoEL+dpv
divwCM2hvhK5ax5MAOTvirWQkcB+PLdmTqjx82PCqsSHdPOdQjCVzvP3fBXHbG2ES2feKJJ3ihaq
CHR6OMuqvalDIlBoy+Phr0whogOlKH/5XLQjMHiOxN2h/1Jqtpel6y4ncmQMhvyKiQhtp00XD7Sx
JQZrKta3iv0NYkOWIELs0DLPpOg66RBsIXUzZZLU0IAyYQOHTBN7CLrQqdGiCOc2dHywOaVFxFy9
CIduCgtqnJ+j5tZZ+ssJ5p21jsOP6C4zqICknS6qWwyvGyb3QevyHf1s/o9M10a84oohjb748zPb
JfJ9V7EmNmfN+raZbDqjGgUFfafGImZQa2rlKUHKqmeHYexi15fZEW6OOvMEtgWyenQE3qSFngTm
udUtQXIV55YG71NYzI7NFL2SlyEbIROb4TyaMjTHRo9PHSxoELHWAZrvQlVqTRf7KwZecKHNFhjd
yHfJmXlootVTNPlf+/NK+z5GPh453STZK3tbuLWkHi1oZ83b09/yBcFY4UonnnbSvUXw/C2RunhB
lKWC0OXv00z+D3XW7O9V0ts8tZyjQCC/gHmP1fs/LaGdPOaJAioUqthy72F8cWnRlK4Q7zfdobP2
uc6k7HH8aGwakLaJnv0GnP+A0q7Ow4KkGttZao2rDmQFEDPll1cEzobFLWZzI57iDmSoKvQg6tij
8uuPsTqu4wZSF2rEa1fWC52vJjTy4UPzj0uQZFfiyJOptyFAPRWt4sU91MYlX0/i4h20iX4kSFO0
dZHKK2rMEObSS+cr0sWGGwZdQoyhwo2ItFivxBoGnwiJN6gvniQmWS7kazSbabrrwBhw8cqlLmeQ
8WaqrO2AeLHEAhptIei7ymy0KQ7GsCdq035b0T5VGFAXpmMI0mpE+NQ17/Zjz20v38DrCmQEu0fe
UBXszk8wipv2tdOZ9LDu0G4bWHN8eW0PF0TqQfmD6mhgEtyr6QhH6W8kMMWWZkbKmlB569RHqFEk
QuCvXCfhXy4+mKfAIc/mQQr2IFTIYyADIkN2g2f14Az8K9EXH54pkOUjU1eTstPk5jkLt7EBXPfM
2M/+sdXY/6OwBjtPRGoPyLZtvTKGd+KYrK1h2ZmAbppGs8iHQvWHM3ymJ0sC89S157XALTeaLztY
z6tFPnljmCvluRHsKsA4cjAHbwy8EmVMhqClCwDXbU1utAfrihIg/5d1Zfj2N6jflq4hOC/hlOs1
3lCAhQP30vvcTGN4NCB2Pt/sHXYP2U9VCUwJmA1nPUoFAsG+Fvdoh8rSCpWthSfrLKu/uPJHqNKW
6c2sA6qWvH+I0Svnt1Lc2qZinG12FMZ0ABbQftumqU1CYsi5VIx9Nh1h8PrvuzdQb4YM5aqCCsV7
nlq8jMW+96hiGoQYcrPDxAuOqMtAn45iVzLzSVUSZPFJGuJWHeyGGrvpdX59ziEudWQ1pQLdPfsD
GwSA/aa/Iuf684UG4i4XA1eQdiL3QxHE8RJXnQUnF/LF/xKhokDZz74WUzUg5x5xmXqXMS1n0w6m
O2t7hhmVxjCtxeMznGJVuBxE7ODXPBS/ltkIme0Z77i6Xz7HannUfODNfXe2EByKRpqyg6PiWdCZ
uguWeae3VRN3SXiI+h8aV2Shen6bat5QW3si0mEeI9RRhXW7X4P3WVy8MP4ZLLK+8F7NOaCvc5Y5
/Pm9XcOT9yPJ434UE8B75JXPMWtP4irlB8VSian35nhvjru5e7yVgAp9bIZONPNsY9xDlxjgawLy
EAXDkRRaHAtDEGeSxtJbvXNG4m3XI9zzhYQU4lTekUGa57m5IOycRaSzRHfX3bSQQMc1URgXaPaB
j2ww0KCDLJ4kX6TMn/jTulkF/5uhssvqF/kydv63CnfF0TbEmGSd+cwdme3znfXnxFqvGsagqx3C
MS/ImqRZrfHNR7DOknnUfsBe2h5+OPPgonMsp3Wo5ihe6ZsFBPuVyE7SWzp1plYf/PlPPKc4Lomo
2/o5U2XV/q+Yoqwzqg+wnHZZxBNbNVORAv5Y0O0YND/cxbHzF4f/RBqft108D/wkU4vRUP0pMxm1
UFirRjphYw1hAaP/B9xxttrY8NEiMwgtYkjnHNZdNnpsz37DlqwJrKVeIEsZ0oSUlxcq+2+TyO38
4xsPVO8hvgorGroYdX3Lt5uhHumfR9KntMd5gJB+/U5N/k7V3xzUHP0RLIzwHAyAyYR+1psA7gsC
suXJ70CXXuEIwOX+XR4WOdcDaGCzYaQ14dZ/kGsoD04y1QGlkush7naS+y1/wTp7vDsQRW29jCl/
UkTROVO9nQG6ATdFOfBVf14w/gHcRwlq/LgIJvtgt4JH5ybPl7d9/xnBSdnM4umJ4YKLZ3u1hGKy
ABBttSiXOzKwYNiXnp5rjcsZyWQfVDz4ZztFg69RdKrGAdmnowQhVR3HS5B/t9sI93kZs++4Ct6x
NBOHS0aTgaA5lj2NYRHmtWmTfP0KXBL3brtkbvtzDJwpP86pwwPtXyKoriiDljyO2QL+7qrlwFbc
H7DouQK48HY7aq6Ztu/vuAKRtw8raHspxmRia7TCQmpbLGwqbamIyTkhWGBoW7yufAtHdmNKAByR
g2efN25NV3Jtq6B9BUlGKyaIA0ncpW3BvciKD3kbGM5j4rHw1UXIezHqHE/qSoONGX7a7addYp7e
zZIbBTSuyPkCc4TWzkiXiC2Z1w/51vB0nWDhMHnCGAZCvVTmJGrAs7+muODW7SEfZV1esCLZ/WoY
t8mTHV/j9QBfN/ecV0p6HIZNOEg4DUrRZp7byjov9xudQQjYt9+d4VeYQ48FGLMjG+mcOLtP5z2X
ctCgNXjDYhHqxqRYjdxOzP7TzbobedpXkJEBfqLdCZF3plzDnhQp8sfqBU50vQlw7WAwmK8NZsMp
bxftewsidndaJP8oAK+6+FDF63798EcS6ciGzM74MmskYUTuenzkQ8rpnTaZhL/4FvO/ssIb9CH8
6XRJWlRBupRe5SD2pqMB81AG2s8BUFyJj6Yd3kNx1k70pMtvlqYINrWJHJ45niBu7Cu6xgKlZtml
dNKZej9zbxois3CcuMGpkD4V2Ty0MQOPmEY0QYub0ADv8qF3IB8aAoH0+3o67TdJFZr5r8L1MYcU
oHMlgEriiVgsNoKk0j+39TFTu0XrynjxYZMGgwbefPgcaHSe0JScSrIevh+hn7W6JC4MkyVVVmlH
NXnzEExdx2fsx6dzf0B63WOY25Ym6F/aBsEOix68Cdj5rY+xKr9WEmvU5LeFMHRownFbobA/QCF/
3CKNbY+c0n0FiTtep621A6MCnlCw4OFRuEwfpUoBVXGtPqDQWVe6Zk1o0JLMClkSkbA/yEpzXQnu
AhXIWarYg+ItBZ8RzIKg9hDxFZodr9H/oAw1xAC021SnbS3VNVdDigFjJazLG4MLFxZ9haG2pgLc
ZNu53CIYVI+LyPh0QLw0cgWELZhICKP+Y8AWmZstSb0C38rnP+1hKNo7/cY8x7HUPnWH6TbcH6jj
PjDTepKSovEyGNgkA5fZ7ADBNy/KwI9TU4AvhI5K2cq9sByK9wAv3VLbhgpt4RU0rBIL1RLrKqOY
k5vcGaoXwoh1Wj8b1H9fIFkwkrEzmU6e2Ho678powuyoX9t48rUXTIsPX1kZIRL2n4FZTj5bZibg
IfrQn7s9aqpxMUwYtVinlv5k5WFb2jg2IN56KeArbOYkkryKZKF5ibb+YuXplLbVxfb0xOKElmyK
NFzlKpnzEULqSH8JSQq3F01uzV3VOmx6TAZc130r2DwjNJt9becPJKANrcyemdXO3Y+Qt/9v9l3o
Rsgg54C91tRzXR403A1/06l4dXknh/VdkyISQfRdB8g9lytBC45sgONdpnyZN7JiZVQpl3xH766r
CXFYqXXyuYxcLvWzlXfeC+nFGayFFE6h15xGsQveKPTvm6eB/oLOimvTIbOIirt82KZpthmlD6xi
9mBkPIeU4LSf92CEGE04obLYvGItVRDmjSgLhvDABtzEHsVGiK+G872z2TqQY3B+QY2rCgjrRk7s
906rX+vp8zsKdxjx3A/1zf4B4mEUVTS/IKgRSUL1rhznKHCmwC5l25sOsnYeY39/lOzmy4Avu2Ro
BtPVDC04xqEIggV9pP2g82zHAU90u8zRdFEgRlL79i97a2ly1zarYp/miyR9Z1DG8nyzzDdmIa/8
/N2QUHa7oTOR3WSc7TVMYEZtLzo4Abs9zslL5zl9MKqW0wWvIDsJC9uswJmo36TmiB9t+wfLDtLi
V/e10gSG1jxv1PcR0VW8yS63GihXRvaqXq/5CnK4J71ATaq+PRczcXmtBcIDN93fPzPBR0nMZrmQ
53ONl4sEhlquUdik8d7TT1RPrpXyVj6rSBM1jt0NZ5pJhEP1e5Fp0gmS8D6/toML26U4OhvsgAdY
/5FHSSrUeF8bceGIEPWo0ObX9PL6GA8giEifw4AsKNpQQrKpA2nkbxyHVuglyVNne1dvmWiBdKgS
G4Lincy6mfu/ubGRYG9X+A3xr9QuegI3IFj/CQ4vcWu9x3h0MfE9dgG1gCP0dp6y9hjHrg7e19fr
RmGzCj+FzQwDMKZChApRmWDJObUMjgnHnoaAao5KptwKzf0OmVNp2t/hfY3ydFSLC8Lsp0oYoObp
QW9YIaFn9EETVGCYmDnZpGezwYk3LYKpkdafdVNeZOOczN9iQ2/4Ms1Oc6xqTtKdVncvfOilyEIC
WAhBnppsMg6ZT2tSBiXPoqANUPOhuHZUZh+0MGVmS9qgYrxldLUzDCNJX7aV7bZwYno22stjZ/v1
OwNATHLAsafGuN7mHgkj+ktQOXosXHO9klc/bGKpZR/jYQVryB7jqdmUn16jfmovkgex2MG7B3Xi
k5A4DQtnKzUAyszPannUdfPBaZpHLs/o6RXE2GKNrliV26tcZczBRQOBQJqV1gw0faSqPVpmmXIK
yp2b1FOCXLaz4SvVHe4cMsKItcHfwLionx/SjXvBU/eMHNPjh2UE1zav5MKWhtUH17b0/iZBADhI
zzLyTK6xrHxehTwLvXUuL/XsDM/UaUhbCbL2AFpAuBzlBF7+vdQuad2x08uFYXLiREXHJHPkmrcl
uxTsju2mh9Tk+wGqBNkhkdbZxYW25gVgLAr46kHYuw0CNveL37ngQGFTHroSQKeqy+oyGDf0S5Si
JbMJDO58ekBSIZB4qx5Mh01wQYv414oEFwjPXx0Nrm7CKNtVRgLQVnJ3siZYPC2WsHSXa6iHzgCl
EZcBPlVw1nz9I/IWrmYpwk4PeJI346tUpm3VedlDrT25QC0hFhX/QLI+XtfmldE+1DX8eTzrHqMN
Aw0sLIOwIh6A+uHvUkG0w2UiRX9zRwY74nFEVgOJPt7HMUXrUEKltmoXehoYaVwF+vnfVqNwdIxO
wxfYlLpedUO/2xwSYHTvQNCY/5YgAbAY8PQkB7z2u0cVDv+/4bk8nRfcVpps6l7LzHRIabrZzVR1
/XW0mzkGy/qNm0Xb8+awXzuzxl6M16FVqtsl6bH0+KXzz+eFtEBZkiM7xqWMlT4ioxZcmpAlW48M
2A+2+EeR3BWGJg68Zc6L0D/EUZH/Qc3S0Nr1NG5OSfLh0QEmh6G7x/+aKxJLFXzUOxtfqf1bdpyx
YA+uoPfw3ZfWX/clT7XXXDE3j4vyeSaaEJOWmOSndjZfUH79R7pRek6xBViPnnGhHZuMexJj40n0
CVTa/poM1rXLtOZuM/hE9txJ16a25R8bs86oz8XeyK2mATd296zvwoOu5cVJthqk6B7XpQBAT/bq
eh10ve8TWs3oT0RSuWdfYVF6+kd+wdSgtT559aLL753PVc+qCb/hJ8mfKLZdWNDcra2O2JkP0n9a
reBOwvCXu2OCFb0k2qrxMvs8lxcln42ahNI4cYAux2/0drFAeL6sR8ng1UBP8/ByJcp7rYClQPBl
mDOGX2P0Ifhngz9lj0aAidNDZgN9Q/e4qmTE41SZ+CuVBhWimA0orxLfs54otLN+RkX34/7TJ6MG
60ok8zZ93VLUH+imlV1nn00Si+lmk/ImmD2J8arl43BHvMJAmnkfEc8q8QBGzVbdKtedNdSwlRBA
2GL5sZ/wJ+9C+pROCP4do1Ch4S2OajiaN+ir5K6mI3dxC3YsPC/1P3kfA3FYOzDjGpoL/RH7/O52
YIPLMmCxuuJ//2NkBvr+RUfKG4UVof6AMYNEkNHXv2LrBz8r1fFOOC/DqxuLLxD82i6fjiFspqzZ
NvWm5q9SQUi1sWRV/qipRUI/zoWW1+OwRTO5LIJyPHotiN1aKf+cOR6dwNvTFBT69OGpLX4d8dzB
K2W4i8ye/9fs+xIohYcu5UQCXcQEhD17RZl4rWzheodEozoTN/aTrcHq2MRzSVaDddQM+bUdCQ/4
tlwaRi9XW8jkdWbacHrJORg2XbBCuOjzE6IlSiAGv4amY3yNLK7GrIKpK8cEhehlFp6EsqlmFDHs
mSRd4V4n2NPPF76nMDrLRyyd6sxv9yLkTfZrLw9vdKEjouw/tVGB6tVvG6tsOs/vuJkwWOLHarvk
QcV6CrxCI2I4RQFmMGr+u18nlGqOL6gkllN0e4vNylh1K7fPKDhDB+sQ1naeCS9fra1ntR6uCtLl
Y+ibfeQ2s6P5fzVlxO4nxCrUg3JfGH0uuh4qICk8g3dCCBm/1i8t17mg2b5dyJsSjZWZKTmHWg/C
pk1LlLSXsLEPkcB7d3/dOwrXZH92j+g1cQNnpfXn5HhMFhMBcf7yS3763wHVIrfBkCmMYSeVzlAf
z+0euM103DXZQx6KmI/GsxbcfL70cFj++mB422Gvjek40xjnNXuxG1sm5Ge7vxVyLOiaL8f9JbUv
coiJgLo4msIZZtAT/EsuMPaeErAj63yEmUW7A7lZlARn9hSE6N7TP9KtTN04pvpCrsZjlnfvt61t
3VLxoDa0aPhs5eaUH31VddH6yvAIHivrlF1WXZ5b2WhBdnbY1wfdvDBdLi8RCseG/t+Ms/KyAOiV
+wQ93kpV3R+YsbXXLa5SS7FPgyEaSvDUo+a3Te2JZRj96OgUFDgrgrayyATohMm1EuFPVLLIWoLz
OfzJSvvbtZLKcPqark8MsOrMoFeoEf4Q3cgjywEmItK5N1ZSmmXw5sllyxrxma5wSC71s35hlZyg
qhaDM1sk7kaL1orYYnl7VVuu1vpauImdL75c82uWEeskI6wAjpFl+B3no9UQ1BxnTT4HT8p7LEej
xrld/RsVVtu1vvP/7myu9SHqHERs9WLPvznh4B77QLnuTRzlcaP1az9WjStPJWH/FXqR6+nIvzx+
lVRERseB6PEZBhPTRUbwBKAvtfxwOupAVlI+HGnoTVZ4WM9ibTLIy+ebweDfFR9FnqwvIxiMyODu
3vYX15u3RpdSslz9mSWUTU43GgB//HtBjbHIKlcuV7R1baCFHOcp8IA1kimf7xTtBXUBv/DatMQg
Fzn1waBKwmud197VGNAefjE9X9rp8ZCDCddslZkh1wTOS3FgaQbsVlGMK50bHwAd04rO81zUfcvh
1RyJOY+Vfnce+ZL1LGWp14js/HOp1KmcGeUUxaO2UNMc50+0vP9r1MWRtvs0y1dkDFyz4RynuEpr
6T1deVseP9pgow2uVJFV0Ctg73On4jC6Ig6xrRgxJ5g8FrId/qexPqeBkKf/8Ik831/SpYJF5CXS
u9/6bbEjgzfd66eBq2ZzQ3qkw1IutzgAt0FPylFkMHTjJgJeI5D6pAiBn4dgSFEajRwSWuxvnw6P
xC85satbmEsX31Nd9IO5WyvHxAKqNUQcWprq2pQuZV07D8fZ79ZY9ZN68IMOc37y5Wd1+HubIllY
euRBHwd8MibdqhlcB8SvnqxDOknx9xWh4on69Mn/sGBICfiBRB78J7St49uhV7MV0gConVO7+Hwl
hkBkmZAoQJ0dOkO6FD0KGmDpVrtaKQlvNTuWH/w9JRLX7/0uWcsuOeL6PZ5iHi3+akhbnl9Xs5Fo
iDrM5LVFzz/+4+uSrNFNNm6au6BCi+GZesHMplm9i4fL3nLS4VJChmvLQqt0IfVc45lE+s66Z1yN
vHW2WqKLChznt0KKeMw/O26z/ZgLXxvV7LxU2+p6PCXdyrSU4XvvNBkGUxjfioK2ZnW/KRTxXm9T
mhBZ2RIfIE/27FEGGeeTAT01lbxSbKodmKGSV+JaorJ/e28ELo4aqxF92jmgl5GHoWmnvC5GD+Qi
b4Ceqx2N107gGkZRIcwpS6p4eb8840yDVHOSLOoAqclA1iCS0rSL26hVUmfiI9qU4Fwy7QNRWPiX
Z/tqbsr2XuXghHX92vmoRN+o6oC5Ex+ZL+tkRoX3APIKZI7OaZIlwZE0VzsqTuRnwRXyeemt5s35
E7WJbtJPJZ0RLW0LbMpRCEwOPXAHVzP3tl70rCMcBBXReR/34foElEtyi0WBy/bhl/UUvLUnnAe7
04KsgY6FGjzfOO25FiwBf90ZGaKGe4MfTlHNQ/3RDitfdLuWJ1PojRqdsjJwfVOSFeo8oiewy/YE
7CjJ7uvZPrDAbeD75y1wyZK/6ouwCgLaDCiSdjK+fLV1QL/GuSwZOVpAHdPe625CL12LoxoTO79z
KUgOZ48pTI1qScDWYz9Gsy6zkE04txI2q3Vt2n+cbjlleplG1mOoKVadzYsN8cYN1xjZs4CV5CwW
fIuah13Xi9jsEzK1GTtcRK+tnXzxteq4CmHkEtQeCEinXb53JcxB+NLrpcticsWhOcRVF6PFy6Gr
Mpr2GfBbG4rsbm3kYnqCh/JWH1Fd39tr7BqkjPcMoWafMtxuqRwblvgkdweZvlNj5eceUoq6B6+f
MrEYb17PZB6abAdoVJ1Zxlj7y9bv+Td4302hWadmhwRUnJMKES0q3l66Uqx0WrZyV0LgmZaZwMWT
3Ve7SN96vtmDok9joAJYCea2JYKU7JVfa9LoTGfYshMXU1e5VycyORUmssG40wOuNu58lGUtHGeV
yQo2waajZypZhRaw7jjkNpdnceCl3DdHZOIMDchLCvjQQUhqjICylN1lEsCoIxebCCJSHzTZRK+r
Y945t0gDvnfGdhWo12kW3YMlmenkAxtTrMJIE7cOYKY4PbauXj2xRR9g0lwJEuaHH8Nf891qrVS5
coZEBpWTVirzqUHJ7KKrpaz0JDyCMi6b9S8XoEyEAxGm5UX1F1XFoZP4sl287/V6G3wgPmoo3FPt
Icd7mOzW0AHAERwAIWHo2sBTRV0yONSmUnr0nucDCXwN/Qom7bbXngYrXP5TngKC6rVFNQZ6FiqG
AGF25lScC7iOcozdBUpRcoUY/4hYKIgdmkU4BY0OANFvxtLXdaj0a+NmcUsCQfYf+FEOJ40fnbtC
WHm5By7gBe5JoZbF/1/Q9U/qhOHhQ40v1bdGn13TVaHjWJwxb9wltOe2lHnhTf9Fq0ctMbkgbnrV
2mM11fSRBsK9hfxpcCNRGg4zpc+oXvsuy1JX69EtAzCYRNnSiLa/ym/cEog1ARXp+KBmSAT42eny
HeIqUU445N5p1NgcZbkLac3wt/loy1l3zp/M5ubs6ObZdPUqxhg01Kq7maKFNwnXqLDpgEJA8kFa
h4ppnQEc1EHRwdTHrMLK5z4W4aJFbcA2UR7TvUxm2pEM1w3YeunRKU/xh0LJt7lQ0YUEjvBd9rNv
wrRL+3dM09/E6v8Xm4Bsk711QRxfLiv2GrKkZT6eb6l+AcckXWapV3tQjFk1KabRQIhHQ4grFrJt
qjZMEMhT/ptkq5lDY8YlYiLpy+m7aM1xBUqNgrhH/RYx0oZ6iruFN1DFT2G1jLXzI+tCokzLjTLj
fPMUKCLyRuQrDxN2khKfALGIaf4IV65ON9A2+TX9Jv2QPgeK1cGQIXA1JCvxTSVP7w/t2Xp8sM6v
jJmo7Kmuh44WnBVChcBhH3IBZSvNBS3OacoirETxjG+eDoUnTbNrjXCm9F9vGeGd7SUKbfAvc88T
7+tecdoTVfqRRuj12EM1P+cTYwHYayZ92KgZVc+H8SnHiLPcXQeIvptYk5v9V61L+NlOT/EpwynL
9glNnStf0IbdmD/LrFJfrCKWfxphuZbhlpvn+k1DWwA6dUmbok7VIM8v6QmR/U3vq/upqv4ymtpG
OX5nF+RhjpMfbx3YZO1eVB/Jb4UqphH5+J5mYqDTIy1o9fGo7+RduFTkhpi73gyhjBNG/lmutWGr
uTSXNwppqzUgKCfFmMJC2UT8NJOtLYxe3g1KWBeHSkJ0N9XTvJ7bHnuQH61ckVso84qrRzA2Zza2
o4rm9BbqI9wPWaPNWJComL6KddfITQ9q1NxkZsOdEmjB04XyMmYZEZqdhLyHRkRiNhX5UfCfnqUY
XuWOxmTtgJJun6nJdP3FKBhC75JfWqzDQm369mtwOTM0PF0phTBJ+0MZfsQ9Z4ITfoWVZ+1+4bP3
2n++EIQ/FuIeT3VlvadCzI2M2p3AO/TpOzS+iZNxN2kpY2y2aBwosiSYYi4jze1M3g45gkbHsTfj
Np6t+4V/YE0QazSsy082y9Pvb/IAb1HEuJ8S20zu/GNEwJna+u9ThnxYgbcPf0swDh4iBzDrfFM2
U8xozUf6GQshaV6KZ/nlGp+TdzgG6BfVvvKMrwkvUpCm0SEvsqP+vhr1VHlCuGOQiAUP2Rqxf+Aq
v5uGWcbBZt8vCQhUhKdHhOhQ6sSCQ996enT8j4u8H+yqM/DS55gdH92YnDHV0KeFO/CpyRNWVmuj
rqWIozPeZhZQhQxZGEnAsQWe9klObvssoV+MRj0B3ClCiABv3tg+3Af+hlVhWzvfp5rPtOSuyZGX
ogetXqJKYLluC4iPiR4RtfqQSu6hpuBIhgbCRYs8OvgMJbhkARGZMD2GpGeiFEPplqXK9JQrceO8
qu4eZJduMmaBZeflpS4u6Q8yeB50R1WHxV4GV8GprOYzZ+nk5WuOOo/IGH67BE//oM+a+f+fnWf7
KQfyzfeyhlp2yzKhn/bHn+GWVAFEsxcmiLfW3c3+KH8gpjRi44IKLDG68w+KB3GEdTp2eNlqLrUQ
QMotlrsTZi/Ox6F75NCJOT3S0bUefTEM4bLzUVSaZSzKpKf2CTV2FkX6rX0/SelO1tQ8RtpzbPO6
vYkhf5gIvqngcSUjGH7Jx+RMrfKL0Im0jaKPEAz4au1iOQnTsUxtpW/8e88j48oGudBRkl+ANOyB
dtzL0moCn/Eqyd0HEaLiq51Teq4IauKvfkbwpkByD1eXqAxwoV0PLdsYZGto11l6+owSmfF5mpS0
MPhx8SkUlBJ8v4dsaOwUj8iQzueJcAl2qNzWpQeQbYn/t2q2afsrSPhb1JoCouNfQL2LRgpVY+Zv
umGWG8eV5RCj6fjC29IrwZWY4M6uS+LhiZq2/9/yvu8J6HK3gOAsHUPjrBEIkPScsEH38A81nMWP
5r1aPkuN8OGrmk5XKeu+fZ6T4SkwqgMdY+wb8gccAKMi6RnTOCa+hzbJl11RBVqt3Mhfg/QB1aWM
tuoT75i0nEDOtStakXg9k19HniN7g1BPoDVZVMU7wgcVDYK4XaNJeXXWkhm05HbxtrDGGZBwvSiV
C1GsjZQt2rqhHW07GQN1MoopsxrH7QJH4a/l/BbZxC+Px5bUvRL5ZKXiMBR+FOhTrooSKVwnGIm/
lDvY9gGoiVwBNPOG21EaptjGEEBZXaldIl5SN0Yv0d1K8toINLt21I8/9h3AI3Xjr3ESOeiNPjB4
bEXhQQfmAI2tal+3JccvD6/evMWMHZk3My4+bnPt7dX/Z5I/BrZp2zZxgfa76sj6dGY1pY6pBBn9
RoM9Z61RhNkZU2NVgbVXQD/0KGXjc8Lm8q5PbG0j2VLXqEsg+VSD8fDbag3hKloHqQJatecZ2mpM
ztvd1qE0TqzATgzzWRPnIYdJff7BjTqoBhI+piFcwoq8NRjgI/T1JnOrXVRqTYDkSv8iCliIAq8X
SeqC0ONTact1KTfQuF5GtuxDX+vG1c0qh8mMvIQ+3VmtfrU+Udsb9JnMJFQhqxxA0CdqE2NCWE61
KetQ3A5MoviRnk2xihxsYi+8VTbkPafctTbllUsldEo5hmqJREulxa/OVM5/J8O3AyHvAAg4xV5j
qWU2VLObBgi288ca0AqIcsGRXDVOFuPEuZ1BrWId+d3YWEaP9KZ6AGmS3BRGiy9HtHHd39vQ4YAz
p89FeIk0RlQs+YMG8mvGih+5yJ+zy7D+imHO8QOvK23s55h/188sbwMXrNrqExzWS1xu5UY9yCai
FkGT6ctdNzpVQkULS0VTz17xD/ImA/7VamzeoczKD2N8ztJcHF+mbSGKzALEdlH4KQ2+NlVhTYj5
JorNaMOpS5V2Zix+5onNCFDBYW/rb2N8ASXLwFn26NF+EOQiL/UgkOy++mbcETpL0PEWKiDOk9V7
SyEyYpVG61PFEMBTiqynlerkypVunuxe1sDIfE3xF7axHKVBhTgO8Wu4qAl3ah5scc/so5GeWq5e
Eh5xSw+u79l0oiiXnCo8i+eOG5fD7aTxCQSu0mZNAly/ytf3IAUp7E08MzZvZU6Sp5plcNm95tan
Q3YVnp3Et3qvbRqlYhNexM9c5TBk6raFuD1DeVUGyWspOS875RbQ/jgJlj6JB87/IbYPXGBh7GvY
1ckPB5WT8MBNB49Y8EQVCtSVbtW70Zmu8XgvqkG+cUBIABrsiKXlsuEE8Gki5eWEpnCTzeKoej1W
Vu6cgqN5/QSIz6PAerzgAQDNWXWsAdze3SBEq7OShe7zuQ2rwIQSPxOg2FkyeR5zfl6ohb2bO1Yb
yqLHmvJNyEQbVCiyZAnXYDK2AUWtLkWNil7SE82evfoQOXI05iEl1aiJk27BDI1q8ad9yamR8Jm2
WoSAAM8tvwJ6ms7SyYQyw6cZMAHnUIPJKbIYd1Pb+YIj0HGsYCe38z8qHE76ziHHzkD7O0IYJZ0m
uaqyNE76PRAgIdAaY9uFxg8jEhCDzfSe2xJgbnCprzT2mpf83JH5h8fEi4QJSvC+WhDl06tZc3MJ
W5PToF+FsHS4PKxl40hwddo4wmJecoju9gXTvdZ5f2hPy/Sh3zpzW0Z4polbQKcXcVW+USb3Z1Zq
QLXMBqJja+heLAPkYHpqRHHmS7G0m03LFEgXLbc/FeFp4yzwCONuwvhr+puhVJOvfx0DQMd8shve
uNeMuSHpv+74nkz8NSX5k8xYfbWYJN93SgiJ+aD1i52uG9vxltKM1SQDsKiOGjywR6yFpWWe8seM
d0npW/tR4LaaUIAHTaSJoz2HBeS77Ev34OBcNjxGzj52kYk8fqhv3rHTpRBgmj8wxoA2u96BVJMx
XASd6G8KMmbd8LaY+VA/Ng1hiVmRDlHqC/egmaCamEhzVVPf5adCYsvZ/rtumL2lMSl7cQuIx+1b
eRzKlrr6Rra0ckj0VTKCGPQNp8AeKH9oXHwqjJakX+c8YV0GAsSXz7xXCsoDjEnWtHi3MWRABw99
CVeRodr4ZPDqE4We15FwrP1ketGBcEzNHx65geD3eH1bYC8CUxpx42SnQNvgvKnsqWXSI4l1K3hl
BSuyYmUV3OID60KNxxWqxDT4XzdHATug3vNs8zwdKUwTiqj8ECaLoFNZ8FjxcD1KzVzn1tfsSxdq
sk8qjwctatWQnbvN8xmgE1QrY8GsMpS6gmeWLqurFEmR1tQ5892TTl6SGYRuslshBNiTgCPpJiwV
2AwOkYFBKUWaGkirFs7R/bh6XRMPwN00L2JbfdNY9sV5OWDfXIF2W4glao3RDsAHNDzbUB9aARiW
PhoJQU4/WCfTXsTjcoH8233oWjFxZIcW8j0xzibyyn9j3msqpCobKUcE08gm27HuqKdLL/RPnl3+
JlVspdoYMAkw8ixfgWpSV65/Kg5rBEfKK0lDS4aJh5OB7CEzFfnzRgZu50SNAW2j8qWrf3wDtcPP
iEVpcOUVcEdCGjMSmH7PRdAAjtZewGvAA0TYuqdN8fUP742I44dli2GK7wFmqGc06FV3Usb0Y2lX
zflHw2V2ZvGjk1I5+OJN6MZlgVygxy2055QnkUaxsCoxozzLVjvjj9DV47vr7eEEK4gKxmbM4+4D
H+8pot8mr4kiKvGsKhDY+rtcOD96Nn0mm2dybAi2WK1n8308zzqT0xk8W8SlTMOn5Re3JHljnUDD
IDStX4lNR0Q03SVZZYNvlYHR+Ee/ErpwAopgxWoNqPnsa3b8cFwEbPBeXqKdSPxUOX0soWzazDxq
I5RGmyYKqmA7TG9dXyQ/m3d+s5v2JsGImgwf+yNh7KND4hKANKdA2qbNgSCgQiJGk8phqIQTSt+6
idnK7SyZuGlMnXdO2/fAW3cLIQWh2eGywDrAMmzgHVsoF+KPopowzbYRlK4RTtAQJIM9CVTwlCak
j7LKEhSeOHh6AtseSh11PrLojpTSwZ45PSmaaXDBLtKpATRyydXavkY/qQ2pY93lesQ8X1tyGfRP
+9cVf1pwrOE+ltukjFmyKghybhFrVE2EPQUm2O4NMkSM6l6cN34105qDLV3Cjc9SCRNWgGSqFIdI
jQbXmzkX92o6Trxc2LV1O7H5J4PGtTXkCnZr1oMLoGhzvpHPb13YiaHOSvAn/drm6lXNucvKRIpJ
igxAxMewcvE9uCtyYUq8B8EE02LHp6TkvrTmrcIfj8tCCoV2qJ6A2MZqq0Emcxu/YI+tjn/KLIT1
SuJbmJ527QZeSS7PqJO/ShljecKjnkvv+4Gk3307tD+0f66Az8wbO4SKqoactfwOcTEDWYNG/+m2
25fXgU49bzi1lBKqTmgpm/cjC5MvQVPFwo4kxvWNH1Ox2jA5mKd2N9AfSP2YVlJo82ut8+MNE9Yz
wDK9iaZ3tfvg96HBLx7L37tMZ6jHlWJKDaBK+bM5IoHHuaT1sst4DLIudDo1JlYaMR+soHX2yNhw
EZWFQ9zNeQFQnqKNO7AHXQ6vJd5qhkVwHFh3O4W6CVEtteVJVqKFxVWnXBqrJe7A5aof2Guv3HOr
Nh2iDc7TExfgAofZYFy+ilLbmnFRyiIYj1MEyjyHvO5twAWZWoCctTWqrwbK856q+59Oph1lQHOE
YHJgnnp691emzsuEJX7X2XA1NoknQMJFQMYP7YrrriZya2X+x8VVYgEBE/nz2npMMtGmkJmS1TuG
Z/Nod8vCdAc6TrHMh9HsylmeTbPtzYsx/8WbRinkY2uh2lT30N/zLCXpxplQpCKkpa4xbh1Ci66R
WyaZosDbgIoXOFIvDRVGdSd3xraZiQGpssno7TpUQGQI5ffHEUbLDxZooFaXgNhghOZMsWaJDBo9
aj7w3uIjPdF80bctQwHonl7cM3L/XnOFg43eZ2bzwFY8tZS/W5hIEGzuD6sFKNYqEofM5ShgrHGz
vri9S8P6hsBFMTliE9p92XACHrQz3IWZGUDnP0rEtcfhX6ZUlsxvsS7Wnz5XltMgSfyx0hcuir6v
XiAolRm3+LE1z0kP5PysGZ44sdXbfwr4YII/OGbUALsy3QfaCVzFA+BArDnyJtmeUgNqi0PF3LfG
+KpCY4yLG1U8otrB6VoHYQh9/jIZl3XzGX/dD2UQHc86dEMXHdt8fiMCg/GzkBskTr61kpl3XajY
/JrolekzKmoPOJETc9SgDh+/Jtc2/mcvXRmqxE8x+q4bAXfpgUuqGmJnZ3wVIMHnO9oja21s3CWE
DWIPyPueeCC1/JEC9eSwtn0B0kBAy5xWeQBj4YVFiPRCmbxXHkws6KKsSg6JfmY+NdmIqwj6Jwk+
qu6qJ5wYdQywPlNvWQ9I7fkAo7iJZ9xhPj9o6+bEwoYKYS050E5bAN5hxGlAVLdLOr2qZJ1c8t48
xEQ5eoQLx1z0+p/0EG+6UW9wx9kh+uaOUkDHH15F5wkopWmgPSUzuOtoCOpPCH4rzaAU8eMtIUPa
N/kLJmR4mciVl9a5JZwhefsEYQII7ZoHE18+IcOieo17shuzgj+3jsq1NCJaT2Z+rsMoJYmmHlX7
YwA3JvQMpGoljva7V0rFSoPSVKD5/By1mBF8hGinp0Vno3v3DWl60w1h8DMANPaDlFYTkYIwVFod
hH0tllaI1W4r1cspkv0Mi6BDOlgUU/qk35Z8iqCo1RDAydTpdvYIGXgNgkbNs9PRW7z6jSv7Fu9W
q9hPMzo4ZvByTx+iAL0BszNaW9P+rxojyIpUw9DjsJYAuMWHMU7w3e4NNsJLg1v8c/8vhdS9I6w2
rexwzLSpzuoRuuDVCUR5NUYBQSXvPewoNbxnIKYIwagPrfJzzmIWYCgY4gKQ8LwYTxjHXheBDG2w
v5OxeyWWsNIturNZpaNFbq/C0zMMLGWivcNk4bitCk+zzpDA+jmvvoIum8zV7cr8sWabFS5DgLES
7oZFBufm+KEBQ1SRGoeTaUBhnWyKL8O2gIABmaKAcN1eKqKYdYYZjHnDVGjmpEjw3tRV4hkLyWkC
sKIeBpZgpTj/CeqeD9wW7AFVaTkLAFRomXTGcCT1k0OdEIvQzcAHXY3d++05QKP+mPVlIQkKv8Uj
ILwEyzJvTe/oMbeWfZIbgtw8FXIhUOMCV7H2XKGxRaWSGZ14xiQf/t/7TuT9t9hiV6SgAY6WKUIW
Hb5j/knfjfYahQsQ4OoLt38iaNG7Uf+3HrW/EfVQm50hfsSw1LkJguVqidWQtzYWnJWW775D4fii
XPVDHBn32zT9FFdNkWm3rVWMps0cvgcihWls27SkN9DPMXYH423M2OPRPoqXQTMZWLlVVaoZW5ST
KSKMApCWgkAu7YYxLjoIvFm36r2chw6GySGeG0Zqv9cKYGQgOhvMldn9Dd7zOqDcJkzyiOO9XIQH
UqglS/AEZ3tkyeEArZSkw9g7v1Od1WTWpUe1NcG0EhDxM0wwp0h7DHWPmIXg7Dck087xquxifvP6
o3NWQyykq0UTAmJD9ZDYguFXwDAYijZ1I19zPP3lXQONMl+RlQCE4mX7l2LLVZVMXHJ1UW1Q8iMB
UJjwzmhbnvlWzT+/DtQZY+c9Y8D1huJB4gE8Y6B3tWBPWMwk8uE5hNFwlxSrRYqmGV0YpG5RIm33
rLBDsF966cmm+A9krLWdNmviX0dW3uJ/crppn+hP15SCEem2tcuhupPmEB3La3TOSvEGPLZchNxl
IXeC3JSU6HONO4oh3LaWT5LAkZeWw880sJzYF8+euyS6aahpXRwCg7o2Mi9TwhvY8w/BDAROZIY2
24v8EjvI2nolkbOzuPKuBd1mELAplNEMQjYk3MJL8mqHHSpYGXGqtvAe2hnch5mu6r6vTqkcKRy6
PR7HfsAz/72DNWM1HVRgy1tFW0W9sXYtdg6w4OLRRcl3BFU8+n5A9ZRvQGjRuvlstrYHBG7e12yf
09xRq37B0Eh01p/2BrhI2SxE/RsoPIjEG37FJUUVSVfJAU+qwtCJCqIZuKLqzBkhzUmh2m7/A0I3
IpCrGxAuNePk0zZylZc4ypqXU8Wqru1imCsLgItQtqXHBqEPrNVGNnyk/DCgHTRxy6/JeHoBc8qu
1Sv+1lYiG0+w+HAqXgjNRZlgIzYBHT4LOMAylfRk4hrd5jAO9S/TtOABHF2d8I4Cko6J2surDGeN
fL9rl+1tgmH2eUkLTS8HEW/bMnPac8cN210Wc6VSx07xLS2OFq0FpCWX0j+oOdHe5VLsjK6ls9l+
L8FdwWjVmluARzw5LmieZiCqEt26gnd0k6US8Pc5wmqBedKrDzNuqm8jP8/pp/fKkbkHofc9opAL
6Bc5T80cPTp4tQhcFrtzTnCIn4dPmCe8dXr7b8CXDqiTcrZYJDcIGVlhPcohu6AMtskzkVbbUxgk
assRbk49hveZ16elfpPEtTeHt6/0TFyJCy/mlrvendM0q3cwAdQwep/wu2NW+dvF0jD3RdRammSd
WAfw43SGKpvoJRNlhCI/VcRfsAR0naUAFPF2mA3c72rav8mZHHJG/lYm6PMCUqYn3v4n5xGvSHA0
dBXO3DLOKBtNLVQ9PgwFSt78ekzqlWQOt53CAh7cmu94aTbxcnrflZTVK8RIgNBibfyNil8S4+vL
jo/prrdGdLfGr/xWYv8/kk4Pjizt6He4ZN0Rtn2exU/cx+MSnuzqJttrAa0xw9nLpTvgMYJojc9Q
/KVO7hhxM8u/WDil3VBbEqvE5B1yj1V+ml1tuVNruSiNqq1iF3VDC7mqW5BA/kGdZc9FaJ6Q3GEG
oxgwtKec4AOQpKF+IW9hNZBgfOR9Y1BpwtYqbzxknhpfmMkuEgePDoO9eQYeHEngtPlP+G8WJpe9
162w5rdsP7yMVXB2xykhgE/PZW8FoCOTW8IwiyZRI+o0fsb+Xz/Ez2N8VjOVzxjwZyJZyNSgt8X6
wYcctFs6Ipo0gXrXw6+oNqmYNDEu8jucz8+qj09A4YRW82Wd4vR1qgO1Rqucw6Ry6Szb4WddUh+G
sA03GApDZbEo6wI8RfRzvwUbwheqxil0cbwKc0LtErW6SVnmx60PO/MSGEq640LO8HWN3ldlfcyZ
6+rwPTs2oojSfq1wwpTyx4dgX801/jpqY9hUiN2ti4bNqRvChTeDuChui4GHA5XG2P98038MUSL+
xJJJPG7wjZ6DvBJ/HhQURx5IdMaOOLTAIE2736NVj4sOD1UwadOLHYe/O0NWqayEzsGFVxTaL1ed
vGb88UXY4E9NKKkUP+86258EgDhHmiiuDcuVCh5PAN0ROx/sxru9abES91Pm9xVZxI65IMlhopRz
LU3Wwxe5RIjMjdHec9Cv570I3o2lUvdoQWhElFgcKdjDRmxjba8tcHb0M6hy+etAJSk1ZoWyvW+8
wd9h55eBFyFPTE/kmYkEukT3u926NB6aCE09DuUj+R8XH7gZMIlEL1gbsjuPulOXAVcDSzELAjT4
l1Qwxepy6Wcz9D1HveWY9L12qVvMis/dYC9aKWqQwz1Wficix2rNKzwE76qtx2qFD0pFcephvCso
7/+JhisFjj1yiher/W0IgdHmsY4INnS/HbTr6k2zIsNd0MRK41agCtiTUB1kKPZkX+xV2vgmIQrF
j03ur6Lbc/XKYJBSWVanj/9V7H/oZYEcRTLs6f6Ax0G1Wcg1x7XJG6wyB7+Tc9vfsPLiZCp68AG9
330oC/jDx/O822G4RqAqm+PbLFX5a6+v6vBBab56M0IYDiQeD6CVA566DnUHywuVTgsO4gXZq9X4
9QvHI5G5d8H3FASpXqOefjec9UeA24nxgA99DZ//uq0pedkV+fTIYGFP8+fHYqPIl6eLYaLj2HT8
2PiW1qBgc+LVRiMPtiYwlOc6FMx3/myE38g4uhqIFPE/ANTk7q87VVMTAH4Kw4LsBGiJv1iD8CVR
1EVmy7O1eV5K20D6sDlSIMaYValTOmlf6LErOHVlUIm2H+R3HQCKz4WeKDgFNSb+NyeNsDJ0zJ0t
e+WnPuoBcHjBMyhnc7wC8HHSlOsJ08QQu4fExhnpjkrCoQZ5PSk13Cwn69XFQmzdm/rSJW5POrat
+C8ColM6uhkKP1MpeMTrxZv593uafMTTnPjwOPf9UC+qYSeB/5caDgbZilfgo+ZU9Hg899x1rl03
o1rzxu0MeXDZhMFis9FMQRW0dbddRREh4T8tn4ttMyq+LahgehYJ2cyxe5LcBTe90A/sb/5K/Fq2
iAw4fvJdKSJEVoTuUIOEHXHdMMT+wg46erWodGTEVLmBFxkB/Im08TgOmgu2WDX6coPcQGm1Z3TB
9apWUbKx/gA+B4QUAOzZ1Ix1dX9ouLTDa8qYBTNq0suuvto5F+hueX994uJlNqqbr8+LCXDotbZv
+s4Mr4o1CPsnfzfr4/gXEKf/Kuh/FsSOh+N7P/rQa1OaIgnzAa5KiR6tQsQa9zWcQwLXYqvQfQrB
k6lMzDddj+/oWuSRxiHvQSW1REw1w8RrgDFpZdUXu1ME67hsIzbKKA9e5W6ktpCCZVCjl/aklatA
yAPveqvvdOhdzSr6JRGOSHJLjvdTCq0lIx3Kjh+NyimjHOs2daPKLeGHDZMCNrmaD6GZ03ARXysL
xW+gMwACTl2zmTXJMPOWvDAPDHlZXI+Us1JYvnO+47/eyUumerbCL9/xjtfgeB9ITMcHYcQkPCLW
l8Xh8LCEeJjUEYURF3dZmiB1YnfO6QHqsrShGnF48HSIK222/3QqlirpIGqHHGX405G3z2dJdNwC
PZ5yBa8vS1WlnY9wqjiym+nLDEZfJmYs6dH1e8l/nltECIGPEqZm+C1m6QaNnzMF47X4xZO2bXQi
8sVcAGpVhGKNtLUZI9zuo3QoEf2Q72t/sb2kX5vlhY7tk4dgx250l6NzztFi29JOMe8eQrUoutgX
mW6yM5cLmh/oMWq0lkgxH77L+YG12IMVqyWGT0ZYsafcv7kCnXP0TcvdaB760B1vKL8qzIXQLAAR
MMOpvjbMf2sIUfnPu69NhVJ1bQGkF2720WpLsBCTxpxb7rr2bsHROw4LMEyxGNb8kMeRDjl+zkvc
LxscYam3axW6iFePEXsCvhDxhSwyGcXxr6IaKr6WviCX5bhn9lPGyDDxqESTZXbSk0mbOoRMxSP4
kAU2OTHa5sRqUUWZr388DokW618X5QEa6J3dqyJuwxgvzR36A0JeREzIk4Ygipva5Idg71zmBD5P
2tSPZxD7R4J4A4itPSUtbyCFD5xurhue+CwoJtlNo+q99n8UM5gt6HH25wKDF8N5rpdHXEmbm+h0
gI28AWJo9HF4CfJS3rr1DafKyjBLSGPfFIRo8ERYsVWB6vlFfm1avWMsybfIkxtm5yT+VmPo1mPZ
yTiTCkC51HNVpd3plRPsrIza0GP4ua2J6NX0hj5Fc/8qXGj2/ogwXryjKehETc8391SWCcyYaBA8
QwIRWYJuPr/qouAYIZHVDrInKoTReI2ahGDGMw+2lVkv9fpklOUfPcsLb2oKxFVKtcB2pXSQdYqB
LRKXJ39la6vcKkedxE77MVITBuk4Gen6mUZongKDEYwCrH+4B0dz70mHrEWjXqp9ngmZH9tejwlJ
ly9tPG/WxQCocRNiJYgCVUFwZ1O1LgFR6nwpvHueqwtL0Yx2Rmo/wSgYbVjgogoIptHhzMoD9pzs
U+TzVxg7pm2tKewY9LQ7N5hZKQ46zF+aXw9XmFRWlKkpOmGemUTbHKPd6fZUSxZELriUynN+ddXb
GjLMPpD0GkT+fbNW3oU5it5F+wFJqFWFN0UhX2oSTEEM6weBQkIE7lAgOpiB4e2FcwnVUWaSwHqU
GYK+JpAcI7TiCJIhXuw22wmXwBN5IBi52bXgTaerR0s1ZhmUE0fR+aOPlzk/eKgC1PZ0VZMQRTTg
PS9duUad0q4BDXbrBncsegKw0BDEvfdIFLuuErLqKAMYUMahDiNBTN5exmtRQrKuVf2gltyznmX4
MeJAfnKpZXVlneM3fTwTqayFj0MnWedexLU9PWM7X9unKUEC8AOiefRPc9Q4pXn7TB0zlCDLc6VH
TtOF0s7G1FfDuydbn2runUlRbSXgpJsttMNayf6cxMAUKzr2pAv5b/Qd0i97qDXAuC1/TGjYngrz
yvGz1hV+DOC0SzfdQwdiS9SMX/EmGuzsnElyi6kRUMWvO6q1EpVgHtJa29WDxyy2JWQeydzpAAzk
4m3uzZ8kbETAxmG7MNplbSQ+JfAZVolwRfPk1M6xnuZAiXGJmhJugeUWt6vZfvfgCsFf4u1m02G5
qPURDyEsuYr+rOELiEi0bQWSajKXTmK39XJJSb3+cAD8NOeOR9AFm2aJiU2MOaJYGNT2uf9ord7/
UfZZyF7kgIMaUNMblyOzavLnuuC/Y8+b4MXLauY4c2sGiaICRogV9aRsyArcy5pdFgu6p8ws2PrH
olRsO5UpN1E9STeZLXrxpDjHAvMNBxTtaFar3pvlqR9xVz8tagUh302Dc8+yBOAV9furxub91inl
H8FphsGNaBNxPHzPvXbl1jtx9ZjcuHIrOYlyt+cfnFB01bKJ8eIc+isltxDswXXyNSOQWTAzbpGA
Zit2k6NvYkcmE91KwL77Rb9SmuODK/Cx22NgYzk9Jp5iBDVAx7ZKN8YjUpean4I4at7uai6u6Pp/
xL0m6NMPSlujU2w9KUksrjhzNDBRolu9asEIJrZOiWI4iiy80vOkynWUeV4vdSS2980V/OMyThWS
tBlG5WZxxJrZ2meZMVXYwrnS7KxqRjjLXEQmIoain+bkLh4yP8TP6hEQTisdD6jhDxxuLmTjVNAf
v671QrtmEQbpMKGFBXKdFP1/hXmplI4bChkQuXSIW2XL2gVquuvgJWDtz8c+KH3C6jj8edzJqK9U
BRuKcAxd11YGX/SWW6wSX561xTtTeXv3p7kmVJNiXY5tfa8hWL9ekDj6XMJ3Od+8M6mziBeKaA33
II4857lSuYoAhmMt1HZu8CSdQwlU75VtIBHS83vheR82X5S8cf2lwJ4GwqVIkM+T+jsp3MVU45AH
6WIS6s414Pp2ZqczGqc03bBUE6ZCGvB8zxt8OFT7HvP1Fo40RizSc5lPgWypAjPSvOn2IvP1Pt4F
3agz/ht7vIBk0I6dnIFQzRq/N2VMtodNzPQhDjm6aGYXBcvVMM8Ce3uLLNMkjzieA6U51Lo/0aoL
GtOIhR8yh5yg7oRnJwY19K+CuYK8H2hfiSn1CeK/oIaXJPvI63qhBVQDXrSHjKKVRAfPbMWK5yyi
C6FYqbE5yoJPICnbRO9DW+CGhNaQCyGOLY+UP+ToVi79n+eSpA67SFya9ePJqCUqa6gK3Pbh4oLV
sAMWymrdkCLksUimBBluS1EPwr5yqrd6IWcu57IcwiskLtvEWPH6RVYsS4e6ZUewBWEMijXhjAzW
U0iS3ScnCjocjC1Ok1l7tVnFP+Ae3uDDponoIvIEy1FpNgC2Ls2VuvTYRQarCpeSU3/rRV+c2b26
18bKgJjEsyxpnKnCPytJOqAQmynKN/O8bMEggmSVtUpt9/Y15BQrWAgvVfeL/hgeg8Ve30cutXqX
7FiDLJ55K3xuWSCUHSNs8g+YbxtJdN/03DBNuRxPXgi5GrZO14GqoYJF0c/xbb1n13LA1vHRmUsJ
VuHW3Hx5HjA7XG6zUZyT+xK0+b7OP3POpPG+3aoADW0AODA5Jb+3sdZgU6vyoq5Nkgg2cgrfqPwh
IC5k4cMAJg8adCjVzv90y9wE8dTg9+JbBCewZ1NjetsD+uqg5LeObcXZ+QJfPSoyMWUA0uXjO1uA
LgZR/472tiLTP5lb6QbLPK4JQ70aSZU3ZlkZdViMs52GNXildlpzsO/e+4qL5WaFEwfIYdt3OeTQ
y6Ofkg7XLiXHauScw7/wOzH+MTI51Bn3rCG6GLa4g2slmI/6VQWkXKUO8WlAWKrw5d5jQZrkjyaS
5PCxqPtvmpQUa8ZkoMDY/LMGkdEMtXR3SUUlVZnxUSidFXwn19LL8FgS3fByUF2mIG3CtWpdZTRL
68/0hPheoHfDIB/RBczNQaJ6lEc9zyHcq5y0vB+IYzI1lwwPksOtsdRkivBYSUowgCE2BHGSXi1+
cXEHYvo6l0eFZN7jPL2xh6n0ehtHH6k13Js4WJA5nrXAbmpQ18z+bXbA0ogwHTd94MvwUsj11LhU
u96SyniaPKXlL1SmigLiCESMwOctl5EZGWmfmTrrvo8FSiE3Nx9vUIiNa5QVGlMizDCVuiszB/VH
QRzyn+VQW/W0FXxWlSnL9FkKHxSbD5BRzVbAaflZ5CG7LioOWVLzUmGGTbfgWyz95uvwVLEb7+8A
doqOmRPzhmkpQFlHhxPh9sppj3XzhAIXSLfy6pgRsdH+rDILh+kK6aUzwQ8Yehh3txUXcTcU22R4
axIiY1CeKryCFmdgFlj0Pumk8L3ZZWYzbXnrKZt+U6gnMd02Qr4ikPTN40dKsmDpnF2zIobNMq7o
ZjKytlJuJLNYF7pa77p8QFQgraz0pnNznb9tpr92WZE7Xu7WOgKfP9j0dv0A31DL/LlckwufTvmX
fmXIdxy1D0Uj+89jQR8sUgurzcIt9shESqPafcTelq23QF9afr1S9k5F9BN0Q9vT+yR/jtYeFe4N
kcvJKx9Jsse2mTNfyGEj3SUIfDk0Be+RjKh03hTO9lT+wTpzEl3zpDTPyvjkC5XlRvN3pdgzEL07
52JjJfJuBWiAAOY49gy/w6KcungmOMgWQnJ/U7xI/W4WMElz4PP7nXCHGDozmmWFDyjTjQGAK0fH
8QFIWBock1n/bvj/NwNOXSTFc0V4B/uc5KTStCB+/xXjdlUx8BtgAJqvGymve3K5OhHlb5VChSaU
fCSmF+dHEdWImqIv6cFTcp7xT9IF+6f5G/b9wkieZaxy71LsT9ClVqo3nKPN5qfKlkmbGULaCuO9
C4amNmI5rpAcwkX7TIEHGbfGhV9ivuWhCd0VP9ytOAoRWQ5MD1ueiJlgb0K8dDVx9P0iASMVG9Aa
bnjJ3KE+JnTZBmp+rPpqPkVWjho9aC/CIkwDEnxRfKku2W1HSoKzr9FSIITIxN/DzGLnVZj4OHMJ
VRbw698NDkpejQV58mmmaPKBPQUiMmAvwrN/9RCBVUHUHdIxCmlkCVSp/LU5Nwc3GA8+HYtBGYNS
8hnyk0ShHVI6FCJNoyKQs0Rn1hAco0wedCrsL+yYJH2IA7LOtTIGAc2Ug0yZcE7jiWGdQdcUNKaR
9Y1riibnuTWpodKeOaOCNUMqY4C+OkHsFJThsYYQgqTLpgHFoiiwPr0EkpMPaqXK6lwHzL5SU5CN
HqZcuShL5yI7dnacQKEQXi9wdAxa52maAsMQ5Aj/E+wHDfuxs5LN3mzKS8vOynOMIsr4YAxP4Q+Z
5K9tZmXT1C3/5y/zgnA+lLZ3u91Loj+Oa0IU9yN7Srvw1+LEg+VjmftlE7EWSmI8DOQlI7V4uDtF
kzf0xTRjnFp0+ez6UKdMhb+6fBcBG7utIb9YPBLi5UgoTTEN4r/3ZznX8c61JFiSMbbwjDBLVggk
TiCesRqrKLJIJZha260uRzesYzPE1UZrfvKzxov4iRskGZnzcEtkpy3jengdR5y5k+5/M2n9uzrV
fVpx3sqH8jJ1vXbQa6CiQyDOL2gCEwlaSzkAW1O5ubTW1hDfxzhyirdOxhid27/gF0XIxBMcXCv3
50yCV6rSQzSGnnu7Ze3G3tlFpAj2lSldBOU3mZ7ivWL3rNzVEgBABXlchGm2+OTj8ebhApPClptV
VcLaauP/lHiu7Jo3+OOb3oYl2XT07Ns5Ntq3R1eZqXV/TMvgI+aOfdZUAVsheQfOuXNqCkuL4Gha
iM5Nt871qP0JtLjhE9RJ3X0dCH0p4FB0dku9T6Ff/JRCuSs8U6X8jT46n7YbMwkjd66LUPUrzWVI
/bOmG4Wz+c05UEnJdvGlzJsFssMQYqcKYlXoMp9lkWuXhuck4CiRQ1vyUXji54Z1M6KQl2QZacb5
6J1ugTsnilxLrwu2HWioaxWWGV8C5ztAdErkZInnlV90PBQDcXNsezFbvpm6v5znulW2E1qlTXSc
EWE9/Wsm6WoSqlj/yUODxAaFBqTivTliC/MEUKUrH+v6ZbP0c9lE0vekvtWKy4rexahxsU4vcj5R
5C/RPz1k/Z8DAg41WgMcMsD37tYITshlLdZWSUfK3FRfk1Wl5BJ+WgmYVIIxBd5kUGknmlMZ3Ivy
G3efj7e76QyhRoc2z0AhmURYqgeQ4aMINJtvvz9E3uuFcUhLNT1lfaop/hyF0fEnAi3DkDT3XUwj
uRgj6xkuEwG0MrFW4zTm3FJHYsW32gY8HyqGdi5VcGVBcv6Qlo5U6xEGJwebzVlW48C29vBhLXs/
RYMCQ3NWxCyEHUHipmmJQkSQ+X1yzHqri6FH18H2yn+kZfRWUeTP5XbpK72y5CgifaSk3G1raWqa
ygVWsoVkzVUcV7OtcnGfnnBqH1W9ntZQG1Omebu09OzZUwVzXLQ8TUImuyJnqqi3YH6gLKV2Y9tG
EhYY2ezM3lzGf/duqDdVbYxaDXldZ0e6COYByuJoy65AKElmBEmxUueCWy8/MfXjYJCFf6hWDIvl
cIPLhycb2vQaeNnqqKnbTniGBqkNcAY0qvFK4YPr42AlPaBgoABeTOylsd7dlBkO3OMT9J4fGqsg
Y8DqANV/El/mGI+DTMn4AcJ1KVEEKu4evzM0i6DqLJqsqeft7IUKGUn0667/YKWUYvWirp6bOa1G
GzTe8gbeI153DfVojciNig/6IfKskM6NJbs1xtahyjFeSfj7hfLq3NPFp3VBX3eWXpjnGoNKTmGW
8v/goZRiD5+6Oq/+7qV3EsjoGZYMPshWmxRjO/AMGEzTk4iLEKeYpFwxglLHED9yWv9OP6ewu9Eq
1KsGbY6EN8Ef+VO3FJk9MoCoCfPqXrvx0OxcvFGUqB2cbGOJAMbSutqwE+rPBDWhF0D37ymcO6Fq
g61dl7lGhZJNF1RhFZjy6Yk5nt6kjk7m9o+BVh0GoFXZ+dXqk5a/Pld5LRDE4fs7wkmqBSFEom3X
kWI68wBlnuXuLktfbT6H6oJZYsmScpUyR6wKkmqxr/lFVHsU3Al0B4kTUc7c+FB0qJ2V4X2kOTsG
eaAcXUoHbMgVTMr8AgwrZ+/tE81NZzM/HxjjF0LHlEwi1r6W+bdD4Ka0BoK3un8XrsUOQpxMByxS
aOpGwvdAEWyI++tMQskXXsIKnKi4ZAUiyCczDwhSp8joFXdR9nQ5HwJ4WkeaFCu0PLSdUGBy57JR
OyIJ0MhHUOQ1CN+5zTUTt8kpnUBVNBF6AWSkVnYHpIZMyID6MUqVd/C6C2N1At/E9QsfWheJVnyo
OAEJghZ5ZBrInchiR2b3IWlII2zz22eiu/uxL5F4sfIKXxt7hymKpLxs4llq/GEJZMoqD9de+0Vc
oZMePPv+ELKQXN+EDTiN4ODOQQakbtVfzvU9+awkbYqWrgAWmcGnfCZ/3nesid5HtaIoY6N9Az2D
luCNMA1F/iYKrunk9uwvD7+lHml3PNBK4KOLcgxYNl/GS7bZMW8w8EvvQ8bYjmFMsTCZj3YAH5B3
bzGNMLOTPqbqg3ZG+TG9qPdm+AZ+v84zZ+or4FiwpS7fNL7LCB9wWxTx8YBsboaa01u/LO+go93b
emlyfX6Ec4nDynkw2B64bQvScHry2rvO67MkO7vSPJVZlagupwP2g8WXJ2WdACQuvxOnlTkE/wig
trVhyEaM9rcM4VtWq+LvjGcgWx4FbeErffy6rLUEeH9DaG6/15VMcCiP4KyhpaBVfhRWb9FAY0gu
AP1pkifiedDjGo4solO3MMZZiCYSx9m+PZ3B/ImeZ9lyeSvcAAnjvZwqnsB87CJ6JtocQzL6F/5F
YdGaKTH25wHfjYFvJly1ZtzmB1eh1Qsgcfj1jhh1kJyEnhwcin8EVNrBV4vkKOFs+gLogjpf+RD7
UIJzgkWieJ4ebKelsfqvd3TiRFxd7vch4FWpo5JTHARgV1zmbDY74lsuapaV3f1xEZ8y5RcM79ta
2SBebJNqzFsgJ12V52NylVAwXDrYmgosUSQkpVjTiEKJM95QaXPAXI8HI0rGZJEhasNvd2A080Fa
EKvSkV2xINOIhX70h0BHbIm0jDMTYuI8hrxjVz5787Fxkpy05hBUN4JkuKcXhbqJIeK1da3Q28iS
+sNbalQuCatay36GktL9lBh2+M6KrVDZeiFTpVN0SGQ8E9704/6ZarOqPl4JHK6HEjTAbPJpGTIe
ktQtpDbWqR2/OXNagE0DAU33uLAeQNn2NZGMBXt+yXiTcFs3MUCSK6JdIIIB51/BKHQqhM94xSme
ilIvv3z07B1HnzHRARn2keqfJy+ngAkRlg6cD+YS1g1AVlCOiNW3p0jG2auPIw8OEZaA94/M2X1r
p10s2WTLK+aeKM8JoHpXJT8/AOByc19gxNuglnCLPZEudebBiNXlvlps7A9sz7ihk/0N9zNQmth+
RXvs8uMZmtzM/iQpSwBINVn8E8OoceLxlt4YRko9fl6yDVgFhd3M2MHQ1M4SXqsoalfswXRmkKEK
hjnPu3u9etjZLnNpblQTA8GSKWxISE+wf9MXSmL40SGBVhXZDvWb5G1sy/LhtjLHbpMuHuUok633
D/+GphLKGzMynG6TSpvMCebHE1Mybhy1sKRx6bteYh7aa9RXmDqJgWcuWiv58iAZb7e9C0pElz9b
FyfaH54nM+Lg7lTKlNO2EnvQxvrgV7IScGFt6FTTVvGOW0EW1oBUSeroY2nRtrfuE9FRlU5HIguW
C6b+MTS3IQe8XwmZdBhWuAAnsL4yfd6kcoG2AW2MWXMC5F4a/RPCPGMwAYPrOR6affgbqAk7Ysvd
x/Ua/tKNSXmf7O/clJWgh7iaxu1fMOygz8Np0vRI9JWlZ/yErTzxFY6PKhmyNNnql6Ncd93gGSE8
5CsWeufLBrm5dEdokX0IHTQzzYAvvEdEn5UtMuiR7//fh9fUUIpIrnzKwHRYZdxjwUOq4kJ2Nf2V
lJlpW4wP4fmIGUEjx7xrSyrOJCHb5GGy0G93MNUtc1k6mS7wmKG/iLSBbGL5don7kheBM72MMjhV
SZ7coF4zGAd63wdL7GYGqG4jNog1LMJSt/MxYmyx5EkxCC+nvh4/kg1sFiZLzmzEaqBrX4uQJGTH
kXqVKDf/KnjRZH2cKpYgERvMJVjoJTYqbaXJDdg8Fe4XLTamvt841IFj7x8jNdRyHfrvQnTBAyQS
T/kMRlVvFWaHjHurFviJ8LxcQ/hKtsgkIEGNgwskMZW6znOfpeAsM020KL4w+AXRgUIj2jaiWYby
pIJiwnbLi4EfCSIwZgS/u7Z1v24Ps1IHOalVBAplbDL35qbmiT/rA0sDnrVAIRx889a725xiIkP6
Wy4kJ6kBB8OQyCdJNIbyAvx4D0o7b+zWqkW01vFZarwD7UaX2L92VMXiF38nEWAetwz6VUFMauQz
w1QVWj6CIuKHjbEeN9oNQoeoK1mep4b61DJBUvfe6Tgl/4D2M+h8pjLfcMyTUZkag6blwPJlcbsr
tXIstr+kCYJ+9OwEhWp0FZryPLEMa3tQ+pENflFJ/qqAoaEy5noCWnt67ypDlGdqMSFWG35L8n6J
jbOKftqX0Vq6/Qeen0AJj/bWNtuPHRNOU2E24s//OmYLKXg7SgaumujHO40H6B6DnTnd/ggCEbVO
6Fz2v4V/UK+EoiIIGHqsGYFyau6aqh+A5uJMS7zsNF9E+cq8dW31CezLPIafGhoriAoklq+z84WP
AQXLojTx76rMLzAYkDZRF3u1UsOx1+xjgwYwlm8SY4kSdot6hsY/NyR/cE28b+STBaDXbZc80rbH
mAovKomRkh0WvuUGnNRd17pIAIRLMuhnJscUwaaJzJwwJmd72lpEOHgx5vZmM7TZIDQLzXuWIRav
iYf0XlKbYSKuVfu2pNLJNfBniVI+WpNtq2DygcZfTyLBxrnMemE93Sd/oXR4fhB89eWSFO/HmsTW
P40v5vECtzKhulmiJ6a3K2Wr58Grn/JtmNA1N7QW52Am+ZVHzVAZawOePeaT9ZGo4GQO3EMI5T3I
H0UKDM3HQil8wyXbzIm1Fq2V/kcNHnrm63FgTjR/xsbfBQGHIB7UpUeZb8rH0Cj02FzQSTSJrb82
r+DYzAyFgC/eT9uHZDiSDFEUtXHaTOPeEqCoOmRoqBc1yzF8Rs6HY0801/Ad9f8CjKvOC0M/uLwu
E9uPIPeN2I1ysPeJBi8H6oHAK6VKn+SZEaYBFYwg2OXw9+NNW/cYbn8jwJ0Ej8n2fnAkvdZitPgw
DXvT9fCteJT6cGPc2+5X19U68vXMtzXHs3nHAk4yniimXSgNamgNYUSW6P9Sun2W+1m7OnvcP5yL
hpXSZ4F2k6czx9i9/Bsa0b7LoL6fRds4qGoXcz61o3j6kEteH7VD/L1kIJxkTgimMaxM3Id25c2Y
y07Skwj79qmySIWg0dw1ZFFVcLXR7Y77dsbVO8AikPsNHH7rzfuSKrYSd9od4HGIoA+XvEfHDPih
0C1Ub3senDIFOlDygOaxTg6bMCPrCzzYwwsxjGJYTFAc6YGOD3oYk6edrw4lndK8xcLgjheQPuiJ
9ydyscp2GJFAMlkIMyuS0eVojvUEpemfgADQSF1F5jk6Rnp8Uk+XvOVWdbxy7ZSW3fZFbuF/mR20
Hs0HzJw9ceYtJwlNple8v4E5xZvf96OLe/LPQMjbdxwb/Cw7fZj2PXw2c8f3R3rbSAyAmp97KJHq
xmDYtr1lB6n6B5vmUl8XAo9iSKvGjFg8gNvZ90PITbA6vRzzc7ZrK8g8ElrRsS63a5U0Vi5S9WUR
Y3lRvMUDBeB+0fghVJXMvZ6xHbLNMNlc6Tk3OvHxIZuf1ID7keyCDbx7arVZZ4ZgPAmZWcM4Rmcw
Ok5t/RxKTEfxhnmC0v0Bcjt/xD3UxSOQGqhrCJFCo0XevfZSrn6pTx+WF0R+NYorOxA4w+yI9ah/
E/2S+UHA++hIr6/adHNxUxDAAJetc4BxVZ5te9plVYN8VjC5iX59VULsIKCVb5wSZyXr7/va1W6p
Nan+3FXwfzQbDCDAH23NveKXF/UTcguYzI8vJ/VkVJazF2MEtk0QWCR0WB8uDphxHotQr6lQefGT
wNSkGGFB5NMYcWvSJA5VcS6ExZSbfThG+JDRKQ0q8OPP3jmeEaXtCVcVQ4VmYGTi1EmP/NyTyJAk
yeWSo+h5cBAj/+dYhKGN3yqHe2fl7OUTdL7iqiMQ1KwOsVTMCHwfGqEi/UO7utK0CdpZZ/Sge/kS
l6IrzKg8EbBfewJ9zuDh1dItF5WdfYeucfLsFPjWJo0nbBiA+TV2A9ZkQ5827CPxR2qTpt7hnFey
qcHY2MgLZAMPDBOQEs/lLBHvoPW8Ugisn6r8VGzwpyG22Hu0jo6NcsK70LWT6tKogAfQHk0i6YlK
xozxix8hhc5UpHlAAP9rXU50Eiixo3tPHZk/tIL3ahO8P65HK54Vev1/vMW6rYWkHdOlYc8fiSRD
vR9L3sOzlQm3k8d4i45J4mWpH17Pg23s+Jq+2ugIcMdT40eHlfBvEYi9pQNge51zvjkL2nAh4QNz
2Xs1tPao4Q1HQ4QaT1oqqkKTWz/ooczB0gOSb0Ct4EEG/zSosIpMENJnCuKI+gqtloFwmdurpZlg
7pGSlgM10Zap6DFg8dOLAzgdlG31hhLsBHLvJhmUVESoVGTxYyDYKeZ5HlCkCYUz7vrmrPPkkn91
SXdfEFK+yFyG6QwkZKqNPiMVtoCazxP1us8+G/dCj9VGrsgXsfNGi0d3AwAoLAJXp18e2k9MlT74
Ea0Yj2b5bD7KCveJC0GTpbJ032QLc3QBaPrkZ7fkloyjjzkit8vJMchnaBZZ/lZC/bYiBKMHvB9P
PD8j0z+KeWGYU45vxxJBVgpCjGh43wNmxi1cLU9l0+8SPnUQUuBi3hnn8199XQMDk1P2LI8pkssO
or+lM/2u0kEzXkbzAV4Bd4AyaUl2FKplSGDXeLswuG5EIplUGxDqwoZQSb4HPJQtKF1MTLFYYAqh
7N6aNz37vEgXfGm0mE1LQMcV6xMyHkJNr4//Gk9gt3pg7RdOfSL7AwK9TEmvdsUuSBMtDwHLCJE/
aAsR8Wa1/XQXut86q9II4dPjoRqsurl35rLFMUMO5lDus85icr1Hkq9DlWUchfEBCn2yRB6z/EYW
re3fkbVXhDIy3xzN0v2G3HNhwNH3YtIlclkaDPEiQYLiRmnou60lrgg5H0u2cpgvSWYLj9W0hXqk
SzAC7y5IziweX/zJpN6bCMN4ibesP3gaspdzYMPwTvEJHq70PYSE8BIsfTmhyD/uy4KZEGbHfLej
0JT3SHQdW8P56kcTCjH9KmJUJfWh8OkW7JfKJ0rmhqRtgwZqkCq5uOeXbWXtvZ5xTZCxvpBBybnt
O2wqGWLMLC7th9uY467v3/gQeW883xlySXfHDVKW5CvSteGURSIc9vz23OEJCT3TBRGHVkBEKQUj
qw5shpOwEVXpjK5gglJitLBfgZNAoh/Gl3cpJSeSrzSs8ESZo5ZFHuHEaC030Y27AQCF6LGxRd5K
qDFQQOkSquHalNqrGSKMVu/hVKxWkPMeFNG5HkPw7LrB02Mdlo/KwKodc++C8YsYWr9asUrJuL+9
xzDqXQRTFNtRGz8sQdkg9MVpHljhhjAWNyM7zsyy/cwNanu1x7uGX1KE77lYDUUxBE/YSKCX3na+
UbmaOZghDhFxnxJfQP8yL/TVeLhhuHw6sVEE53wH/baQ2uORkre7rSu7fa0WaBIj1Xbd7c12nwUc
8WYttq7k/kh7S6XaoGo0cSw4nf7AXXvZY2mNCgydmCAqDvO+N/spCc269NK1bg1Z+/srtWhYMtfK
VvbOqBEHU5ZDrZa/yscWxGhNumvFYm35HDCbPyrW+BHBH3+Xljaday1IwpuGMZ4i5b8bCLgmKIKg
rjFAVHlwWOZ3nRt2sLFFacep6r0R4ZQOHgD0TfXB1ZlCRJ2fvps0NHpP7LSVRHNEhKAz4SKaMwnI
9uFJblqAiG1GDcM0jRiOyxtf2bJ/P4/6QqvE8rbGms8YxvMmTQy0uf1mg6swg1PB5do4DXn3GWui
2iqVFcu11qfZW7gPcdfFxdHCWt2JOf3t9PBwowkt64fOxzxcc06EXbsNJowUbxF7d2ppOwjwEd6x
QSndIPBQl7MYi0tG932gtb1LSvA8geucbw2hpXcJEWEfAaR3r2oaEphYizJ00mAOrNK+k6PLzFKY
qHu3FPDS4kfqmux9OTt31SRtIQHcN+1CwoIIk7EgFDEY51gWRyXSHCuJ58IRyW/87zFCUFaDAqE3
oZ6XcerHonyH+5ZWU1rJXDO65b9kb+2X6QJuID6MPom66pv3L7iiQeJ+uml0qomhf5Vy1fxzLt4f
p58fgRunRYT0gCwABpMfVfvFCxmYuOMgPakMmqi0fzOHmPhMJYU/Xd6xjo/8fseyLV3AlcYyLea0
PFkPupS4yjijJ1hYhEfiovmbLqSP+2DvTeHSxHylH1Gp9L9jXuGHjAqHsk6Af/d0u7NvMtXjvaab
I40A30ALuSAhXXpCTqXjq0ZcM9xgQX+oL08rwUTQO5bcubXcowUTTCjsykeyUqrXP6VMzzFSubqV
BGGjq+X0GxBNrAMS9GTNDkeXKPgnHgX8WkanBrM9VzUCKaXbT3ZPM+8jErOPMNH/NSxC66+0gCGE
uzuzMjPw+has11dDQjJRCa8Iq13N0KolOSoq55mOgap0Rc4pau6Nzj8LBLeGCFDJrFfVelFhfsQe
DDypuPl1qVZCh8TSRejv7s7q6VNOJ3bnSqxjqN4fDbQ+ytKg+Lu/TkUhhduSp84lbmkGtJEwd6kG
YGuuSzpJjnnVNnHr2YSkx6HAZS5MdpUXtzDf//A4aQvrBPKp3Kb0372miVFKRBoLWQFaOqY0zHsK
hVikPpn3/u0guDHRJzOPibGzj5Ex7ThsU6725X1HZxGi/lcmx8QnqZU0q5CU1DIf8s4zOhP9BzFV
drQkKGwN/dPN2bLF76w2Cw2or/subyoI8y/89muhMkc8904Wqn65zQs/KuP2N1xbvECBlt+NHMsr
S1tVqFFdd6L+B4sfxXwkB8cahu5iHS0xoRJhtEYthFdc6G0DXWlvAP/m7CG//flQGkrKDnbC3BTB
0P21JcUoi0twYfnbbyEPWMPIKKxGIFQ0fIbdz5wOgrjY/KzzwkNqeSzEji0kgIqogc6fjz1sZO3f
7/K4YKo624bZdRePsE1pNWDTsHcbbJuXPhjdFg4oR7irThoX5CRbebXT93l1rbk0SfIS0cSMiVB1
fpzLiFTJXWGlus9PhvQrUaglKhX/r9qmx1JC+SS3yVHTnjUerWz6KXzlCoJFT2FRFk/3unlDrBQl
sfQnEy681aIYURtWbhL+Nz8NHSBl2OZSjLzC1kjWstB9p1+qrWzyxzbwfRlnqwypl9gXBkEHmHKU
ktnWx4cLXytfs37CFPKob5qKG97TnimfTY8SqpGJDQI+KNRcE0ZuCy7MrhbDlgOJFYGl0NP8xuSv
Rs/+KSzmY2+dc9+kEernA4jW1NDRS8z3jInkWVdsccn9eceuWc6ED27ujwvkmk3zK4DZ8WStYhw6
NuMZfbIjaOOUezM6o/3vFHw4H7pf6Gvy935w7RGyS1Fqx7UVAD5mALb2jVpOwQo6F01QIUet1v74
amheh5FWux4OBYao+AvyeSqaS4ZcG+/+2AUdjqbzzs8l6M+wAiXfq9SODk3c1uZ+7gk/n709wn7q
UgQHx49mqurudvs0XrDzhFcj+F0rGQYNGxFQeacWWCW3Mkpczsht3ns/xJKrAK2MX9YDHKe/nNMR
Slayj9Bq+zngA7OxFZq8aqi98aX7AHCdFG0rYH0OUfrtfs90pdsZ55kPjf5FwyUI6eAVdKiPfSVL
mnWC7Tf1iDDIt/ZwkKjTwM3Z2/3itLlEB3oQlu/OmOPDX73TXzeAkwGHNrgcYGU0FliM5+9kwtiV
/OeR9W/bLo8so2olIyqQho42Tp+MPdGyXHCapkH0LKwghnvYGvNmkSP47DVEurmItG0Damo25NFM
uT+f7Qf72SlnYjNElO/pfmmo+tQVgN5I9til4ZbCmILlYX8B6Z8F+ZfGo17eqTQMtw7vkWaOxSS0
wVlDzBGXiUYPntP5k1rlNugI38iETkMfL5/V90cvkqwyHSOWq/Px4cVetTmviZgfLM8B/TGht8pN
ubeDqrBb9GjJz6iHTa7DNsRDkLK91/NFLugekSfLs1tentwgmEJGAgBVr1sNhKfIPgW+H3YCT4kB
ISEpbn56wqEQWKs9U51bufiY1x06Lqr9w+QYUW98QA4sPGPnRTV/XMkyk6cCW35g40roXV2PhBDm
wKHeZ7ucvS/cc4TTA/rhArDrDjxg57lI05Y31aXw1ZI1lyhr3xcVv+RH0HLKYE82u4s3t/80vP3Z
HjfnIOgupjnehPapLMsPv2KchiAHSNhQL8QsZtMGeTnSQ72coleDuuy+qzpXNGq0LkBLQV7pPhXK
e7LXxoTLxsjsXaIkpNIuK2dEm7uWrZiEvgVL4jMQ1ZdUdLD2XaoLOUsSwEAkPglbMUXRlX6gkNn4
ZoVZLA9CA2rgmI+9UeHcfHkhYvGex87t4kmH1bGcmz8UebU4GF0zGmFISxyL/1FMv0soUAlFDjTn
hJ6cWp4YyIADCLN7oWqJPJ3oC+mlfmnZEuVEZr5fGziLy5L23V0OtSlKD4KEm+PMjDTM4Gk51SYg
FZpruRyJbew6xP+01C0VgxZS0bELTEzVcvMkqZnGHM40Evq0VuLQvpHM0Ia+jTBpLdAQtg/zsPCx
TTWPyIFtpWG9G0tuoCFYMKarsBGbyNyV5wnENMEDQsXR1CDMw/Uxs6DkkvQiQRD2Mn9BujMChQRT
1DynGR9eqQCCL8WMkYvzzQM6XB2TnlA2ov+TCWQ0M8l3oi2PpwbzrxrmTf+gvbvTnCBOmZezYuC/
r5zG2M9E5hD1Z+rhAw5LwMw9EpTmkgjEkz/ZT/Nc4TIYqiq+YSxX9todv2/NcckNVBZCBo3+XS6o
Cyu4FCRa+z+2WFs7ghTuHbfG7fPz6X15FKIm3uwuc9IVEobgSKSg3t99BFiac9wPBG87n520Z3Gr
KxRPdiYO2PgL6JsvBpA5H9vhjB6nKys+FELpBbm9JTTSG4nDxGQ/LjUz1M2dlpkVrGAIrc2MDlK4
Y9b/fV2+/Pp1dwiGgeOT2t8zVkVmmsMywg0Czk04ESV7sHwual361hY4Fb0ufpaVLios3/EGVyx7
jw9odfAbgw3EUwu98MdDQ+eJdCl3ely9W49sWjdQCtKV+TLzfFEsRsKLYeOZGuMVEQepdsCaYXaO
A2aSRU/oYV555+jka6x8t6auFJASq+XTI4ZC3Hiqlso0H7mwB5ICZrVX8GXKc7u2aWxUPLANGL1N
DxyYCXqGsLoVl3aPrnegBQ74vfrcvEbb02C7kltvogsOVgmlMATvPnqaTQIu9VooS2ryrjPFQAhd
A1gzP9Bt/6pLjWC9wy04843oBfOQRJk9a7jTor2T236R2BaGvyDFNYpAcltfKAiqjasiEZWjokay
quyeXB9czU6iDhrziCZDDSrXnI5Y65+JlbDf47YTwX/cV4SnH96wQzCX0leWMbRpmFB1vlH08Gc3
yBdaOJ+icn5EuVn2a+Jn0+rvYgtflo9yfJPZ902nBI2wXNUg1YCX/EiGOEoKNtdqyGZuWUeiTnxI
zejhplftIGtorCWLpM+q0/0ILkf+xsjTe0HyT2wasI6kT3V284MmluwYkcM7YD5cerNpD5F9Gh26
4ljZMDmZhFLDqT8He73Vf99AQG8l//dmbpCpgnSKLVy789iYkLuQraoT3xuDj+rgoM2IIFzjKRSq
TrVsSgvZJ6OpZxZ1c454tAur7iwuswssafH0+bRSD0GPzQJJozfwHG+adNJos5AuE0PVLJnxw3wZ
CYVOFjIpEzhpCgESDr05MXYP+3g+yX0YRnSIOlrGK5pEoTYY0FD6sg8SRILF/ZDpyEsW1AwCW//f
HYqZivVSIUPUGgMm+kl1K2Gnm/zWnbZavCJPK5aq4AwA8tFMN4tR6D5ooNhyMeAHaC5Q1msZy0c3
0h04vT9xRFzH7HAIuFZKbeqQdVHK/ZLXlZ6QcY+KdyK2Erhye0q+h29rjtc0Y0QSv6FqVFcbPBOt
sP6jQPg3M0b5a4HydKQTxVE53EzRMUXlQs2V6aFqNk8uKX35ZuoKdCl8jLR4EXn4DhnJaj3tkhYV
RQtBDWlq9gTXvI75/FkDh67y23x/icjuRTAmCUfHRePovcOV93moPHY2O3ml42EDLqSVCJv3DgOF
N+DTn8z6lV0fs8jEUfFDfutWFltq61cF6g5Elv/+yhSPlrihOu26Vi2ACHIm8bN0lqrWqc5jDCYM
oU1q2+07oSiP9kAQ65qUgdV4qv7ejHojUCFMqnaIMn5gWc5GHKt3hr/pyc4nePQIWtCPLZiwWkMN
uLyqsUGVvn4Nt3FR1fdVd6C9a9C/q78SHnDKiPmL578DaSvr0WPFN6C1KmRQVzCGzGCUdWCoxlpP
an3+MkapomQHCpq3WEkv9if69nq6TQGwJmNv462W5w22L/8vUYhb6DCkHBsTjTJN4J7vl2fXaF0W
0zAaALfN0M4BY1zL+3AXoKgMKzWkx/cpvSwQ0qup27STC7MelG6ijQjrsMa6CrWhSVescpUemjCE
nWXU7PU+dsVQLdrb3VGHlR3UPZvn/a7nK4cLBWuOGU7VwmebuvVMIJIKtW6OZGhh22PEiStQ+shl
1VnfWGOSSB0LwhyYEQOTtk5KG5nkanOIWCrUNdpgSqRUAq0sh7IsLAwsYjhGFCheLnBrBg+bse2J
E/Epf/SGf+Xwu0pWEG42HddTm7daD7rgEy8I8puFEo5BVqCUA5Wi1wwtV4/gCwrDhdXerxGT8PYR
z9YCpFeSF299+lebAd4BdoRfP1lpLU4rIBaJeDhJHM76ACcYVtbjDMOO44uj7KFf1vqBLLhVoa7I
qB28O5d0FI7DA+FxyhHFK/nzwd6jZMZkz1bQQ2Uy/qIcC5tbk1I8/qOWaTilHkQb84LuZZ8fAw1Y
bXx+Pwtf+hfNAo+Vup7+0vyRsk3iKWMHU8HXkV2wzSOgHQYSy/uet9uDhVMlx/xOz7I7BlrzZ2mx
M9Y6sL/83WBldatL+64LEo6RM5e6VaS2kaham9m3mEEK06Xo5cmi15fHt8Nf+eYDn3Isyl7aZGE0
yobiNHc/EFsU+Z0tlXdqRx8mUxl+gI9q5UnwE1wux2li7yM8Lsz43uUp03W9oK5nDjoUgjxRM0Fr
z5Mmu7PylUc4BQsVcW1xq49HkcwUswb6FNXNYF9daKnujij7fkzRgWxO2OqZMA/0qS179rlOnKVs
uIyIzJDxunHrgRA3aN6ec35+nlqJtWyvGjNPht2jEPeibPRI2KhiwKXWmOnNHi8yoEBvyIda9l0J
2b3HLB5iZxU2wnODyFu8qeFJn5Rxgyxr4tw7AVSOkhlvll8JcW+eGQogvPvGmrxqDxoEmILt4wj1
dQu3ObKYFD30iyD9qSYwe8YTNObMrLHSnBZCNtYx5+ipIRC6wObNLYrAzbDrRJ1lWPBuSlhIFglW
FQwJY5j8XoMkBMDQmcD4O6BjxtpDsX4XK+ITjFBE1CE3WwoCQKdtI2142UXXwqfFaQgARzMbi8IY
+cUd7ZIWrD99jIs0otVbYRRunn83qwY0LrK49WLnu1BBRJ9e5475lCverik84RFVSzoXxOYnKlPI
/74/4Z7lS2kx2/lTwcGDDNCkizdx3A8zCcx/I3u+lm/iAChXz1FTWQz6905ObaueYV9R/J76lOt2
3FwONY/ohyJpOMsnXSU9ywzWSEJdi9dnBqPpxtR0edqcNG61TWIUxx8wL8zZHnzFbcbdbEAHKzV5
j2J4613wC5/u/zjPc4fvJ1pQzw6rYZh4a6nmHoeBrSCSLAIgozxYnGbqkTJGHMjxHgGDU9fTyX9u
nFfVdWw7S2TmBVRPipqfXIOzHECadjjKaF2BPcUX1KfbV7I32VX7ZqdTxaLzAhaO6ScaM3PmFy3w
ylfsizhHcwowPYqtaAHR3NrzvPZAGjXRSBZqvwIUbYdzZVKoU5jR7wenyfmO+GTc08hCMW5Iy0kD
RUrZlrsURxvHKmKeAIfiFG6+U6HRhimg4C6DjZIM/asm++MCRLfg6Xg7B0NwObcDhnHE70cbsTY4
JBIR9s3ZXvDzCnj2Gjcd8Bn7gfjQTEWjqVYqbt8d/Elp/sEgpodRr8F+YWv/hJ/wrpDKZZxGKcKT
tJn+hLpwmMK/FhcLb+zEZMr0aRXmRI6g4m5V9fKSfuNcqLtX0qngvqceSDL0jAxBEIGEikfEGlkK
18rM3sooN1m27pgJKsOMvoCi5kogB9MUwX7B+7K1MjOZq94/bvNiaQ/F80D3g1FlhzmG74YUjDyn
eF3JLp+jiEBSVII5pVn1Lp163d4BteVnCTP2S0PIkMXI2QSO/Awws4N0EEmjwS05Q22I3w+Izag6
a5Jse3mWlEOryUU3DVBJbrjTQnBB8mlbfHm81G4JsIaZRprGIx9UeLKBWPjtkbHC2YchzJ7YlNsX
WESgcyFaI6M3+vCkskrQtogundGPlDIjI1FFH3z8BgGiT2y5WD4Vlj77634x2mRMYynEyWZgwWyk
GS2Tvbres7XEqv+1QrL3sTB8OZ7v5TWxObfFouPSHvgAS8lz/mnJSBqG5dH9dInPsBvuOKDBxH0Y
AFfx2EJLguCMFVBZNetb3dDLn+ZPe7n0c68/piOyxsnLb0Slg+8D/7AkRFzOfkuuZP03dorqDl0q
FgTHHjNTqbFTEnEg6DgndlYrfwJ0IYGQQYHBmtiDDMgIxR+MY0Myf5aRtoMNKpkmPPZzaPOOZ6aQ
v4bAGtawOKrdw/P8d4W9ttSMZp3M+mJkirQNpqtN6iLJqsAB+bh2XsbiZyRwcXQfF4E9xn4+b1kQ
V0J3qGrNGRCbNvLJ/xf1Cyp3ThSgaidlPb183qE+oOIAKkex6ybAXZ1e+7zSoTfftWvkSzl2VulQ
6n9UOi/wqtmepNyVjc0vvAEb7c26RM66L2OTo0BGfxx8PkF1mkVpliyhed/ws3Bucn/JkzyMH/77
oLouuQqkzlWh//15BV5xnShnnYCT+DgscwmB1k3VTMyeu/6bNl5BOdpZMRwkOvKd2Zv5dOdPQiWp
32msu899Hd2FunEi2A0GN6hRUeBIPr7QP7rLkiDb1MLMVv83nttuZREi4oGzRloQE+gdA433kME+
LjRsBdpJsEXJaJG9q9+JqycE0niAsOXPoYpfE8llhwVKPEzUlEg7Z5HCMeasHTtedFnN2jGoVfo7
hDLB91JaoIQC1CEvnSdv84G1IrHcE2vPwM9z5pgPfID2HLtNXAIG9qA5bAYmvR4jLBACYA6CdfIs
y018T0otfnBOZUExiIZ6CYi0oFTqGot9LiIX0GYE9VDTQRI3zLpe9EL2UWAPD9QpsrRhvqtOQqud
9mmQwRwM4c3qG12myRZTasv9vXh+BRHzpWRRjHdr4lK5ts/dM1g5hBgAvfU+2sEzEoq5TC4reNh+
4cllWsMqhgTEcrzfmYCuJnEsFnr45y6yMiiTaBQmF9auIgVZ7VhLLQ9qzeFW8sISfwX2h5TJ0yH3
5/Rwn93JsGhemkQTjd3wjcClc6DmUobbLK/vq7wtMEjPv8nvxOj+V2a5NHSfMoVY6AKC6yTwhssY
cRO0CgGLx1IFXFf3dpiwCqxlsRGCl1IBnxJMLMmfOPxX6z9frgkgpfcGeqkEIBuaf1LweRi3Mnb4
7TqyHTGuVN/iuwnsm2dqc+z+8R/ROqeTbHYPFfJWTj7S8QSj6/I4I8TfQ+190bXZlALYE0kmR/8y
Totj8pi3TABt8d06fwOP4nbsrxF3q3s329A+ScNbQ3Vp6yH/OJ+PZPDoOUNvxTiaMYsXyT7tYpGs
S7R1UVn9zTBFsNVEklmR74NfxZCVBehR72b8ZEqWYqF08BnL2ibpZuHSknrvS9qYYTDeK4dFdLxh
PU4nsCS1GMnJc/VVcAqK2eNzcDWuSIWEvi/txMALFuVfIIdy9/UdaLDTVrrJYSIdbiHpxIC8wbS1
5Sol+ZLb/wY09f7JrHbABQ7YV9cP+NJ/Q3PYiE4XgqxkgebZge4AWUpynx8noiQGJ5qa16QUyfD7
1sfNk9+f7ZCNBsmE0uyy8EHOdDD24ihSHO25uWGtM7FFtvwDeD7WhvKGMzmutbrlAWNBUpR7qsqu
wYI2nM/k1OlohSahYxjbWKMU7vG0WQDRC9EhQYzOaNnyMAMpKJRotqFp6supTjYgO1wUMjrgxNXA
yJqF/KJ3UnByvYtxbv6ZgrVU0ojK3PHaOyCoPiEqGg7JK0HY5nGDX9tfTBKys5NhAy5DhXkL6nnF
67zPbxOApPwJJP7VawQNNut4CjzpQQuaYFVTAKR7MAHEzOgKM2KzSHKQ0FPcv4jDMJUIM8HZjTY2
zkfyfenGjMJZuWDtMqDLB6H9VX1M7vEPcQmjJvQ2MxePegMNUWA6gbEUgrdJpD4Zx+6ZZY60BZqp
1VxC0A7wfdCmKmlaU6l7svosZSWs6xlIDve3jSMTMWaBfGaxsKYt/TuleKAzeoMHR+As2rMJr+Bp
Qd70aLkyF8qhXjNZS+VSPrriTU7KRDMroWq+AWEoy4j1Oe9HcmjqqdJaqd+LuX/EUsTBVLAPkRMu
2kKZ6VPpQfa/rhrd1e7njBb0DTEffmsA3nd+bqxOiyQksXRjPc5uWx2DshX/mb6TbaS6REUdvLTB
6MMuuSPChJWl2Gi0mscCu2ueZvYTUnlu6KruzKcYVj2x2OGARRTq/HrZl6EvCnAuG14S2G83NqnC
Wp42Uz1/3XZ1/iSDruJkUfBtXXRldOyF5/Xm8CRS3q+FoyZ+sc7AYUh02+OGijPLcC//hYWcsUk2
C3/K/E1HrECNeJqGgOAX9hNVdeiWm5bI6a2eShaIzHaisyeD5qdHKQwiA1swGNGVMz/hqhibSO/X
yBrz3R5sk5lztNiWJ/6T8BwsP0UzMpFrbHZcGbA3kxSWghbdyR/e7PYthnHM+8ZVZgww73cCT+PD
9/oyRmW5SwJ9n9gm4TmEJTzTuihPYPc+xH1dPQp3Wwgn/eZPHcoGj9/ZCYSowe7xixe5Z1rBONyg
C8lOmIgGWOfpPm+ecyeIMI3wqStF+1qOBmCg1VbrmCDbdRQnKXD2OPPuwLKTD26YucYO6WZCIlHC
nTiSH8wSKg81lyHKfOFGO/h7LgIWZi6Z8OLjkhKA4NpB7ryGggTpYHH4+no9PY66Hh6zrHkF1fS+
YC8pH0Ii4RpPK+zgMfYF2xiBN27DxDof3ZLULPFiZR+50w7PEQB7npXcqjqSdBLIkhwaZQrSLDKJ
AYQOpqpVRrCAwIlb/hDJB/Q3qXpZQ7TwUPsLOzdHsuXCMrM8j56oenPrvj0AWKIBfauLPd3j9pLE
sA0JajYjyldcUzfcLHFJw8mql5dpVU7a16iCcWmdUT7sxnw0/yfk+vUvUt23yn5Ovrr84Ohpd2NV
ePVJK/moRtkqSx0+dmO5hovSu0aTtzxmB6csnSvtSzTuXyzWFNopaAom5z9AD9OXe5rvTEjLUsH8
8ige9ltJuTCSf94pU72TWc9yGpZoKrsJQAIo1vP5EXDqCO64JUTTfDjCAsu9m7N1Wu7Fswd0ElOZ
CZ15GH951uUaRpqKK5ZzBNVlW6lb9BYNYpvLCnPAeskqYSN37p7oGdjszbwNWJogvPwKu7tqK2Xq
KYCNnySssb9SDDtv7XLdomjJ7LsI2AmJyfO7UHnXSXrmAUINFp8Wp3Su0C7cdojry3fTp6Y1jO5V
vGG0fPE58Bb1fMXSbdRAmff+Og6HMmn5dBYm3NVpck3uwKK2mLKxkGEFIuCLxyuSMF6gaYtPnnOI
SId5X1bQiTkRURFREDQMcO8JW1655gofUhIW+qpySbC6gP+dZGryDOgkLIrIMriagKnTKa+iP6Ax
qZHpoCF58VO4UqaDYE7ivUzVRzSOvPoeTeB3IoiIDvJ69oXPrtk5O8BIAxzPpTMOL84TR8t5/koN
CLy/UUzUJ3LPp4cw2xOQL6oElG1Iz3NPYiYC8A/xrk597A9ZVm6Wdcp2BvPoieVsjmpRk2NzaXM5
Im9g9XgyzotTyF4aa1V+7GG0GYPiXinwOaCTGrgYm7MENvWSpo13jWre0wENF5H7Nn0hCMYtRl0X
Cj7YfpwCupE0oKYTHgTYskNtcKg6CfJi0rKwyha0vSPXh6j3Kx2+gROrPO6hpnofl4cWt2NIXHEy
Rho5fScmWojonubUFsyHmYT+iTBF6MoRpKK/eSgQSVQ4WCLArYcxVp0v83fgdAXZtvLZbJMzhP0I
AEPuTQscjlmNa5qm+7ldUoaYH0yC+ujrcdi6Iw/42MX/naa1+PL59aEtz8WYkBIgomsZr6J/irpx
DMeNSk4rlHHswpGF/1yMrl9nPpft1F7UkhJ49en/cNiQEVHDC6UXJ5miSVKNZSNVyyFFa4AhUq9s
nGeo6G5PJQbtCc9yu9DmUMPMeJh399lwmtIVqHS6V4q9GwkHnFPKVPfmP4Ipzp5s2q52YGGzowfg
AOh1hJJDo27JcsLjWZeJwlpcu9EnpdVSis11hB8CQiH3nPnIoM6/1KT9PN4JLXioB6c5Lghu8yHD
xOXGudpkB2nrBW8p29qhQJuLgA41au68YRzL4bphR/OPj3sx21XzFCms4NrxK0zVWjhhMEJKMu2M
sJqS9Y8ONPTluJxj4XELoqv59xaNTjRk6SH8737sRU0J1Ahq3mCi/sYpEk2efzisketFl37+QUoN
DkMHcrLOIAdRsLhkalJiX0x7+qRMQlXHdNBEsEYORmaw3b8OZryIqHhkfCJnOEjQRxl4C990S4/H
6qVKBS5Up2wZiO++72sjzHjfZEIy5S6cjHs4B9Pc43OgHnozQ9G+50IACG8J84+b0VH3HSHUivwx
TMuT60G2YPRu9mzKRymYL8c+HrhCA3v1I5Gh91xX6F2bPa8Ur0cB5E10IoBv1A+hZSD4nRnoQBSP
bOXRS5F9Wmy7xzTm24dJ//QE/YtY/NHlGQs0v5QHFBAMvBlwlwjgszl8RNJWPkWzZ2rx1WC/V5D0
E8jNZCt9In/N6hE25GJ+uvdaaFnAVO1VEN9xfDlKG8ZOQamIbaIJ9BskyVJasGeLKWOe0L2/yfNc
NqQKcINTV6gV8g1jkrlgRbDAHxorntAflkFiisZ/Neh7xu97P3eXiHmfZWBaU7GiQplhcrjLRV8C
KlOF+42/aK/UszWRlhFNQg0mf3TyXtjzdOuCFc9tt3QG97cQTac9Ym11ahKynaHz7otL7xauUyNw
4BA/blSNKf0WI3QrG70HVssNuIqhQCFDa05mammtVYv6i63zREEFkuggAsMLgn0pF1Cd8Y0V7iln
aPpiZedk7TrePWKRCbA+Ku71NKaDIlEssOk0Ymz2sH8wY5Hh79pwuYgmFY74dSXOiWFmsKmf0aHU
zCWgTD+13ZZ2UGfftURtlqaGQoIszLd8l6KDyIds41VqH1BtbllinGtkbS4cIaSBEGheRLLja96k
A6q/K891rIb4vKe5ZJFq01wFHk2VXmugq2Vu9sv2oovSsfeTudP2j9JOqoe6gGZ4pcIqPbhD2+Zf
DT1FGia8EhUNMeik8PaL6wk/i1rYmshP2g/uG5sQbv1hC+rDubENakUcFTK70f6pk5zdOBOGG4P6
oOCOXw/mnrF1TfhBC9ducpjX8PksMW+moFvZNo1V2H/rCLaXV7oNt7fNU2a7jd9JpW2LhHvkf+1u
LM792iFd/iD+nsPFuP2BIOBliHSkQTU+6b6+6bH1jzJX3fdIKUup28e/bmxgNrXp9mE4Yh5mcgND
jxvL3RsOP30iYWpZqlw+bCct64NZFVkLS/VcO8opEfyj+dllUg/d3IqpRmvLJuPDrjiVtZHC/69M
X8GpizezIBZdHPlW1A5W0Gzu8lf7NDOysTK38NNwHa4Z8YZGiqs0wzdRWAJhceNYh0kHqcm6blUK
WWvTIQTCtsWK5oF3Dk+H+SekbQA/nyjmIR4GPB6FS2CST4gioJHfnFddqevStEd0YEz2jyezUHR4
9lZBH6D+tMjhaN665ejLgzaEmbAn7Zb7zB/ezgZlC7X3ZlexiXCSKZfpLB9yLGqJrIma02jOV+pR
ZzbjpQe0JKIKKbR3ELkq8y3G2T6Elc+d+RmSsqjjw5dA8OaUN75B9HFN81LitR6oqLp1exLdygaS
16XkrfeoOliDHEhJEQmy434+QDI3NCkMAMIMWF8atbZx4M/qTpUwQ3NyiZs6xDt59gAgIBPnDF+u
veOyxJMd5fazkP+FSBHJEEaoQxJJso5kEarYmxGtGhkDXlpqDKgB4eie1jH9kkvesGv69W55NH0J
Qd6fQ/sZDuYer1XLTZSvkgLRX1p/rBknlVFN/I9lnFI2WVI/ZXuQvnG9uUBzhNQdhXTUwmRtHy3u
NSWLrgFMG7Az4QV4jUX9H2hbA12mf48Vj0Bdu6qMAGfsruZZQgIicTB/2DNubNiUh02xSNPiBYYE
eCAaX65RI6pDiFEr1DS5/JD0Zpryg9RTtrgCrUlqKxkLjECclEIrsIDGDxYIGKX0nPS0F+ApDkw/
iIOJHHPo46CCz0uORVDUArJbNzmiTKE+ZtnPzZunihPnxet4q92C5GW5jagfPSj25y7tnhLosngz
sez3GFUkzZPG6+Q/NyKzWoboJ6Nl/J8oTaypifdtofmO6khtgR48IXjZ36g0I3wHlg0KmelskUt+
rCArG1LGZ8FJYVM0WtQ2S5GXx5eoVe+OKg4afrnXiC13/4QarGhKW+YasOejTLPn0kBVUF4Uhabl
tAqDck1NFRz0nOhl/9phpiMU3eS0jZZmEEYhvC/AFJ3QdPPZ8pZgbC7VCXb9DBptKspgk2HYCh70
lBecJY2Cx2PBw68QCCmj+13stQnMj/FyrmdkSsTk1jF39KbKQvUKAKKquyEJubnEa7/MxCOHJRfK
YPUj3p+aFXH6atync+3kUVAVIvZAl54gCM66lMphe0UaIuJ3ggzzj3GiQ9CIHYGB7hTcz8CBrnwl
ljuMUbd1bP7zdsM8T+cFCmeA7Uk0kJ42S46+jkzzy1tiy8RnC7q1u3Hiar3liAUBs33CUtn/W/9/
+C+CywthybGdygQa9QLT/nEVBarJCkQnTapKoRQDcikvi7B/9pc5LKQCgvNWYjetqJCFTq48NREG
qvKenKP3VgoaQJWLC990aeK6TxcvTgrB/9xkgg5l25lNvyClstYAVPM60J9Rsk0EoesPcE9S1U8j
PmpQIcvl5BHTX5TFOJJT9IxSkSLCN3ix43BSifjU9Bv29U2P8dwwcr5WxtabVCRf2QE2Uz33aRZT
Xe0nE0+0WkfoDbpcIwtr6PUyCiCREZgNqrsHLG4qRwimNBp/Xr0yCFrRrpa5/rzlhSm+WrjZq+1R
GCop5R9ve45xgMCuMCFDoFB6UW2xL8gzq0i9nQCp8VvJLBly93i8osATGh10zQ1hfChkOl4cpKXG
diq9O0t4Ui2zpf7DvDo6c55+/QaIs7U/Mm57SfOdoezhGLd3RFus+kC0NrpogeiRdGpHcoeuOD1d
0JbD96CshwtjE3xL8wp+k3DAeQcGw4gOFSGF36BTyqZPHSvox5kPX//XyPlPLtXGZgDMBQPnwPoz
sTVO0V9yP2l3/CJiUXaHkcpd/ng7xzXASdOMNYkxE6cJyweQfv/Pyomn6DHuRpL21JNDUYjUTPez
yuobDjrjowdxYeVcvy6Uh5R6mp2ORO1zwR5FlZoiBDFb42WExrBpnjY2eX0ZB/hmVTUP7xT5umdm
GzZcDe7qBf9d0xpEaMeYhvEmqrpuZQ9ohFNwiVko3pK5iKwar3OhLOzDXrgX+F3lYzmr054ISuZR
xi3pfd6EjBoApxC72LTSUofvV4I1cOvouWphKDmmK9oTRHEMut6ck3uIAQf/RKD0eL2Lt+0665v9
ZFa5aHdw+N/voSKN652AjhoBgpRpT3ViusTd0BH7sV7ypTE2RX+ORCGXmCpdnmBFAHm7ZXfQC2VU
FfH9cq33e3sLOrWDQBvKRJi7Bu6SNy/cygJheR/DBNTsdifoSQIzM39o+qG8fBSXbGFMGlxWzN6X
mdoeFYRb1OrHynWBj7Qg1VF3ACmBkeiix8sDsnvsynrInZLcqKeWDQQgSrcgu+7JNoEzLHhOSaXf
mxmWZKdIBNjNfT5wroiwhlYnpQzpH+EbwrbqFwi49pQP4kd/DvHj0q4veY5JQtHxKe9RrBCSYYkT
p8ugGaFeuYVhf8oqPDNAEAf0sGFZ9UZJuI9XFc6kp8VYt/eZA9TfkeX9S8e2m9f6LdsXryvfTUiy
XHMIlXqD3rDsHosEVf/cFv40lfH3AOeMZg6EtTbDiO4sWLwXcfJmOYev+Dz2e957UUcdXJifOIbU
4fGinu5Yg2stvxIacIcERK+FYkVJg2A1e6Ujg00YrGIVjHFAwmrdsz1DDDKeiYtgqDjc/1Mm0a+d
A1n95ZABYE8EfA3BO9tT9fFwrfezsp37Ao/kuSx7px1tUdo/gA8z43B63Mwmuo1A7CNy7GA9X1Go
o5sXSaYOlyYyvIdMxWIwz68x3VKyCSkM3B0s1TNYrqGR/mC7GcDBGpQfnnzE9efxn/06b8IbnqNO
4M6ZuXXmhe0UnW+k2eEfbONxJd03tWpiVPaxOCCo4veYDst36uiFmIjTamwmLzQ+Y/xr6xzaw2bw
jAUFqxgGY+SGuAPoYnkcS0dgxUJ0/vL8OL+jzHKJlC6EuMo2HighbEbvOufWoWhTqf0+0i1n2ua1
uXbAjA3Auf2r5w7EJltMO7N3+vjjY+RmBko7v0CfTohzVMSK5ZslJPy8OUFylCYjObG+ekxwmazW
O+oFuccGdVOceSXz7ViQk5NOf93u2GvNjXnuefpAVaOi4eP1ROXmRluyFF7RuOQvgEZ+gphydo1H
sGPGxcvSiEjmf2qmQwm5uG8mImndx0iW9qmpHwTdtYGHrl4Fpy44FjyNMC+yAx107W2fIMQPZJ3B
T50ULsy1+Ic50SdowU2o0AsTwW23S7vUL0s1/7h4rXgEqlvELkdlgBKvM4xxaWx1MJgdD2oAtbTa
KJzm0gUkGBsltt4x43vosCdASGHiSahM3Rp518cwjFFh0yLddSNzisZypxBC9aNkhyLomWy8uarI
kjA4iLaI6CwaoF9bQLzAPmoKPqFaxVQ0yggJDWj/nB38VIw8az4H6FLIMp7UpRnxk+CYsjeT0pf/
pXWCjTM2MA0g+yb9tk25PLq1NLTOVB0rPkgmjMbVLG46z+unok1XWtkOtqG6o77ILcniF7vGhGAy
AOlaG+fnrSxHo//KX98ycoFG3BjSQ7Hj3k/m2I+zQbw+O4EKmwKQucuYL7qRBksOYplxXX0ViDI0
i3/ALVH61MuL1VmWW/nt1IGWPPzAVGTvJ4ketGC77ZQzoRZ2rkKAJPryRJyM90Vxpkp4iM01qVlf
ZWXuiGzt0zJyJJvzD8OkRXxY/nqYaNOKSTiBOm8g72U4Cpk3pH7aFcqcXsp5HhkuWa5H31ibAk5z
hc3CK90ZXLAs7SfoZB57yt2v0aoFJXMogyy2zvYDZyKOzNBFRahSPfS2l6hbjGMEHQP8AZnhRqa0
GHnGAyTjUpMBQDStxuU90YZsq0uYmtVK4br6OBivr8X9ypxeVXQ2zCPgAGs6vKVFpK/mDQha4au+
8s9LmQoTTGSJw493smqIC55z10wSiXj5cCJ02umINQ0ZJJ8OFEEMz1kd90hjnpvg6Fng5s8flE19
mjm6OMl0m6x2K3pPp3C/tW0fXGziTJKCpy4hAGrZPHnyArOaH8LivSMr9J1SiuzlYfK8C2mmcbLK
sKEig6s4Eea4eqOo22EB7h7S6s0GFZivhjyZz3tTFbWEQbPVdO1lhaXhGXgDr3X/ilh+hTJjmtNe
f4Z3x2ci0IM67xZ8CsmeCYyle8hXLSS8FfW0uAd6fkzGDH4FiQF92ZvnNlBLOri0IdRTXycg4XXA
JUy9b8MjAQiiCHQ5QpyqO0j2AfULZNEuUYub1nTOXWbtLl3ClWNjQxtgrHqr2+YbwTXv5z3SXJHh
LRERcPWSan61qZvTT1vGOKMj1pJKEqIk5ZogYnPu8TaR8nybYk7toEU+pvZrAgUzw7pmMMCwDrhQ
wZM6h4so3BMbrqR4BTYVEBptOfR2xNg//HDYu27nU+u4BLCYTusvvgjScWLHWg1fgiv0OQh/Webw
anKb2toEGlMBg7V3IRY+FaOfHmxZx//9c1zj8cbZy9loqVZeqJAmDGELR01l+X6Zdtn9FVJJzyAG
BWxPxdO58Ip+52j/eBmDgYm/BKa3XsvPfgpWMsbGnaGNFSUEG4qfU2BcuEvG4ZX/RgFGoxoeK3Fp
uPQ8ndTFD+VY+sZu8qQm/HmPhVog1Yz0YkF0pSDc2DgW5zM0Tt8ORb0YaaxY0wJSNt6rrvqdSKwz
MHbPYpVG95U6PrN7AWZvjw7OGYc6tVjJR9oatdQiaJrn9kNjpFsXkzEWPS1x7EKL/DKWuvvyl5uZ
y5L1BdkmiB0IZo1/Xpdha1XCYnVDrVIVYjVm3ORoV/XsO35te+fDt127Ed88iIyDKZx/JnhNN258
GL72Hao5BnO6PE8iKyCe1v1ew8vpYUvOlVet2FaX9TvfmElBUxXgpo2LL1xCsZEGS7cQiyc9gqug
09oQLEFjpAp5eEqdq7JXef0Ka1CYMlbmjlxbEJWzWvVsQlCApKc0nBsqWgA9l38KXCLc8l3OYhSB
F7B6qkUYH7jkEREWyDK4MLO3gvrsQ4fqWvvIXlXLcq/hLMZULRN+MdnrUe2sYugRUQMvSBUzCw7B
cePoMzyLjjB2HLsvSHLvvCrZYjS//tvdbQvxyKOcp8obmZt20SuQ8XCpeK4QGWnmBKyizNFjPR/p
a2fF4N9/swArZKqoh9qVA2m/NAiM21ACsvqMahQ8vw+IHzIMDTQqyGLl1elYHmVU0tmw+kIW1CLm
RcuTNTOE7CZK0TTwwMflVtN0od/k7MaBbsJ5DuEErQtL91QIslWjpd/uq9BXKG4/sEFH+UYqM0q8
dKkdcNYvtnpSArOPFs96C+J6kE5apEAI7t4A9mzmxsZNQfdGfsydQNoR8D+JYoGaCOhGqkzIaK4N
8fNby7yrJPmn0TilGBZCQzt3w4y15Gl+pce2SjOTsN9K85BXkkcoCadglZ0AXQ5GHtiaRGEki65x
Mh7JEZQ9ulXUIL54AI1rMbmBYiNeSXh3h9nGs9f7J3w9ikENzZeEyNxeSfoXi5HWIP6McHH1aVYM
inO4+uFs4ZREP9+URAcrtuc1awumIOpAV3nbHA5FJohJGhcNjHeIq24Qh9dQbSVCf4GeeR34kBx7
o2YLxbpLWFyiAkReMuZr1I/30JK9JUcPYF4qUuWUOKTs2onUV/RGNfnjjLJqBxtYkLYNxK5Obqlb
GzLUOIU6KSt8mye0LI9f2UW5MynxnwWonSdVyrNwfw+Enqk/nmBuo/Dn/mkpWEsB1lBtejNpAiXa
nTr1gX1iNYJeQiaRQAD1Nlpot+clRBghateIUb/7CiiRQRTREP+xDRbmvH+xREsXFHt+P9HZwGmS
LVOBw22vX1mZyhpEnyVeJ8j6AFxLagCinNStRc9HlcWDowcvi6okruIRo9wDN/kExPt0voXp03aL
0yUtkft+dC1RqvE2pOGnSq+ns88JMdHmdgJ2ir8WRQ7PkBPCqVwiS9prOV2alX8h9CGYSh/JZyJd
E7uqvDm1oI0qj4Hz8aMCpDJBhvLpVHzCF2gHCZD4QVV6a2WkLdBL3df0PPyaE5e4lW1X318z0f1W
XvKgAv2vKPrLYC2HdXeym61itfZac69OLFX4412U25KEVjc6dUbToeOBAIsx1dMxFMUtqwRpTqZZ
cI+8kVNjbn32WOXECGpN9fdRO0MvyZe2KZ6qYcpy39PNqs1i+nuLdl0IVjUFZJJr2vd+oOP+gABq
4cXOkdMv1kcHJdpqchfuaYTnrwecC7zvwu6wyptKMXZCi942TwZ/o1TccrnYVBN6PUnyns3DJUtC
4eUdz4cw+Ww3ROdQKqXhKTFt5KNUgLWDS4tBVL4BeA9La+qaoUA2N18RLZQhu4mOog+wXGcpDomn
RHHXf0gHSn11HRYgUR/2jG3VIlMeA6RpAapwbm8qBfcYjSIjqCs3GuIZTyGzxZhtJeYwBUop6je8
hpZQ30uWX6ixWNHyhFn76r6G0HPfYMrhDKve0hwb1czbt1aqzGOhwSapfz6de/6GLRWd3gtgXJ08
UZwxUI2sDGt8uUmE0DYGxCd6bsGoz4dEO6+3PyfNsRyfljpjcnnb4oWRzM1Uk9FmoGmCRUggolzs
aOWCMAwh2ochrcoepmY9sgBS+rmWd1nRnMnSY4B5ExSgKVxQy83Zo0djt4nsKVqb3gNQetwvtqAV
OyAjvvMxXjM13lAf5yt9u/BMcVOizY8vwBxQdE5G8keUsXn8/DGhXHULbVgkb/YTAwUVe9GzAxw8
vRprtqFNhhIf1+r7tjLuAqQ+EG190oHOw7DfS4j8TVvVN6XWMWBIORm63Vq3g5gaVkVRIPuMdWUw
gXI2Mrt1Jk48ZB96TtYMmLVAXX4XpBu8dG2uD5MoU2gUB/zJOblcFP1UWiWe2QDvVjxbC6QGIFKN
yxFA63ohmaJI1BI90rPVRYPp4llSQgsLfvhLLlwFo07QykTEwbVXuE2uYoLr5TJwZFaDjRLPJ6pa
Q+lMnSv1EdfvSKJqvjplGAZtXVKnGPSy5C8eV9aSF7d8DYtt/6IqDO3mDsjoaSflP851eSqnPwVl
F9b0p8/+0NaKvmPamTlNvpfcUb0aUZe/PcHDqxFTqDe0KT+PhTf7YvEAdUsDjFjHoIHD3QLu8Fvh
A6UoaBLy7dct/IxuRRjPlN1y2YyPuDJ4wgnrX5xnM/3nbb2igMzKvfCVMbVomelPS0PeKC56uSQ/
e+YdI2Gr91PqMTHz1QmUHpSdvFxcTxXAw2gANfj6tYqpIVgvnuYWfgjnEGdiHlDtP9ueb8u+pgKF
4MuehG5cM3bS5ya8O+y6j/FJ1EZ1PlRN720eLiSx5LpINIR+9dtX7VqsIxs1/noE+TRCLiRzcjsX
6YEUtOcsh9eTV8V8jdB4zRNGsEZaHcxTP03vK2gIZpAVk9WQlgYiiFg+aimAQhGkhOTZ7yi0h1ab
zWJkaUPWIwMPqtZIyvtmyHQlVZK6isLEcI1+YGyohJ3rDww5zzOujoqFirfY0PjrYaK3256udBAb
Goku/u4pyofPPEK1ZaZs8yU5WJwLdbhNCN2TuIwurzIW+MC7gaLpnjXTgQyzAXjjKTHPgOMKOrJx
3lhOQ/0P8CNmwbPbfhwGPfFTwL19ehPnHVIDMZzF8hDqEpXngH0WC1GlmyrAH5Gh5wOJY7RGRMI2
kRWs3GWnKQFAw0dLNGeLoZ0ck1QLjQaHbBRY8Og5jYPgSBb59lCauzwgGXNUi4su2zSXiTIuEIl0
1IVLF/sMErmzkGaqIkwFIt3/1A08mePQt7UEnN9S77gzfYYSDw3Du2ACw5xzcKT0+3BPIJN0eeqL
nxkhyRM2j5iNCNctf22e3GS+1fALBPe47sNF773Y6yZNq0v6JRkpHw4DR9/je5KpxckaHAQ+Ym6w
S1zakbakMEVQviWWT4+o3Ukish06js017c+4sGOSS+mItcWIisjOUUPNxvx4O4DHzijnYGlW2mdV
Wgx0lnTDqcPdbg8HbXtEbMtblN/Y39kWgtEd0Ne6YEUO8uvqkSGAUCC8LthQ8HN9BvGtb07dxykh
pRrxW4jVTqk+FiimK9hEFXcl/+UMRfYxzHj+OtAsj6cE5QVVITQ2YZNi4E7WRRQmWkzDzoUu5cR/
NEHwqPcT+i2L9Eik+g+OAgt7KtCVvLqQQD/S9RgdsRRwGa5H3IMXnSlK66HZKXuIAFtSACPtJAmJ
ERlI6c3iCg070xtrmdmIZbTubMdYZ+CAAumhDL3ku+6/6YGNpzDhnEcWI/o4+ADb6UPLSJCUk8wu
nOLmqcKw1CY6JD/THaccIpJypj6pY/HwQTskCqfu1yAQYNUI4BL5046kUdnLpsaMcC9iFCLUs1aN
htCdcEBrjl3rlK2RRDDIFagMeVYznO8OSOHu4wC+cz8HIreZ2dmW3vqqqHY0mNFZxk/d7GrLuxS0
zAv0D1dCSLsrEBCd6falNHBx/L2R9xuLm4HCudgszmpUWCST0eg1ti6mjb7hZGZquQVihe52HBvT
v/HPDeqpa/hJSHrJ/CVjR2sbtZJGBcPvaY0mLhp+tEKv9h4hwlYEBAvcYR3iW2N+UqOueZcZXAUj
Frlum+dUU4SzThuVy6hekE45DFp3pUmjbjiDrm9FasKRdphDmrFP3Wa5/YR+WnR4zbiVDABdAmxf
/lLOfOGUPrIzzRhBwFEjvB3ET6dAH5VLB87XV18dOj3dC7AiSEoI1UhTjnRNodxJKNNLPJA4NMsZ
avtLxfO/JbInEbUEyib9M5r385iEuMvepTikEi2ii0oerR1UCY2+I8/bAsru3heHL+EmLEWYza5Z
o3ub4fWLkp0DTH+MJFeqQNa81gakUI00CRWpU02OTLzBnZX6mr+VyYK9z7rXpuGMljP0oNycEhx7
4djehPMctbAMzn/2ngRUfy2VGeAL0BxD5HN0sct5Swqbjnk3stJSyp+DBoNuIGfEOp+E2pIO03uS
dj54eNZx1IRgDX2YMBtOTpXNFx1JaVwDeTW7tiOjX04obdK+qVVCM9qnSTSaluFwKQJDUQOQCsS1
y4zA4UK3pBGP+Z116Cxato2qPfOBUZEvUqqMze7vpjc3y3UUqrVjb+uWdlopvPwVQx6Tt47kmlzb
rcYR+TZYRL3riAnWw620CxFjYwrsuaQ5JwyRKJGn8L1zHCWZ7W1kMPdHMuFRjZeRajoQ4sWukaCm
PKA+PRwtn3ZfnoyfwWPHfxxkIlTVoOnURuNCz9/2twII307KUSq1E0nIhoVKHoCPL++Cflb8FfRq
3RagdKYn9cAbTaOItIMq6HKd/VCMGOlQkhlsrsWbzxe6m033e4eUnhy5pP2xQAq//Fpt59YdFaNs
pMXU2c7rRTguV9snlVQv+mDCsEgXzPIQ4+HFZQG+0q+p/BoIRWBtQgVbQs17OeTI0FMb53vUzS1c
8RvjZoe1YMyuXntEliEcU5qJYvDNmMYKCK7n5omhGG1M33yaSny2E9AHSvVRgYfqjOIH2Tkb14pd
W6uZxWhbrGARnQxqGIgIuuYqvQYD7JPKgjPAfNoZYQlD1vpdiGYWjv5iqSMMMU8IUa/N3+1XVUSP
jbVbxs3g0RmTxxEUTu6owdpL4ZLOsVzL2HcTx3onNFXqxvYZ/EtjlVS/f6p97YotHiapYjzyip0r
qkf/m1XzqXwu2i/eS+4Cqo/D0tpahTDSkg6UztwSzAK54B/Avat4OwKuFYfK7nP/dx+nKwSirGOL
GcakvBtuuP0IAnZVuXoEwaTFE5KS0wavPk8U2xpHPuIsLh+VXbxl4TcOKj3jrmW9Q0dJsunpp8Yk
FetvDgzpaUTEuT7kEDLZxv4BWGTHS8rlyg22MCRhf+zadL/+wJBp1KRq+hlTr0oqs/NUnjq2px5q
HLqHbpZs4b1Pw544iydj671GxJzf9CGGxDUxadbOLFu0yl87iMxp6mGh6LIkH1mNdryKCV1NBBbM
6qBwy4kgnD5ZWoWDM+8yR4hCk3s/2xkNbZNgIiXHbD/FrFfRTDjAsVwGpninZM2ylep6F10IYeEa
GOmClJWEmdj7nGMBnV4xL9z/4W9qisxnvFU92NCWEJbyMPs+I0WqhACHkLk6GjZOHflbP0YeuJej
Df8wpCkO3HMCiovjXk1wl2BUm4vPuGyAOSobDS9vfbsO9Si0LaVWlk07SgIvP/f+i0TGh+0QWFx8
fnMJ4JatWOe0D+O8LDPNTr/bhNrYq4s6cKZCWrwSX0prIa27Vx/AHsffuScGeUQ1J+WnxcD4RpDD
TrCcJ6+AvVb3ToNurr8ZrRLODX/seGR89VgY1pbVAjwQUC4DBzuBWVQ4odPfVMLu6Rmfc3S0WuYk
JbDz0dCyxaBZ/4Q8aqqop++L2H08Jpu+z8LPmHU6hKnQe3TZgJCCE6CJabS5sI9s8K5Ikia3jvoK
ozwXHQumX0HitBKO0bYQ7DFFfdrjQsN5irzoFjFO/WhISiBUf3OUp5G0m+Gx1JLICJxO4azY1xKM
fHbA3kfBrtdqbgqMyvsbALngHll1K8YAFRnoZaThxlYYsXkiDrJ8JT/GaYnDpKX+YBv7AUOKhGqc
jz/ko+SX2D1nRDow81KzI83mz/bhmAet8gUu3DmHW2b7jVPD6f0AC82Pb/JpMdpbAj0c6K/5E7eE
ZN0/hUXh/1gzJUCjYMjECyn9ZYhKzJV0rh3tCe7QBTVBtdQGVARXlbcL3M6AsxfKf1AZynW7qOZD
wxyo4YuRVWxkwU+PG2C7MD6m5PcpKpHTWLzuJPec2tkIUw4kxVofeKc+iJI1y1xLWMcoGCwKN0HU
YTf+PD5RhlqW1mS/D5d/ImHvlRoz3l0PTuNzfyEHiN1KYeZqQMIHTaubymVWcWbWyHPjogETNJL5
pWIoDREwN/pIXMe6xz/1Wcxa7kKlguKVAppt4wHnzsjQE+Y4c8Dn2PrjpR24YOZk2WHYdh27b1oT
rjkREuEVl85QqJ/1RK/O3H2/iGAoVMpouGOCxcPgvDClXCbwO44MU29cktS/w1KxMbycCDT0mAuz
lbFT8LT70YQDuqVz5Fjf9Lt/zm9MXBSc8zdUbBJ45Wy/t9IFlxk5BHXyG8NsEgtbS3WZiPoX9nvG
PQDtEaozLIWKeXapmMwZRNrS/xXPohZcbtFAWv77i0CnvG62Rx7xGO/DVJlgEdsc1tiMug8EVd6I
SE0FF4GFodbG2TkIsJ45HcZq0x/vNW+ofPyjewL0PdbwDF6Fhne2yDGmDDyx50c+174mlrgCUeNL
+OloJUS1KN5D4rDKqj3PFQZbrahQzbBh+qJQJaCy8bXHFH5VOldvF6GJ8nYRZbQ9ctun+5/UnVY3
wZbv25EgLHWGtjueqK/uj1vyRtPdWaaFpdn4cdufMp8t7TjR3w7JXq0LCS+YEH73qKFXVIlzbP2J
Kj/dggMM7DPwS9ioIxhY2/vtr7OlgF/TrQTqmmJbVwpl7CUC+nX5kVkcN22/fYAiqflG2GPuzbzQ
oCAQnADkhZHSqZKaN18TcOkmxWfQWc6VD5HA+wH50XaLbEE0BuvMPXtUJbE42866sVxNO1iq83gP
81hpV92DETdadWtNL7ulp5/SF+cnb6A/2uXecPIroi6jQ9BJ5I4e+noos/djQZntss5TdQs+gDF1
u8vwJG1baCvWOoTt/BItjoQdRslFlyjVYTx5uow+8jtT+vo77TOrFDfcuvkpqCtuXzU+wCv6ncRD
EHp3C+54dVOL0ns8FGY9Qc1zAyLGhctQ9B+VZCX1QTHIo9Cqhlw4tozfKaf7SrJ2HTNwLC5zXMUT
DtiFrpWgEgZ5eqCx/ld18HThMoy9huXYb+0b2i3h8F4Cfv0Ez860fpEiS34UC5mt0Hu5xE6zpJWd
/7ue+foCPgMCVZj4EYt4O4ji4lKuRKx8G/7zRkqb7j9F8M0iLbdNr93ib5pVnubSinu4TpAByrjq
c+/KHuFmKUADlU3QxFw6mrajRd0xkjtDN4QWpx2D6rsKyFqQT1Oj/fCoNFbQAWjYcai4S1++bNcr
ZqVs0sX5jARItGnHG8ClBbBkGP84W3iJLV88bVHHg0nukItAx4dYuqqylUxHnto6ELO5A1q5k6/N
jlgAgNh8rWDwu+0XcZlZnb14rG/CdjrDu3FvGLUuIsqSigODR/pKKocc9MNOG5TLgBKDE1tmn0YM
OsSYtBp8hLT9JxT9MJpFBKstQLToJ0xyD3ptrE/wdn50DX+h/pDsk1ZaYOLE/+MVHDiwlLZm3hSU
aZKbFRu+3H9RBPuuB03ddqN4oys16tHdcxHBBXp0gUOEfNQfBrAtnvkn6hBNtXp6Gj8Zt0s8YfoF
IeQWjE3I2TU10tK+XZH/tUiW0YQimHJZSEVB6F7hb8wEZpk1guaMDpaDPlYJp2nI0EnRh6RqYphB
Bqq1/8oD6B27CluAQF6u8+1u2O/rl6h7DYTqj619egXXd54lS5s5xnpk6GQcNuB0U6cUo+ykahBJ
Y4zQMG/d1BG0w3jIt0Rfx0Tn3gGDmAVBrlAtMaNUz8KXig2Ngy5bcOKhQfd+zt9PbwlUl6cYpVfW
V20DgzmsUE0DcTzW9EvlldiEnvob7JYYAthpnY5PkvxT8fckkMk38cQwvuOxAxmw5xPGAD+4o5YD
iKntlZW+UuLvgER27Nl/l6Dy513Eo3HO/M4Z58rL5UYq5I18LWNRv7sbEsTlHaUL1jfroaSsorjO
9x7KnwUZjQwoApQT9B8noqaef9qGUu9Z2FTfloG3vhBEMABatrPeOGiWe18e+85PLn/2Mdq4Jvzp
rcArw1hJEfTKVu+Ni2bm1EdYoX+8csErZftoVV7zKl5g+7uTdwBGOQEnN6NXzP5CPCNUvRBdPG9t
QvIqF6SqrQijU0VztYPDbgOyWDgx7o8bA+stFMGfTlyEsGvBAMeF4sCmaTzDMioTSgn34fHmtCrp
uhiyCRuZ3DZ9GJUitC25fic/Ox0J3aBsdLFZfaR1fyCHlIhnSRlKMzyo61bto5xLLN/bR13QgrhU
qBc2LKQ/gxpLxjK8HyvU9gJih7mDFfsvgztSW6r4IW2Zbea3WUVcV7dEN/3Zzi4Qng0xva5nlXpP
g0y2Akgd3N8TDJNPSVac9LsHG1dnqJg686SMvQFpxLMA4iuzjFSYjSTnD5SYe/LBEK7V7z8RtHdy
gwRyJxzSHQotCu8FrkQD4gZOzDxqrk5jWhViqvV8lvZh7gQ5iL6XUn7ue/cMEazmKwfp0ZfkaMxR
UgSTGc5+GY1FwtBiAlYn80hgGLB2p+58XNw2sNqHAsR5BapVVmSvh9VUtnPbMsFMHH1nCaCEsUKH
H9FLG8CMvZpFYdZXn+/CNrVLQmhKtalkr/kix0XOmi0LFJNnqYk27la1IoOXRShB7n1gFonPYqSs
VTn8XsdneeZGyjdeXdIjOVipWHMFrNvcnVDBn4foKG3pcjoZlBpWkTjej6iiV0ILBHc8Q8+ly48p
OkxsQKbqnytrdGSYBJlwH/NnMiMFu8vGTbe8Fkv9p1oCENxV2/051exMeeBu9yvkV4uK6eBMzl82
cKKyl+v9uX41XxoZcORryEMpkqwluRiw3krP7pBCGqTPtFQWaklhGwzWks90WZX7U9KDGK87N3q+
NLzfGnzahje66cErYNnv8seSte33KKDp5Kb102Vczjyhy/ZvXcBtEXeIPdoP5whvdVv2+MMtio85
Wyi21Nl/+SMYvUY8mFwI5g6iEkH8TtpjiNAq9DrF97mn3AiKQ0jhl7Xi4oO2rA1FLjKnpnW9gsos
0sAc2j4nzmf3O1kRXZ3UF/IxYYMDp0BQac1ZYKyXx5Z7qBHc75nZwJZN86v6z2tZPlRV5s6gQ/JJ
LJg1fzpHiS6G7YbE9jYsTk2gxB8GaQQVM6oUpZ8gRwgxw+yWPOd9A/nDf1kFwRk9ZXy9u8N4+UMn
x7Cbg/Wzppo+fwoPNnseMLxRUz0DEaEutQDRkKsxrRaPJI1/FVnTUE81lCNI65HtM7GG0/jc1SQF
Ft1Si8st5IuPuZ6hfAWB2QGAZ5l7olvXMmKta3kvutU4nFYNAlIw1OdfxnC0cBNuH2QQOy8dWNUV
f8zrOuzAJUvI5jmIdf77HKzKUJY2XCmLUXkAkV/43XoE7Jgz19w49+1qQzEPQS3BsLgXhI9FctcZ
PyJ068oHgPmRii9fIp4XXTNQsX+xyAAkLiRo7rGvdwo75c/xg4p+q75ld1hW+6j7wFoLEZd4Hcpx
rwoOYG6av4Db9p/ZixoTZ7nPqmahlNi229s/P5NC+tQOGxIrDF7kVvhGDwxGWdPgp43ryKgDZ4Fg
tBuyjFvRqUSCX6oou8d+0zb89RS7IA/2vfFmXu8WYTh24otI1+PMc1b77SREplVCw1Hu9ceamqus
1EdYoZQ19eZxRzovD+h+hPUmFcSPrZz+l550dQUA5hZtNJs25a+9PApeod1I2bxnmsmF3a7Xi7Fk
RuO/DE56HQSwprIE/lgcyy7k0h43vQyeNejj2DPobVTKcCJLKqD1dVvEhHyQRWVy2NcQBs2SPU8v
Y66bHSFHGOrysEntQy7wJeXLp5irOKPOv0mICG6oxg9V+EKa23l3l2cIixWONEgN5uEXr57MdKlg
b50z21GKKPhMI7iJ/76axeNACrfnldv0c67DYxPF8qdkSNnUhoqmkENFubJTEdGzpWqwx13iTTf3
KZNus9eQ1Sy1LauQqNP/kxGaxwdAW3ZCxCi9qfxIsDWcwcgAy+e/B0lZtPnS5+v6z01HyC/OoG1S
tF+GK9kOvj66Y9x5bkAx368DBPS/Guv/Fz8hD6UhIxAP+6xXcdHZiblOVQNy24Wukqggm58IRc2x
1xffOUVgKLCBir+SWH4oX8j9mtMVe1Y6oL29TrKv6n+SPqGj9MRH0aWqcn73dVxvXUwIblh4yHPo
rk3sys5jjbdU+SmlC71hrNs7JIT2xM/x5jva3uDBrMZsXUn42gcX8wqqefClnJdKCMCBCFktT53H
aHJ5xdgnEH/XIRNqsjjHZSyOy5A2yAM+Yr9VvFLr7efxtu8lq0kNoCrlvUt6lkM8rQ8b0Rms20ii
6E9l4mTAPQX9CTdE6gttcFf2Q6BeVx0f/kxaGVWlCjbtKBEYkAw7yfBG25q+3mJCJQMQ74pBdIvF
HtpOP93xMBCyzdMaX8fbQH7dwt+PWyxJSET6RLAKJBMugO+HaVRxGzW50g/6lEqjzQsG0K55FWe1
HOVTViuWdYYF9hP6bntIbKKQIEJFd+h5poprpAdRu6/Jj7rCfsLIUXhG3u83dlyzkCg+nZNN7ES0
m2iVk5PsLtlmsb8vDFpL2hrU5SPR2yuCYteoJyUWfl//5DB4nPIaxGB9JgtnzYix7EnWpegsGOl3
7aAlcopPxEjZlEHZ4bW4KVZbX8w9dN6QOQ5GwaywNn2jReGkQIwa62iuVlSs+qnBMw8fVaTD/Jtq
h2iLfMAawp+E2WhoD0BYGfCJ+/89bTRSYe1tIuyg6UDGFpW1oNatwuY5U3cOUt498kMEbzWNOTjT
Cw5iWdPwKEmkuVUdBpjay9+7H5fkgg8DBf2iHYTwtMRNPdl6oOPf713YkMl08WwuvjgdPjqxjhdJ
IWOcjDRBZwmxwvie5TKKZP6VlPTroT+PNxk+vDDuVTkLU9AnH0WeD2qP9hJqVRr1HA3Pi1GuD51T
m4zLL8fA2P+XxcNFq0QzNIb8hCt0dHJlHswUdKFj3QolR+3c9R2bbxnrsmWK/t6AvgJbexSTiqQI
DIqv3K036zxsFSEv0FbiCktyfmJKM4//9VOygEDYg0IWtmRaetKundb9a3DLIgPLOi/TV/L23Hh5
IPZ3ql5NR/lTS8SFN/H4Vt2gHdnY6+hnIOILAfo+ttxWG/jO59vbTuRl3jBY7fD5c5s4LaeyIYz1
HM2ZVhb7sCuQ9f20/p48ojh5596Jt1oNaMzWM45v0ea8EBF32LlN7Ft9CC43XsepJSbKJerMz4F0
8DOfOF5/Ncje890a5C1jM4cINAZT4yB3U6TzTQPRdOju2e2zGVNxNtPuDL8anYSLTQ9JS+0boYmR
vQ31SBm91dZEdWzS+gdqUx9FEuTJ8knFHLmxo2dPnW3LFuytv8LXp0p6U1PMUFFM26cSPC8zISPq
qEYL7JqAmFi6/V1un90T4IIP/8Gf1XiBgV8kD6UaPIWfG3E+aaG3TOKn6oUBKo7ag3rgzN+dGMqh
99Q9dBk2Cks6wB2WhNAukagYa0ywSi9KG0z0zKjQZCZmf/7zGxV4BMgoO6rcW9xcn3czNz++VRW7
1Isj2zTg+ARuc7Y1wJFcnidp3zJWP33zARbsMJAP0z7otHbTeGLDCkywZBwYebTTudjaDwleaiyl
pZXhCUF66fMDI915uJQXKh3VS1NP6MJ9SUwMEZVj5EsNn31iOvCz33EnJ5AONFffVZJW7UBWlf2j
8hjptrMPkkX8AALSNcU/0dz8keyI4LyarvZLT492lEH7xNuEZa+qXUWjPU/oHzNfJVFX+x9LBIUZ
zkSy78aNbVwQf/G12nMPlaNrcTLtvwOWbM/MdZnZIKJKl0Jm9qtAD0RBNUtKb8Za5l2MZ6Bzp5XU
PmgC1K826RbdLqsqD6wPaSC/1dJ/76izPk2BTw4uNhs0i8i91KNKtSW2P4+V92dZBf1YooKJKGxf
TQ8GPO9Ay3OT5AKmVz7e53KA1S4mJwT9fSIZOyGHyBbfp/ZLWTQwvsLQPTWI/8VuELsABmW46J1z
ZpikxJjRKKtoLfCYi7RCHy6ArD3I1IriaftLfJ9JNzyPDRLE6S4R7hl1vSVhAJF2TeSajsKHexAE
JS91tF0vQs3lzTnmGrb7YZRFkMdrQG/GGp3ha7cW+ZE/yoBSbQzzGv1rYOOCL37cjmttdeslE0Ah
2Ybg5oGidb6O6gvmmfaKpkk3pTMizOn+1KXlyETaq7DkqgFSHVE5wkt8EMnfWZA/iYfAYOjwCY9p
WKbEeSAmDPZZO/8V0hSed6n04+e0gEfWHfSoa460KOi9X1O/Ra46UqZi3Nxm797+KvCDM+JICCyq
VaRdV6JXDgEPyIG1cmx8G9bKwRatTFclNCLAhP62D3k181SmOUIEkMoWrC22RcOGxR5vHBEvaez0
TZkmfKjUziQDEy/+BTSTEFpjBDQcEUZlP7sV5RW9blSJIvVpFWQW0Onc5KOHHOJXBSQC3XnNOJ/L
PqJexxar8I2GLcT3lAbrABzacr2uCAHl2xf9s1d6UFY5vdhQqSbrCsLcDlipXkUDogff4xy49kt6
MhV7pfK3Uc8ybIzCxjzshheFjhSjcYH1h1r89zDxJ/Qu2TumltIcLcZp23+bwpmhOJXPBLcFZPSY
JGJkjUCHIXML6uOWL2nYFDihljfQMz3QjWv23vLSwXrQSM5mIkFw6gu371TvN1SnJz3nyIWUURdq
LVB9XoR2cCjqVZEsfyY9cxMddd+gcfL61R8e+FEmL/LQMmD90bjzPXtuEOoAwrB3CLtELSzcDzTg
Ht9tv0XAufDCfDouiWddH/Pi4jcGG29mm6sBFfIguiiIhcOfskS1YC9xdlwtSRfdshI1i7hOWt+U
xIPxW4KU4LAdyi2XvXrcQJ05O7IovjXwFmifUi9afstSdmCCtf9DgHDzauyRMSswFloD6+0Fqjln
26T7yF3bZGVPDUl70S1CViio2a3kLvAPMb/Gn8aCuPHmFajGnW6Rqa2L1inRACzgP+NLzkD0vG/h
dh/EVZUEzN9rqkwfF/mfSQVD7JVnARwIYJ4vU5yTw7jDoSdCfQ0q4u+cAPxruJrndmFYtbSQtkIs
r4rJoXaf+P2GDRqZa7e2PleehjogLXDTw+FexnLBnk09dcKQlUIP5UfCwK08omo8KONQl/5VDcmB
zNkwkRiriLlqO+/ULmmoJbJUSgMVbfRCg+wRazFLOY/nyOSP9WDJ2Zkt1VbQXR096Qq73uwWvub/
YDN0tqBHJYQZsi+PasbWJ/YNvyQNEYfvFn8U0AzRFLSaUJBt51eS/f70BiCV70SU2iQSFyqgoaX+
ZSG4cM8m+0KsXdehIdbOHX+xuhebbFUqqtQMIRZ7/KFCbzy61ahvY0UMAeHD7dMJTvNn14+NcmWo
zF7Ay8SbsY4TT3J6Q5DCthxBGxvTrRGkcwPjD6T6Ro3G1N2nGzh29jOe1K2f7WxspFXyTYENbNDe
5LVNZo7F984zASd4vsy7dzYr7YkAF/VVO9ZbLsUI2gifFRkqBlQrdFEaJNVDG0cApGQqcRrHeklH
jNrHi2MpIfub2X3TyLGJ57NsBw86HP2pBzNfYPxu2cdZOLWX3pO23YWQcv4Sj2u+8pSVOkGoejlp
9YsMFtlKXSUVkeMNfna+1szYctzzLi91RxNlP1eZXoln2HNtxoFbIl/23RqadIpK5Y3DJwb4k6k7
ZCQE9SEtJc9/yOYKQ2otT2EUqp5xHbMzaJ2SQ6Ukj5X8RkQ1v+N74rYCKqfJE8gHcktO7RojzMP6
e02y4xx6irL9+uYBYoHsVUuNtw/YGiWxLAbOR9w4tn3oBjGLQT3gM9IH5TMhC0o68vyCd776akac
QvACRFR3v4lmMiJPXhzVTEqQUyoiVocKIGrs2/o9HmvvYK4WpefMCVoFg+thiYY9OIfVcCO/yfaI
uc4qgrT75G8ba95ZNsOxZmNwq8JRb/52pd+M8om0h+ghN7iXPv8kqUzDSF4Ti4vQ6SUL3mChUNMv
2IGPOvasCWkclqGwSTzVnjm3gBZJVN3Ytf2zcwsvVwCWHU/Xp88QnAw3s4+JapcNSOnc67SfFUC4
TniSHJJBFvAUWLxyzYedHraZuhpPn8uBjTGFJJN06BHjuPtP7KS/6Psz9kaJtP55VfhcbhoygYzy
bkNaUlokdUI/+mMLaWM59C37m2IC7Kad6Dj1AKyK8GnfSyRCaXhNT8+Nj2j+iSyDFYvI4CCYQIVO
LbsQc6Sp3JXwM7y5acia4EjmzC7Uk4RCBbEkTkNPJYo6nXW0jOgkDpq84AANFgRBaF9zx0XsAOY3
yRNYxwdzUY+g5nc2WncKGtTUTkarqUkizV1u0TLmGAjTwsdDlMnweGYwfv/+hs0ZaZ8XV0cXBbHe
suHUFzZO3Plv+E7+otTYaSVG31UpeFEI0Wh+YSCznd2Hxcs9sUsE5P1r7GkR0aXpTJT18RpauXhU
OOXomtfZ/4AIGVSG8NhU+zbFH7tbjRifTkQzXBV8NDQcfuy3TUiip6ePchx8KDT50QnMFdylCOaB
HhrVdawGXKP6b959HS2SVZb4Xg2zKZkf2cSCSKJUMLHgr5iij6AmCgVHsJYtJp9tOiKPq+b/fQTF
AV/natkTECy0FDG95oo4TyCaPOrnxtJck2bW38W21U4r+AGxYBzx0h85kAvYkGD8z3VwuOhBu0Bv
yc0R7lO1wWT2HKWIrb24io3eSgENNW18zK/b9E+/pnzH0jSrEx9QsYBlUbe7IJ9knNw/hqdQzG38
miSTTr8yiEf68CxJ0FiJ/7PMsNb3A8E3yMyBoe9gwR1t+LCyvsfTWoqG8GSPOVaFakYFZhpZ+ZL1
YczcQxwAtg6IH9finZfznvqHqGpHIdJzlOX9vNKR+wCbUI8xqFO62R6+jhQ89cjRgcRwzg7B+cyW
LElQ/UHIz3WPr03NqK+6tQl6F4o272gz7fSKBXnpC3jxXC7FW0hwsC9G0q4Qiqb9jwPM/+0dwVw2
dZ3BexL+1D0oCxadvYyvJKOntLcZgVtxHU3pTbEw5l86u6152S20K99FGn2om/+lyQHqXugX1a+e
Hd7XGwr3e9hHEtbEayZUp+d29nII/AoeIHWWMSuTkgUqUJN5XRd56+F5FiXKt9AeUTbnHzPc5OOU
CxDaunClEpm1jAeDtlNxqPlw+CDnqgVIkqGUQTDClJNyeXjL5SIk/qUBfkGMRt3csrs/5gknvF4F
S3CvlAy45jmZrwDtx5df4siZfRl96YJG/xAXFnuRPe4x0RgO8JapLtT1jfcFK0vrnokpuuWhXQ6q
zkB0IDo/UQABhJzG88hsJ0L3KBoa30r5po/9zS4sFWD/CSfOP7BMc/MdcjY2jcYdIuJtl3nTFT62
qM2dbN0zW7Q/Ww+4GJ5lhYb3ovMUtucN9VQy9PXD/4z08jumHkGqJCohNo99zNF6je0HIClek1+m
EktuPnUJGYoEK325I0khiGt/f0OeQiYv+ZfXVxFb9Luia4KsVbnnJIrM8MygDdVcKbw1xsiCZfnF
s5GmRVEVC3i8sDvGCKj1IpJa0wSRBmg8yq0ynHaQRdZfIcX8lV1JknM4Dag+eNHO+LY9n1IsKDia
UzhN2A0Cj6XraUmL/dJAk29qO/1RuyTs1xPBZJaiygC4PINYBWG9myVhBQirwDD2AQ4MQDDH9Glo
zvfnPIHyEC4flZnZTPO+c1L3W6xQNmho//wOKh26YfVz5RJJU2g8O8q17NDGy+xYmrQnc7la9LfA
Nyr+5yNGIkbBYNEarddaJK3jSssES6z2keSwR4txxs8WB86gSeiM9laEhmwMKqAbSXNG8Sfg1/yd
Ba0tyoGOlh4C4LxaHQ+0aDNxo6cDi3tH3FcLHFKornptNDwTgQg6q3dRG3rOx9BIuWh0KRq3Pwcu
0TjikQMAAv6WNyoAQg6GpkCnBfQpOAygkjEOXh+4e5eKQfJYgQF4KW+f1R1+KfGdIMG3fJYzIbM9
tD5v98TMnPVdY5iadjAScOCO+d1jwrfmsIKGFRf1L8PYqcek8cD5T0GGeaanOcnk2Znaq3x7KmwM
dr3OczlBIj4sozmbtSJxgXvoIUQ2WcY9aS0TwQniTKCW5urTP/ib7PjwRFQqKi3JmJHgcnvOsYIl
pYf2bIbi7koq8hZtMtAnkktjfoX2Kljp4bPDkyvZd7Iq43gmjg5U9Qy1+b+k48CA5/Or9LGM6P9q
Czy3+ACso9uA6zFnZUfy8oV6JXYooPVZVSjYl8qmYNYGV4ifEFlfwsdpCrC8YfxPLS+zyNCXD8pu
6c6nJZNOO+4JJnyVI+flFEZ5ophlKlpTP0Nyl6Gia1BRgc5qD9gkXx92v+v/z8czPVVFAbJfhdiJ
npUsHNLbbRgdlNHFkbjWcR9T945GOrrzTRiwplST+LAeG4S7mKtj7OD9aGP0vB/qxCQZCi1twqPW
VFrg6JmdlIasqTl3u0aV1b1b4PG0V/uguqk7H+ibdBdMyiua0HyPB2CSIB+3C0dmtiadcVyT2p4D
/a2kkA9f8Zj4YrFCxJmPY+Edi7skJXnaY/Vzq7nq2kSA2qehFQLtkKX/Iqn6GNO/jkCoOkp1oO96
LKWaPKaW15h28T66KyOjy/oh+fhK/0A4W3EzVOAXu3tjp+FrB4HgiTizqv7PRhS1Qt3nXWtqGhN/
FshgeC74yjL+xtJw/54WwAeCaVa+fgTVaN+dSf2x0YjrMktRDoLLavaIgsmaWNs2iJm9oJ1YlkpX
ZlKmNR+N9XShyelKg4+s+L1yAqWe7jdP6nI0F9NdNXAN4cGBi9wOeaU9urQZl15ke4HLk7zZwO7H
ol8XT8db3kGNsIpxrGYdgUpQ53xZPbaHOvsonqaRocv9o8/jXx4z6Y3jp3DyUM7a9f7dcvQhJyUC
Nf9U2veV/dRYHOweTQmG7MvqstOQSS8oYMqdmXQ4xBRcvPQ81KgZ0OVA8FviAtTa/qOOO3sE6FJW
piAS/6+aYthWfaLHAXRl2dAqpSa5PtM/9xWrCeByYjw3MV33Yt/kM3NI4Vx1xFR/ph6icqYhFE5s
aw10KwhJGyEnVm87WKfu7mCYoDZnbahc2jhV9LAMdNDYEzQy7tVcB7rhEUdENEulqZwVoxn8kOYF
qjW9SeRE89fk2y+BJi0eCauQ6sME1F0BXbhMrJBLRlimlnq816WD79b5waFp4QyK+s0HNQ0ybm1q
ISiB+ZaTRciXq2JC3GTdRV1f90eJf14BA09mE6Vj8b3GyB7dxV/6NpFPjtEPctYTYJZ6Qj/1ChXz
rwsfCNre9pqFKnj5NKaR0Tw5Ah3yiW1AlFkamUXj8JCnyMS7wk76ztUtfCGCchN2g8xmFt0LoQaX
Hw9UeJtEkAu5oCzrgL/X5qL1jENuXBftqGDGcHRUXTMGvOB443VZ4ghfJcFl8uJlJGP5m4NN0MY8
18LeRfgCixTFHasTzNF94JqdmzIOlOfO8/UZrUwnYbml2+Afa9hzr0Yd+BZXNwt+QCrfnO1/6X6u
41P+tcOvHPVcnKMQn/v9tVmklRpytfuy5ibUTlsAN2HWg8HEYBHxR4LUgu5M28I3DHgblGDgoIPe
sUHKYpwZqGHdY4fvbHr7KLOV6oiYJWGydRoAQ0AtXVIhpCK/6vCqQgWKv7ADHM4G0FnyMJdvDeTU
Tr3FXiZYrZuP0gTs9xirEOxXbECcf9+Pg1y15BaA73g3HdHCcGvdkanoaTCJSmRr5haaXjFDfYhy
fNFVp0VziKr38i7Yg8RObLJA+BPnc2nc971Gm4+RgZGVlvkY1hhHruaJnF7Qa27q0+v7aukSZNN5
3Lfge1R6DtrMPqm5HjLSIz1tGAcNMeo8Z19cwdAi31kLTpoYSe07URwLpTHobOr/FVkU1keEczCc
FDaRHKB8LlGR0PPWVbIDaRIAWKQPFAR19G6BGFVMQB3VPMKy4UqNj0sUDs/vAxCIxlU1cxm8zq0G
wZ5foJCP6Sxy3xVn2xIau/OnQ9Av+uquLQNDS8Bk3lk+wGLHRXEgvJhZtFBLyHU2yMLXpAiClRms
PnIIh95Id37x+KRz1a0VKoZEIBggAaVEYJ61G323S4Tq43AMucAo2eFzal6DhDe48200KAhX1vEz
2EYOlub85GEJr91eCN0MubVK75jSTHNF0FjBT80VUwc3AQbrBv+xKZpQw5wSTcsrtPAYkWCDXlRX
UgFeMS+t8CK84KepQtProZCPyHGPT3GsC4q1NVyPQpHRu3o135SA2ep4OZI+Imd9ctncVJ+BbsCD
NuSpUWUgUV4IItSCoez4sVks924VepvLmSoiy2Lv41Ya6sw+KGrWc0Z83RSgfuSnnlimoSR7XZ7D
ICR9IzkQQFKZg5S1FKFgMOGm0w1BKC3NoB0o+k8JweW2Kv1cWn9cmzblhwv3xdRWMmuxnjS1Gfhf
0g8MYE0ibOewgYn7BhD2el/5lV3vExC9bQSIGCJhcxf9I5iaNdO1iDrMEqVvASQvGtzq7Lwm8dZL
GjQjz3aC7TZVQGyJLc5sEm1pGlphYlxAEC16LGt2EBlMAI4SJFSqWEYfoscMskP4NcDkeBhzBeJH
tzpQLCv0U9fmpK4JV9wXlO89IPfil2405qWOmaQCG8T5Zmgl5TVtBM5QIqK8i9SofgdRxIRDEn7l
JL/12xkKroey4vX963WiXrjt+KveATL6MUihFMVfXPfcTcck1fZeDKYpS0oM8rfqVFmygITQ3NY/
67aZWDKfhl3JAYkkSsGcWOGITPrwpQoF+iZSyasWdQ6kQaZPQQju+YmWhZnCljnzu0nannX+xOJs
8DO2yI+XC5p0r0TD3gD+LydUtgZBdSjtn2YYxbmIf/rptHreHVR8ANSZRYXf2/m5FZ0P+anfXy6A
ySWF2gl/MBWlVYGX/aeAKMvRY7HlXCCyU6yzwXpDBlFeYkQJh01yAA0bqBTbsE2Frf1B7ktZj6oY
LqAIaIO7I93UW61ISUyF4kGK/cFP1WD3O+3t5hmY2yFQdQ2lKckVWo2rgAbfkWknaGc363YT20BF
7/4OC6jUm4biSfT8K32G5PCKYgBbz82RnJsJaoc//cKKrYkFmy33lXVL+mv3/V1R9Y8uogYEyTr8
rmYYn/jvt9HArKJXhkMbySDo0lJnQz+OJrXOzIZCyvHc8DV2cQgBNCSz+wkqW6MRaii6IIzvanUZ
mtR0Tv6+Qffmk2gAD0qW0DTT5SuHQcj5+uajY0zfgnMPguxzkjW+NHUuz1Xajh5vM/1aOnLDTume
KMvTka6+FXh+pSomBNmOJ2YN+KmAoWRZAtvXNmrysBaR3tHSZxlHJZKXRWV+Ma2Q3fAs1KV0iMy2
IZK/VSV+7nQR11aJkLrkJHGusgk+6VaBR28qf6GKPuQMyZqrF4uci6B9OUzzej0eQhdz/jvKrmGe
MKQQ1ldabv3HL5010EDCI2uCekpI6ozQE/i18IsQPp9nkoa/sMLZ+rVyoFOZXPfW5+gjEKCbMHst
RpCP8FQtj1rjoqqFuAwpHn5YfQ0uXKOZDcQZ2nqOnUcM3RfOcqp6VwtfVZadOfEf9dVmfyN+vHN0
+ObsmOVoB3o+e+eZzNNzsUEB5uEmTL48pb1s17OUPC4EP7sPpNRXL3OO0eA6pbgT/CLXUAAfPkUs
LdvKbIwt+dh/2c18b1s2tMlpF0XlUVS1RygvgFOlA5yJTqoHX3cNkelX5j4izg8MaSpvxeMSgNA/
tzjboTbvnaBKR+CSvOPO1kz9ixyGBqve0fl2yP8cu5HR/JTzvCWlKQSrTJlxEbYsnOtAHWFpHebW
vqaBmPQ2Q5V9ZZkjOQ7Bzuj/MzxVBF35txfFQDuBVf7fL87zsM9PvE6X28tqXWM2yuctUjjzUaqb
eKfbtIvyUO0vRTrHzawGHgPz1uXzqLOtCcNn8C3O1wOZ9759zyIM1CTMHaH0+BPzSsxp6tDE6xtC
G969woSxOVdTSnzypwaAhHm2VFVdv0Oq3LoZxVDcoCVD1bpBH3E3vEFj/gTkxZ+ZS2YH0xq0bk9N
LlL7IQwkwmVjVItxiuHh2xAHrsBwAF+4RPR0Qep2OLzFjw192s9QOUYS+F2dfFUN7+8sfysmK3qz
XOxUMAUGIBJ0TwRd16NugThN65hd/OWJdSP7CDXkGCi7Ni+LCtwxgsL3s+b/9KVwmFRNC50wildg
b3DZ6kBUe9r2w2ZNzFeIib5CEpapNImfg1u3LmXCgTwibFHsb5uealtKsBupHa+iOG3lAWS6Jkqo
EjqUwLnDNknWT2lq3PVDcSFt4BEDRYbM/AxnxmNi3fIIYWi6nJb/TavGj36JGQcHJJZC3yU9HI77
ZoXcDliM7d6p5r3sDlVvH1Er5fMb2yDbnIImZqNMdRzdw6AsEFBg0J8QyEM25qIApLf+Rnu0ogT7
9cXFqekwlYAJLV3CTvQCYnu7Gn8YFnMriWEewCCyzgZ4+qqGvudRni/OxJmLy2pmvEEMq4oZ737O
lzcHdETSFbyo0mRu1kkqXxNTG9yzlS2dWKzeR48A3Td/9xpz74NGLXp1DzUa6o6CEa4QkYX4RD9P
LoCi2hD+VF7PfX4RefkJW1MtTYXMW04ux6sZ73iE/s9a8CVDC7K2DWDOTjOBoUeCEfoSVJN6FDlj
/ura23QHI7l1YzAFjrd/s3PI98cW/dOF1Y/4zAUbGj2Cy5dhGJYyd/vq61++6/tcCOfX8kH6Ou1n
OkzdJ18FNUf9vhbdp49px0jPZg5vXs1UXVMArC4ESRgArE+oE/sqFhDylEdc14//Vjk8WkfGzOmb
0tUihPSqyW9MeA7+NN4IWJJaarz8JcYU/VpcHq2l10LrwfSttcldvB1jbRQjXebQc0o8eD+Bq08m
qSAkm5EXMTnBQrMoYOhMLIrBiZgXRgWcNmWmkyTRNLnT/Qi5Ayz0wYmwQzba6dA85cxHXixL+V4n
hqvvTUQe58Cn+Ud8GJ0LcePQGswBh9LbttvfBO3TX1sjFyL5PBQ7QO7dbhuY9X660KpAD2MY2Qhz
ux8uPglnnR/gym9Uo8+IeQnTY7jdz2PKvNjPHqqMOecxnb4aohqO05NVaSE0Bbf7RoCwt/apZpti
4qcdnulJPswIyBD2EL+YsJfD+4xgmPUVbmScS3GAVVcXf+vvXY+bJ8dpaCTjba6wnUeOK9sQVvKD
S+ab9W0s//ZfXYJvenkrJUY4pCrioalJinIEzTWiBSzfjKGUKf8H24d8o6HYDwMbWql8NH+psoWk
4C+ugOAgZXMdXaJIY8ZzAw39GRGCOsaBIYXZyve34Uw3PQTZNoPa0MNFxUOm8covrI4hwv0DyJWs
03eQxvzMW2ssIdjRgvkFPp166gZYJFXf4boLPskF9OcL8QdvXVL+uG1nTC+1Fz/ocuzXl4egmotj
u/ai3wp/EvdAnAkDK7h2dWh7ixZon8cnVavcpSLoMLFKPi6g/0ebIuSr1JozJJk1yDshJwcAT7/Q
PNpmZjOxUBBuUcAKE5O5vdgCtBCG9a/wj/UHnwFb8yDejJnyEzD9PxHblV/W08WIV1Rk4c7mJyJ/
/mpAl8yqVAZEKwim4B6LogdE31TOj7cIZFNox7V2Iu0Gs/QNY7xerNQmntd2OM1FEAyldre94DeE
7b7kfFwzadG1fUCE2HX9tXmwf78SqSgUw1O9HN9ERZo50DdC261JOdDKyTlY6fCSEdrJJO/beZSz
GOG/pjwHjJ7iwXN8GDSxWMSk7AF38hnRCrJWH/r09SKfWFz5KIWYkpzJ6ey3DFPMyVYERBGEmtFG
ZNCwfxxfU0KZJToQVaOQZWyFXKUV5IU8mV3DxpwpzCpL2mhGd70nJlUfpvAnZB8dlWJGAl0tnA2a
XnhoQV7v3x+OOAQqYAhz2PA4zR5/iJKa6V9F5hTxR5YNyi3IH41PeShfVdNYmIl66u9tM/mPhjGz
bbLVSuOPBbY/jRGabycJ30bkRXrB35kqDg+sSlTCfHaFFhqWc8EEqaCz34GLjhAMHb9yiIy7rb2s
I505wV8ip0vL1j8XRok/GGrz2I9/jllPJj2rTgomIZZX6f9OI8AcYDBEGQuCD0JX3OHO4KbG379R
REouBbiB6VinRtmTVV5MoYO4vF7BE2hGFX1uLbg3phIW9X+2KT93xmyVmMD8AiBNWD505E3Sppny
IjTWYFqaTB75wWKvvRs4DPTWam1U7qf6IQ3Cckf8pbdTZhtpfOXI0FM60Mck35Oad8LVc8lOa8vU
TiSw5qYW90W1EAFDUbFmia5PErotxIuMFKNGunNQOna0OLFDi64NxKu8zil8WQx8UqakiJU47YKv
GSPFKBmjNiazvLikyWu+Tqbw3vou3Y0xOspvuc+ky4Csa8YZxfNr9h0jteemRG654yhMMHTTsDej
bs9brDP5jIlsRV3V9CX65RWM9+ILaym+euePf1hbUBS+sG7cEq8WOs2Yv7dsanAkk9mK2OIXVTad
1qBQFu2onuOfUKibg18kVs2V6Mf/q7JhNCpy6xHYZvNGz9TJ6a20DUmwhoTdW+7hmPtWbUarQcD5
3NlIDIbPGk/Tr8IrXsi9YB+49m9II4vN8JfHYL+XVSat14fBG398O7ZYq25Lg/EQkEe7E5qfhiNO
riCc2P3Vqgn1dfs4grrCxTLElGQxL6gthBFsHjsN5adCLzFvaO77TRRZOWw9iUJgodu8uOXJPlgr
TeWFbx0lforsdu3WWM8tI7LCOi8KGaL0r0iLNOiCKiAZaj9GutDfco0xQWhq+iwao7nEpaRXgSkF
+LlhKu9t0Bkql3IjHdf2AVrbrS1Q2/avPnGcUdADzjSaN1SR+LDNVwOdsqk9ukOG3nMLa/MZFo8p
PczxSzy7MYPDdlgrBEpgig/FOl+Ox+1JkoVy3grJdGboF2PSgFA3II8N7OgkASMHAzdGyENLFip7
6QDsaMJ2gDhS1+11cNyvT0tiW9iZRX7XjjcQWJi6uN/unmDFux6D1zCMmGu/qn3SV9MyJaSVWH/a
yJIZRhXGYSvbFPvMxCht0zAMTgGjT+bYkgfgiXINBSZu+ulegLI48UrI5NIkbyBZ+rWFr7u4MnTN
12ciavm/DRs/w0+TPRQXz7JrnmrM/WEEa1dpYQFeGv78B/c4GsEjFR8IVfho9OziMo8JJPh0CJgD
xJYzTJIvgu+e0nappoCEyMS5lbIJ0Ez1OUDqV229If8TE2AgLrYdL5jdAa9mOXRW+jy2jIQkSQwf
qx/fnQ5WfKPvoAbGlrUHCAD9Ut3bjLaH/xNaTW40ACHJaN9c+RWlrR+MYqeUT01RM4evPxECEESZ
czEIs77r0oNq+7imHKxusP59JrYqenbeiHyWLwsgzFw3BXMH7yNbbwWFN+md4VBjz9ZYvuMgU/TT
+mSbuggB/VLIJAuv1IvMeWwkkEnzBDoStgsLiYknK59tEhtzBJF0FQenCTzAVXTqZdKSG28z+bla
TeQmuBssThfGqAeFK50Q/rJoynUfTlFb7CMYOFTL5uqSznprHYIgys4XsHThHzMWC3pWTVjbJpv2
Rl71n6GIXTkdnnMKVIFDcENhJ2C7uMcc7hYwj+ydu8VgYMXYdQCgnamXzJB9pqLvQIleoMa4HKuV
j1stefmRB4NK/I+mvCUTYG1MY8Gb9zlQjJQAb/Ar67UFaQYPiFTZu4m3LSvYLBefDMnrtUwT7bca
N6DeTPHz6gqtqFmnyFidt6BmxoU+JcTaeeE1yv94EYKzsQNIH7uDcI5B2vKXizqEXXjwQqCCQeDN
4GH852oLhO+C9miOptLpizyxh9UKIAIsSp784z38w6LHDdF5yScX2bWwqLHd94h4sFC6M5Ipszvs
Ql4UeuMMR6SDiuPYlKynEazQwj30z9aIFf2lqgX9gWjbE8EUmtwj7H2eDUm+2h8JT+Jl9dxLWDh7
COqHsfb2jPQI8P/+9Q2ys68nrriR2tMQqmB4RaiJCpLLempFiLEvVnC6fEOmwEu7lJ5JNb6sB7Rw
syxDZHppkx7uRI0Pnlg/GJVktHulcF6cfae9Nug/DZNZYf3EL+4TOijSv6uH8Lut8veUzG83vbAn
vsH1MGmew84vRAOJV3kiZSVGeml/CpFR8l8D/8fBXoAz6Kv9u4+QWKJfRk3IbwpNqow+/teBhULV
gJFedTFUghtCYtQrr5baGcadpZKa0HLk6agssbnN9yOsIW8u+Iw9ewcghYpSM27M8GnhQbv0kRRn
KQXv4cZpnYB3wq46lS4Y5qDiawhWw4sml7qoPm6SGyORyW5lbtiMFlu1YUtNK6ctf1tdz0dhcjBW
XdXCwGPVDnMFGqATSpYeFR1SyHLJpFU2N1+ks94rmKoFOuuwRUF5vVzYyWD9M0rT49TyTzH9T+5i
1nCMUz1hNBOkwqa7Wd5udMfzCW6qxYwiT7mw/PNyhSvHt+igPyDB8DOIAWmI9QuigVNgnG4bTM86
QYF/Q6I0tN0flAGhkntO/8URXjs2owHT5IalXqnvyqGHW9a9yk5ECZAUSbcPazAvSNJBIQNRqFWe
0JpJW8rTQCNS/Af2vsEC2DlmxY9WtwndhQXb/5osubFYDOdNdGfNiSEuBicpXA2/1HF9z3NQhBmk
ro1i+rI314XAlWUGqhFwZM9Q06Ljz/1FgLmLi69YKn2YGE7qYvTN1P6YVGzClsuR3Xu3k+CGFGTn
FJIP84Eb96eqEiCRzArJHFAB9gIKnr52FCQ7KOwuUjtO5fKqqR64DmzpGgAdgWtMD2fm+iMshyls
6hnldmectS0atGHgU/ch9kcYtKHnnsAGU0llP2nTnePjUJ4VuDOPLPmgJgwW20O54c4dhNSTk7Tx
26+evzm4YhcwKuapBpPqpIMD8ohnE8DaQL4A2kaj34qetYy5wXSaEjAxOak86uMwEjk9jbZAFXKg
vGKD4iEuU2Iv1uXcJwtJR4mUqTvoqb22+12wlZjsBCew+Y9pZ+gu+HR3ZCqh5w/J8S5NwmHp2Rri
gjZNsZS4VsKnWyxH0WEdFPbLlVv+6zbsgSdKTtOAXBMaTJkO4o6Qbw8WAhQI/MqsJx9Xlm7LPKhb
96j3Bk1TmWFkjTiCY5IpD1mY2pHIsbQ8YjRlQ8g3M3z/wrqdEUuCKS/ldpYgElR8eMlqysttlyeT
JkOIVKgg5iU/XryMZhyim6+hGDu/bKEol1m3bAPEPAAXBs9GHshvX2W70djB+P433ogk8bvq5JGr
SNcdRCzYQaCuzLXnqmsw3sLa373PjXqIsrSJh8pwHd+FXwX3h9W/AUMtBrCJyJBXJ5dHx0mlp9fX
LrVsVfO0ciLIKmjlhQuySpdWIz5YNKp4kO8iUMpH1P8yCcn73pIBU7W/sj3jDA2B9h1L7Xv3KrWf
YiIfOnfYnGgcrvkE77PswMWRcV5HRMen8UdqrqySkp0zQShdjJ6b1B+qp0eTlAlNAEo4Mh7FJ8Ng
bDhGWRIqiFRwGUAJzLp3qkLsj+FdG4VCRkmwtDFMpfUp/ulp8Ai/r/AKcVT8gUSQ7QvSxruMFkLk
I3ATZIddkwjUXcTWCFq1GtL8B6RdCg8ol1ymvRudYwSVfL7IApMdTjy126i3VRDjNL8dhRQUCpNm
fvlNEM0D56Is20nlPR4LYp3W2e+flbdCbziSqYZsDrOMV6XLmZMKTKLSkCu7gPG3yiMPC1/3dTjg
gWMdFlpNftcUfPUeUh7y8sBv3Fnlj0LjsUJv3RvdoTeZI7jjpKsmAOHNw0ODPU6jgXbzdzvbqwPr
S2Xkfgl9fdpqWLrR2xjSpanyZMDlmQyeiaDuAGeieAUxK6DDDb6wfTS2pBFq+DPGuBD2yt/2Gp5s
uH21mdjwcJFhzkpzfZG7cMWqqAj7afcd8mVPHGrATxspS/E9bgJoyOR5zUEO3MtBKLE8nQ8HaOUe
dR6MxvYBexOX0FDPdLEq9kJFepoSk+dj25zUx0Gyh7Ejmzmvu4m20E19Ua0owLw/UzNGwfSQp0Ft
gqT2u/J2eM8u/Uz0g0ptnWgvO1Rkebb8AubnhsMAHzeGSpJdIGIf48nBSHMo2CY21WPTxAlqm3/K
JVDkfMCl+r53f7AZ123RywCbt1/wqJxFLBulYYzugzD50bDHGweC9Jpe1HeUSYVnt8Yo4yBko7Jw
gwNsUbUDHK9qGOqZtxmOtRcfV+z5swCawYZiQ5e79yFOdbCjutkR5qbuiRzkJPv029Nmf4oLwf/K
khLACujKh42Cfo1YlXyzc+9bIUM3BtYkJWRnH9l7h9FyRpYEpXwQT95u15a494SHpoL9heHZkSoF
re1rFEcR/Nj4tk1TIIbwn0kmXrhwmfLV7ykDZGuBuc/prE4l5YCPZIDQoPqLGygbMamcDU40cKQ8
kqj4v8J/3oFBtjnKWIalvUL4Xg+1g8Hu+SbSE8QnUoop2DR7bj0T2+jK9LUqvw2HWBUBHANDRlC3
K4Wx1moGjKqx91n2nB1+VsdafAtooW57AOIf+9s4F8m67gWn5kMo1hiPaZPhtxRqaJvNV2aAzzGb
6evGPMaLET2J/YY3y/9ZBPU5/ZoGl+m7V2x8RbfoxifTBgcSWKbBSTQ9jHxjk0tL0QeNd6eaYQ1E
/Qw6ZtMHAw+OsiywJYh2PjXbkgBzRcNfbJ8MHQ7E53h4NV5cRkPoTWKQ/9vcBtQzQj/Xf0CfD+Ts
RvUONJso7VCEbib3i+SGuVUNMVexAKkkIfxj6gdGnK3gPX9J8D+DVXJ65cP82ghb120Y0n10cuHQ
T0QopisJKasUzS7ocJ9PH/OIvj3HsY6omIyPlseOH5wAsGFmyR9O2YZMx9ZO9mLaHI+FX+mf6yiC
0LeNB/Vwm0dZuZGHsZjenaUM0btyzHnXZMbCH//4Fk2VaPdAOSSGw4ZOTgmUPnT9A4NQrJEHD+Wu
JD8e3fWVZIh3nSnb4eD4S4zOUDDmYl4RwAKCQUalnXu4yOMTrUWOjPQkePstu+osKBT1ggmo5b2A
odCTZZUuDb8EBnPtl/kUBfvX9fvOEaKU17tuMWRSjf7cblCvYM5bFOeOdijJ/gXwozrHZHXqhnEX
pYlCBBwCkKNAqxF+3q33Loy5jHipD55RVsFmVW23+nFPFSpMpKdQ+UFCAzEXfOYpaHDEX1KBQKWM
uA0up204DtmmTRmMVC43QP06KwkgbbnhkgCxx9pFBWWqhPpEi/F8cBng5fT2sfk2tdYrmrFwEFKI
oOWOz/RU9St4Eu3heQA/M/JtFmt84w9IH6VrQRNlNsyt2oD/iUpxDWMrqAP2vLwWmbZZ37vsYwmR
M5bo2oVEzdmM5n6vWiTKE7PI+K+dXhJxLBjT6OK8eT6PEQD3P+nQ4FNNU93FChxxVC741zGsYalY
O+pZDul9nmbd1nx4HJJbVTRYgmpCEUjgO88IvfOcM+V0oUo0BlPazrx+LcR/WwxAauI0KYa/0M/t
7QNR3xGQJMpTk1YfBKpeLKXJ6p+l2wMwdsOL8LeRrA8kZQkNXPSfAxsoE/LeJlB8Uc0YQFWnhOwQ
ozetfF3Euf9QT5hQr9xw3KpLvzjnX8pVOhKs7IWpijA2bREWh9RpQKbYvWA8DH3ZVh2soGX/zqTT
29VV1zfmcpMQTcg8LoU/vLUsfXvfq/1AFJLcO+ORZpkPftVnAlNEAJtC63X8Bw+ScyaoNV6Fy68t
OuzNg8833VzXqb12X/9vrgQk/Rp2lSXJaDUkW5KKs+5ZO/QnNKmHDB4Ba2tG3cQitWe7dY/qVLVm
6pSpMjo4LQB54UzGh51FHDFr/AYD35Ic59NyZZzZsSQEpUotebJp/Xnd2Yh9rzYhE6wrvXw24qTH
kO1RbPK7wbeNHLQO42qPu644WTtc7koCKmgoy65joiDlr3q1V0yJ7Y1NGq1o0vcnvuWQ0TuTlWi8
jjD48FFaiQejQYic/O2jV9thGTxdaAoJFkCsKPal4SkIIXt6Z1YWyIxwA9t6MAzH+6xtCQoV7WdO
CAsqeJ56rWU5upZyx8XZT0tjZ2pW5SUC51cqvsKlfG3bNEo8n9AtnoVUrYCsOqsWBlBAtFQdVZ2z
Rsl6ADOlCCWG+4AK51DAeTUJ8sNQjN9q1htcpznivE4kWGhm67W8vYQdkHO4zvE7qnxPJDdtyIis
eOfgoP/2HK4CcYzKOik5U09WlTFK9ctNG+tg8dUSdA7gd5tAxBWoOWd1g3j72OWVo6uQcmAjTrB0
PibuvyQytvth+5n4Ip2gOhXUFhsexzTfAPjBaaItByl81tHqd8y8Eh9DEj7DEd0mPHDyewhtzTKE
9o6502n7Qsk4gfI04kfokdF1tzOXcIGebg2ZItgAE8ANJp3fUuFUKBpOJpCG4TeUQNAA7Dl4citl
4Yww9JOp/9eTMJ0Tmg4SqpWLDobutZVpZwXnawwyctcO5dKDxx0IPpG9hug37GdqTR5g+DAA9OkC
8CHIYw1pzw7XNHvPTUztGpE5LK+k3CTVtUkpATdzuozJNWkcZAX4q4eBUQOHigLRSkXLS+MpFk/H
ac6xNiVYMED6mRctESc2UD7xSsFQr7OybamrnHvZFxz7Ix3KifcP2vFPzsCKcMBZkF/3779rfBcv
9gJLYhB2lZYXD2qsNNydv0OVCAyJfUToZduWZKBicEdXSY4Ud8p+AQgat5BlR2j/LaD8xZV1J2ul
d16jvXn0g3FLODEUp89v0OLKf5cHOoOk7wbbGlanKjRd9UURl6Y7omAwSTaR52Os65wQ2TKa85Y2
L3gp3eqTBRtDuBTEA9ec+EZVzi3q2DJw5lRjTW97cRhRNEdBlxfNnd44O0a0QAzaQlt6/nDhdoEK
6vR7f/mWQ5A5KCIzqpE65TeE3lvAAuaKsYgdOZpx8A9f6FZHwR96+sHxBq0ScU/jwFxdnzaJ/eVp
oum0O2/RQs4rnSCBpQteRFq3sJ3VVJcNovFKrSWEi03UNovuvbfLeUZ+imsizRMSc7+vrfirkCy9
OQldCeTsfXGnMqKhdbt2X6UGevxEWNrnFEgI3J6/+y9ctDuvyOBD3WgJlw/q6ektF0blk8C4b8vY
kaNgwyytVyEZGLqzeaMBYHzuJRw4TGJ7Rr0EXuwI8uDe5xbh/lv3l3vg5m7disE94/evZ+l+OxxB
nAwDBmQaKxegzk/qt5jDo5Sqtq6DNOU8kX3y+8gL/dH5EmyTU14ypYL5CnuG2SZGfbSMHf7M/vKT
S7mW7foAFeD1Vl3dlLTHGsmzPDhx21BiKyUHGl5k2q++XdAFvCIXufy51eiNRTU6yN13lSJaq2T2
O5AmPNTZyD2+KsNVoZGOKDIOdvWPbePeu8xdt4vkw0nzIXPQREnuX9xGdPEjF4uqrxQpSkXbT2bY
Go11ohJTcCnyXgTKRjG/IguK45smluylZi8CDk4UVHq/K5H5FNy/oKNbUnr40JePwfKvN2QON2ZW
H4S6uZmhszbzDwvY2bcDcQ1x1xQmVthOghKjpFdjRp5G+bwdHGGs0p+72lRyCWAAn7VEjGM+DM0t
eig8bEM+cI1NoZeAnqsxbSuR4nJrwjx4p2tjpd/nCzdr21zs2jspS1+q9291rTTAd0wB0WSFcbEj
zpL7+ju77XwM0E61yzR6b0BeiKUZyHeOBhICZ0uzq2NnI6I4Hr8LNUMXbxoaL/VVeib/1wN575j2
VbhzjzAjl/UhQcSoTO5HXHE0RAJq1cd7dBGZEf9as9SceCRi+KRESYJQEP5wpWTsmMDaEBAvS8bs
pyVJD9WSnsYnFU7sAwnaGZBU3nyUkHbWSh4RR5MNNg1fpUHFfue7FG1+U0itrGYx0prMUvy/8FGf
kyo4aV9vkj29nzTHiQUU9x2HF8yxKrTD42KnEmUVqWtKvIN4ConaJHrm2PekHTKK1bKL/r8uZS06
AJIrkQvx0UpD7RLCHuADCcyXCMOv5gzUeo0iet8mA5UwFwSXcAXwF5W2ovyvrg/wQJQ/5iJT+eo0
IoioM/TsSS3D9QJd8ZRyLVDt52C5/aW8wutxHYjNDkddKYEla4PW1RJbUw/CWmIOUjaVPbR/mzBa
DnpG/Jh/kSOfrqsIKwbj8VyqBTMKdHjMwoV14mkpydgzG63Xtkds2vf5gb1uiIK1TcbMJKrzstLp
PvIMezkN38sW76+7mjcGjaN9bXu/cV6PI3b8zZT9CaS5OTRuNqsZsrWfoXM6f4FNEKI/iknAnH2s
4kACykSPZbB8uUBQ8vrYr3xGxQxKertepgdNcR/0tC5b3iK7SmBsaR+zRgW9/ryJ/GvOPAiz+ra9
xKAVtewsuhQAGaOLw/1IHc1W7E0JeNl7zS0QyVVC5DMtVngXUUuV7gIayuXgCZFFyOM65WF579fa
ptYQw4yi198eHgQ8+7MCpoGOw9IMPFtQdjXU8qmIwmBXtO/vfo/eVo3fEiZRvPvJCHXizPe4tCgh
rE9yO+Rzp/d4YEjIMwhFuy9YHX4pqDpjHoKD7ZICm1/x+fiET7GoqoADY0lXlsam36WWSmZlp68B
XCoJkCJVFeWEJVSjNn3bNgy1XucpuZTZufUglefUumNXbVpcJ8Oz17Bhf1Rb4jqi3y8KhVOYKXXC
7j+RX4OZEAzsljemwNOksP8/0FbAGDpzK6768Q38m382sWLaHfbC8tTSQC57sVcM9dL3rDW/rxws
H5AZDQ5DhL5r4uDrEeBNDOZuqikSSGi8R8gXNY0tLBJhKQLDElQXHYIZzvONL2hqyTmd+0PF0Roc
SxzFlz1hEWebD/He1QgozPRm7LmMKSDqr1mbf3K2oCTJWSBByqVIKFMdGzLtwxV5PF86Pr++X67l
0c2FMTQfY431QAqGCUL0qdVezpgU3XBtlTzzQwZip0B6882XMmO2ZUilm3J+pACTfWMkkCbK/aXH
e06NzQu6AJCgyiJ29f4qFM7mx1gRLw8/ABU9BC/ehuIZ8/5XuXQyVNkyD8nT1MG/sqKxfz4zwqrJ
Pjx3oN7sKYU3k3dl8gcpjVC2+hnwP8QFcnRD/fBiCno5/CcYiJwSY4jlG/UTPIcLCh+j3x9q1BzW
kkBwWLX3TS6dYmCjuMckgi/6UUW7Svz/KDDon/rtuIJkvuKNWnm5/BcmF2BiY4vddUvO7HH9iiXI
bCH3zU+GxQ+Ule+Y8EKzlvw0GzupeXfycW3r8a2UEfivpIX5kHeMxz1v6TOcGp5nn5QHoyPh3fDZ
8QxEJwp0GDms4WL8S60PuZZ8pwaNncD9bdDnQQ6jSszToj87qF5HbzBXygVZGWXJDfX3vM9va1Mv
5QttioJUL4ZRkf/fAa57D0Bi1nQfTJmJZA3mZxv2tsQk3DCxA+YJPUc5HrFBHVgGtasIVefF8Rxn
cZmrrwzDG7F/QGSHS946EoaD1Z/0OY70raOM/EWbV9hPlEgOE7z55tJEpkbX7kx6kC7GI6Rf7eQ0
DAX+lFKhIh/ejWVh6CvkFJQJmLeRhgVSde94cwlcpT5ncsTR9tfXwcKM/wK/AUoI169N8HLVzqZF
f92g1x6b9Z8MktWVODiHbzMza1BHNLKlJrACpKgtKGkd8vGYrfj2K9+047Z7h4Sj1wyS+c3XQQQJ
IOFrJ9mLPhBnRMosBIbTgLa00RemuyQPQ9bOy4mqWghYnpD2JQTOnivN87hCqonTU8/+hBj7b4bA
8n1rVkuMwLpvnAiigolSL0V0frJjQ64W+J6+ir0rhgr593umj44mL3iXBi8ks2hpRUZwDWWcEomv
YE4AwT/7KueFAYOcZVdxeQa0JMpFi9mcGbVTb7d1H3sR7sTlPttoX2mFKCUe7acpPU/jIwyvjseX
LZ0i214TnG2PDz/wSjCTylIlixG3J51VImg5Qn6Giqu3/mPM9z1I+FnODklbMJKj3rOpIjox0p1T
/apKvzcRrhmk4vxKLo9KRkrJFReATPs5kIxBpeDS8ms8TXYu509KD7dUTUPBzIcN4t9bvVfmA2Ra
d+Ey7dfrp7xisRnxQew1T1tDKKK3nftQ3enm75w/EKU4ktoLS4/y4qrTvV2G7s1xJfsf7J+JwUqL
aKLIVEC904u2IU/NaEpWqGi5181EeKZjwk9u3uTZQ4rCaeIKA4miH0ttxMpTBdBUq53allMLbf1Y
syieCtqDqaZZe6PKca4LUYo9EYfjn2U3bt8a9+TGyITGvsf+3zKmLqzM8qRb74wiA85dgx/f7wFG
MNqKpQDwp4xvbwPXVPfDNx5foQLdU/STBFjWRklirNKtfJKput5I9IIKZI3v1GFC1TiZnOMcd1FT
3wyB4fCdZnfBaFShjWWhq4Jh9AObZOOjswWBh7rtdcwCN97DFJYApkt4DlYsLjJ/dNkRKc64HOBr
wyKrB+AzmT9MQZomGtH9n+5CMMcjjQs0p3r2BRWxMEkS7p8hyrjjUplReNvaJpy9+Dl0+Mc5KaBy
ZNjdJcKDvqxfmfPVHDyFrmEbDkSrdzcO4POV5BOm1PdvhyzmeheMJZiJqqc6SafbRud04GVrCjf7
FoCQE5S0+gwHcf5YvB4WGQiE1rlPqBvkQQ4gqJ+sMiYnEqcP9/oAW+iErjzXLtC1PlTLWwGeRZsC
9aQYjRc/Yd88T0BFPuxPoB9Ep/DoOGUCOQ1UAawKM6Gw6LP/MygBwoA0qzRLWNsVM2QvxL52UOie
eYAoRjVL4gDKJpmbS3xM8q48yC0r2sSsr9A2sWV6vdbMCYPAOSrEqY0LcpXtNI6AEqosP0hvcyyb
5bgFc4lMnaJHXdCIdlogfjf1kWNkVZE7cbqifC4iFHg9upUMxsNw26PJx3s60t/+U7QTpCn7frQC
suy//x3WH3Qv/DSmwX/3XRlpDAMh2stRY6qMkG+leO3oTCi1mw932XTUEnzmbVKpwK+xreOhSQUO
hGjrg8wxqVAKlBzKa0N/KO6k5vA7Ihzs/ztfZvf5uu1raVmsAQgFpbEATDjbigU4PkgAX0pfd0FJ
P4sz6rOj5boCvTxwdn8YFvT+heq+DMpVOCDZLOjLzSEB4RPe+N4zQ9RalzQI+udwIvWA38C5fGk7
O+CQpFcQZFkTJy3QcBrJNoUC2ekPa5VR4qsUtMghvM+2EdODGE/JWwcf8FlDVN89tNHQHl0+8ixd
a7/Q+4PkpBAnHsiKYRvvLK6b8c9S1KMGFFjNB7nGayBFTI57KbBKMjOfjSvLBtzNbT13HXpxvP3N
1gbT/b1kCoow7UkxP3WIbu7LxyI/zec3rXZKub3VevydG7YoG0wuIdIn55JDMXP2bAMJkHyHmbtZ
XUxmdfSDUUxWi0+DjafEqD1bH8ECKUSAVnQWCKLtLNq000ONg9x4WuyeXLPL0487lpb6ieoVshkb
dYhbMBLdlf9aYps9zVs3BbCx2YJX0En5CnOV7ssaeZFSOTiawPEYtUlX0EdXL9K2cxnVcaQ04Pav
TI1am6U7Fp7jq107jggWzUhKqg0xKT0lM9zkVMP8htsuY7UwRUYP9lF1U5sCMcqm5L8HV0BwnSEq
IslQbbyT8GkVNhem1DCqX+/zSyNxofKLw/0Y5X5098BTWQNFrj9Aa3QyFjNLrCLIpcTda00CfHpp
PkQ1odW6sUOpg8VGe4Mrgegohhs58VNERjbuDsi8w+mPTkFeR+zZP2GTomFI0LhR3weWMFA52Myb
W8C0/x1KU7dh2dd9RwW4aywxQeQSBY421SM3VeuN/i4Nst1P1z+Qx6hlS74EP/0Eb/Yrd/TUZtMK
P/C8SqDyu8jR7JZY7rtpVDcdo83hzTKcP/QMM7oit6EDX4OTKCJ030l/N+o72Wd92KKyxEPYQRUI
BGzFUNLDht8wVtueLJYDRNwBKFtQ7LxKe+fOLgQSNePuiQlaK+enSqDcFSFTkkUsLf/JNHYYanLe
l2mMXakVmK78hgjfoJu4Io5C8H0ALMd6CktzaXZKnJxg93a4B8Os0DZz/v0NeKh/wSjREXuwmtl0
uTqQ+wsSPMhPopHbDa49y31oOEQamm9XufYXFGrDFkY6KottQCfKmF1ZylgbBOiuTR/WTTLy0Dhj
lJ4Gz7A8n8+X8RROP3JOgiNvPZni5XJusebDsZUNopLIf9Pn+ZIBwie9soUNVP+LQoM1UaYrKXJc
XFMW7h5Tjxww7PzsdDzhfVKYE5eKWmVJdMeUayBWpi/4mxlJqf96PBxTRLc3MD4nfK1CJ2mwtLTz
bEFI1TxktEUx0Sy0cjr1AolmgCBuCCg8V2slhb435tyJ2E2jjrbyanMYSleovf3cgX5zlyaeYQ5I
pcZhebO5pWyYJ5xikSc2oiomaPKME0VXHKj9NZdnHtPNuKdUUbIrRZJ2NxZyxFsk0MZo8M7OgYLL
fu3Jln7rw9lCsMaIgrAaxV0duOY63UZNSSgjWli3vHGWR1Pm1+kly8dmqmKjjN0prA1RFI8IE6H0
uPqlPnRKVhRO+mtlFNnuTo89yYqG3mwjx1u56su6+bbP57B3VZ9vdJQsqoUKg0HZq8ZYQaLeehEf
RQFZc1RyN8efazmLLHcUbhQvpXJINTISHdhp53v9h452nORdKAlBNAJ0t47BMfg9o3c/yMcC3McC
GxdNjXeXxCp5XaEo7uCnydiTgdcGUGMQhxmw6w0K2dqHgRNZuKR2MdFcAmG6x09oGxYFlZvafq7H
mVJwRAYNFv457eSGZUjbM931CnMWFr/l5FSvJyRBXPtbmCZv2CHBjG7tAB963DvlebWZN7ZiDdOH
j4nq2lnukpS+BhSLtRcfmDdLgncESlWnlUQ/Y/gZgRHtMGBQQbpSe/SZewfWkNb81cPlA9L1gwvI
RJb2Jt3tHkOii394yPibX6ePkiUH2ermFqokVxB0suFOcnFKJA8+NGZu0Kb03VogkMcFvKXXUlMr
nc89N197aN7/LQyZJb5NhwE34vWTGF6fUnKb+gro2Ybu3n740R6kv84u3xYkem8zbuGkFO99g60v
08sQXheq1LDimLYHfhI8BoRUZin6YQ4jEGhXU3o/kJmAJqe8Vj3i/H1veiPjSpPPBHDhQB5DcSSy
u/zsp1/XVbvWk6LNwSMZJno3XHjKltweAKUk2+8EdYS328LMyExwu33vm2Vdtut1cNxBns9YXYkI
QiKHdB1bu0c9V9Qn/ApKe8rjpcpfQeyYLn8MnMHG6Clvy+Lvc1pk0gYBhnp2vFM2OyB23ZTDhCxX
ujq5Emb/LsB5yIwo15Lu9QOBYQJ6N3+8VHUAp+r5ySCpS2SIzRcLKVzefzU5X+E+LQP1OfUyNc6+
bEdrQWCcqkdPhLf1kB25j21mL4LoEpiYtBI36qRVo49rW6SWo7nT8ywvvGSXDUCiCIH7PCKYvICH
vmCCQXDoLT/7NmFTxfuqPz/SaQWhmDA297MyDGCqH5DlQhq5JAXwObglCbPP3ItJ0YWDoDjlNRlr
4EUaQts//ZFFtvCuGkVtSGuKYvCCygai58dQ+X0kNJQhRfgB34guvtqlVJEO6mjoHbKVlJq280bm
HfWuBlcN8d1QJd/vSOTXiHVDHfvnxrfWyDmer25e+ESTvK+3V8xneRZ5gy8m9V/4mVJbSvb7AkjC
07llwzmzyLT/dtBavrMvZe8PEQ5PlANJiPtyEC9MWLB6+S3TrM8Fy0mCbO377MsRqDo5TgItai0f
VvZeAnWg4DzqD+HcLFZF7Sgk9dGFxQ3441XJtXrMwSK7BGHhZAMLU/xEA2nWELJEN4DU/B7cRd7+
8ETww/2fZlHdhZYTN4w2jeUFT3QJRbMiD7Seu2Q2NWuKZpsmACDIeZqrurIZr2FvsYuRSTs1gAzn
sFypz3zvcaVLgVobL5YN+LS8rt3qoTYyV15x4uyJUJ1GyC3scHHRqhG/nAXAN3nldK8icqfGhos5
PUzEmbtn2PcsYRj2Gz8BBsy+iZazg/gKCbs63Ku0+MC6SsJLDEP63vTu7aVBzDeKrDxuxu4Hk3sh
7ar6VAb3CL+a0MMYNXYSiDx38oO3U9mr5QletftKIIwFzYY/oi92VDHHsC1dK35EmmRJfbegFHyp
P2/nsD7w6UAKAGv+eBulKip8lqlDLtKQwQ0yhpJze6UU6utEwKAF+9ke5h015vIzyFJvRvByMVvH
aW15SXd4nNqP339Z7xsMYnpXgwHkdu9H2yu3OYakXihHXTGraN5G8OO/+y6uMIfWisyGqZSWwWzN
1cBIcV9gDGia7nDt5h2w+Q0EgLQpzV4bsvElVxUiRPW0M7LLi6CRE3d5LO2FQUDrW0UaIi++PLug
bUKB4DBliofsv0SilpLROVwh2vXlRAbehNOJoTvMMs5iSgGnxjwJA4bCzCgv0TT/TMgXgRo4HMln
X0LqHcmZZ6thWTNk5RaSbH+ABKC8+BKgIFn97Uh2f1xzkzHWlVDmQs/yh/8iRi1pqyPoboYy+D0m
7s7wtx4lfJmrl++KoO8eDx2mCOa1JynOibv8LCjM5desM0lKi0s0OZWmGVH2W8zjC/eLiMsOVvi4
WCen5Gfcdw3uXNPBqtkWL6MtfTqXDjYsAxyUi1LaLY6+oBq6ffPuzTx0Y7FwmqejePJYC7JgEvwF
iSynhGsvipxZ13giP7NAcVoQyPs53YnXA68fIn3gXQBKmwPys+geYMkaF8hwP9EDptJjrFxUjG7s
ATBPL1gLaNI/L7XNumb/mOVXoVDUbsnWbQbt5MS3uSqOAG3sDXQrEsJ7K9OfZjlq86MphaPRRT/9
9KssyfnGrfgZEb5nWUs/QbuheCPKLaqIScp5ZVZPN4T/HpbSFF6A/21B9GIoWyaGBq2zfqNlGqWD
HWwiQk+LRxaC2c9ngRpnYXUq6QGw899T8Qlfm2xxt8T8UtNX1YT4J37jRXHNBU5SiVfjUfib9Qg/
+eJ1Bm/9pt0ySF4OX0YubAJWgDYOBWF5zzCa1Wfl11PdxFU2MjnQ2cpaTM/i1ufekDORzppeEMSU
x7dkllJ6gml0oGZ4zhakNB7jicRtPcInZhqpF0RcFWg/4hwAZbHB7GCp4oCeGlJwr4d7DzCM0ADg
qnxkM56JcZjcb2iWy6L5gtlw1rDYWuD0CVtaBc9+U2rni/xLHqa+A7f8Hq/MQ/rdoAmOuxc/73Wq
PjcQNIpg+libn87aaaLI6i0BbMe1bX93+M+W3ZnpmKiD+4ve2xO9kUjpJgZFVeTHEfd/dsWMjuvu
ceSF8ALyEJVzGevMt5YeCpAAI835gslBtVF4JQqhzFLH03Ic1zGTV27Z5AeYjAiKBHW/6QvwRDdb
oJA8ovktvGt3w6oL2fY6uNZTWdYD2IM18DrotTdTGiw1j/mNTThZwv0Y3qjApgN6sevFAO1ervPd
SXnXtuNDifnIYCzRHaq27d6h2r0KR88GmUkRckDtmeqjfN9j75rdpZ4pH4+ANt5wcUPGsWamIo00
OfowXOJB1QxbVhkvaWGoXHHvyzNJg6dCclkgasR3S63maMKMZBaYcZyTnvsgbCdiXO+ryNKRS/WX
zcZGkzOuyVIAeBl2nJNZLVEetX3vd7ci0rgbjFJA6UNA5KhtM20lmzaoCrc7l690Vbx0DwF4DmOI
dKQzhYx40m0TLmxXypSeO9IV6vRfsHN4JGoh2Thapb/LdIHkrPNeo9wC2NcuT78s868fhTzNfYLJ
jlpblpHFCOT+PqTSlVeH3iqrTkEBTEVFHkog9VOFGAkZ9g4DTCCqMsOM3rAIw1B6evbx8/4c+rTi
DJGMcFvvvZffjJQoRCgpcXrD2A/JZdIfhgHYBgn6AbzFiTkye15Ms+4iHK1WRkvThhXQkGuxkrib
uorugT6ZpwivaaGm/fqmmHBTsN4SxwhymR4FWwuqc+vY7Oxc4IXmDlI7W481XZ7FDmr5HiOjJhSt
POrc5q4o6dOv6krt5jJIji07yL2hDCEu+KnL0q8aZ8UgycUYfUqyULY1bPi5YqLoK38to9bLOH5L
IY7SHM4NX2of0IxIo0pjlPfmoCCKi9M+piQsmc+lnltBqbK7M8eqm+lodQVjE9qGzizfighAUH8y
QxsiibQF/J86Gcc9lQvXcWdEJ2UtJiJjjRFJmQ8rVoxzL4+joj5CFvY/czAdJEbC82TVBwVQCQfh
zCt5bsoUzGhlvuVAgto906RDupe86cMI0JfEe5PG8DZA5FzZugSfKxiL2vPna8KPKhGU0BVMi2zq
jE6I3+upDP/x0Af4CIoC3PWfr5hp0J47Tk08rXbUj/ZZ/9E527A9BgGgefeSa2ss5BbndiooqXlI
HdqFkwnk1NH9WKY0Ilmru5TpQXvpAn/abLLMALOQ7dTZeqh3bzF7mPsvyf7cxn2RGw2S2ZI9uc46
adwvghyxDtrb5RqhYnBU70AXGdLWTCHJHvv4AhP/WFA2PDw+71r8EhpSY9RjMeXCHwHZB8jHc8Is
dJdj1+np0O/CzkDoknjgbe9pCryOnBwaaXZWpagtaogiLS+Rnc+S2U7Sb65iwlK5minTsX7LFiul
4NrA7SuXjfZrpkC09EWonI5X1vYJEsfkZVHZewGFjhyIrkT8i7folpxoLdMuMI0hNiy97v0LsolE
AtO7Gyqs7Ta6ii2lNT+hNTDXFq+Qt5yPV9N+zcOaoEXBKasUkn41GWMen9s8cTlka9WSa+MLV+Fb
ddvgRJ2tJEqG8/XZbdDJQUoUxYYTZSSQMy69YDvCcMBkrPdyHRwFgICG5WPY5tzi5Vuk086KLumR
rhUy8Hff4RrSOldljZQYdxKcNU510/qRzzMWfK8faE9t5OMhMJ6TlmOylx/5GE/ypvmzLFBLW/q3
dCxv12tdOoVu+aAkSWrhf47I1XzlrPVFHfFSmt69gobpXnfhcSyWFBxqyYHQai5oJ77wvkH2IApF
HlnYrO6rHPTXfyixGqtSoJ3dw7zv2L6aRXiwf9BNYimi0jTdN2S2fwDt0qJdrh/kAO2fG3xJd4zM
MEBR9gg9Yta35POGcfIC7tOWvhLzpMEhDmLWZsDuP/AV6JDw548HLae3qgZL5uEypA2AFZumCVRA
37JHn5B92FBpM3+VDnYG5cfrxvQZLYwcciD0JbXSd5NH8U00clxmuF1M11mBAyreMLznO+bCqvZw
uCUknrqihej+KbzXqDghWcHz4s35am/hBtVthAJkcvd28LLK4TCIMwQRj6zpotURuqA/QZiTYMz3
cM83YEndCxGBup+rAk3N7NM1C5Nd26AtkTLQ1xWU6KinyxIPuQzzxcrnR5tiZfrX0ZvGa3DiipIx
DfeITlAauPcnpFyBpuT/s+Xlq14LSpbSQDDmyd9CnCdfWWTTsOuRRU2lUcm10umRc3kSH8hijJSv
vGKLGrKp0Du6IrWfpY//giHzGwwKJ+557DNrQQLlB3557SH5udaKv6QjSG5EJlSORahfAcgnkeho
VwazoJfVdYi+PnZz/tqyRqwN5hEe5XswkCTpzuFTvEbLNY11T7MU4LRbsEsUcw1g3QECZ8jZQCJC
bjsANOnFl3zKUTsA//+ARpjjauR8G0tr3F8qn4oZoSiLUHOBIC2252pK63+z+fvPE8q87/7nBE1h
XrKSoZhVB1s2l2KQtkQl7VGKiNVSanNTp52JcslSAEEOSQL8AOn52Hzqv3HntrZ/F2OXgZ+QmHrr
QYUvos6wxldMjbR/SEeKB9Y/MdvWVMRSyWRjwOIImnuFrppTVXjCq4mhdyXSUADnFx5tcpENSCfN
Otukjar7udBcVOg33YPXq8Pd+LgUEDAouxqK5RaPZ11eCYmCboQXaSvA8IHOK+beVRF+1QJG7dj/
ny1crNpjSo7OHBWcqFI2s6FT0F6vP4r2+/aypwlmzGhkGu6TPp5yefaVVfFNGGcEtcGBXyTk1VmM
1W+nb8e9jnB8RAM98BFA3GwvyTG0N3liNMegGNPrdcet2adNrSf+st56RO6X+WqBDdrb31xJOWGB
PmdiMdAc0msXCVZ4zEFwfToBoijt7fz5E9pm/T0RjDCb97sFDK5cDBMy1AcyAj3l5c8ZIdzXr/02
Veuu74yA2FbbKX3gDY9PY1mpf7A+YGAzyhHsSkvJppJ2EAmaJ2k8LijH7qMa92dudXk61/JT5Vjc
r/ckviQMWkpcyGUlgA5FnenVq4tWMhb1WEFkqfyEPbECEt+R2URYGXzXt4+wk7PDc1VgTlh+3max
nOuM9pOXfwhP6yjLPI76hos0J4VSGC085kG/loszAzmQlb3frBh4kXL8Q56C9fjK+IwhiQPMsanh
pbNjD2C4Lapl1G6cXxrnEfBEY0aEgfoUpMi3TFGFbh/8/dDwdYY4ocKGScu6gOE1H1vVsovK+p2N
zOplKHvcANMWWT42XIe8kKhy7c8MzoJBR0o5khlMCqS4oiP6qkZO9DJAwoIl1eRjHpxa69bYO4gE
ttQCPXwEK+Z2hkPPlKlCmmFyb8m0NZTiJ+E6ppeyVw2cQrO2xbbav5erWPC8U7vmye3cDG86zSjQ
ErEzWbD0MgBtQHjwX508HQumPiReR3GrEYI2haEMPuIsqKjWJiTvRu6SBI3sAP/bOCJJPYnuMHj4
dFX7kzDIDZu+BQ12gO25Ri4zXfT6aBINOu9XnQ3mE8owQX50Om8f48uaxSARjRVCfcHFth5icXuj
tHIIqVb5ydG30CuHP/eFyhmjclzU9re0+dHnQ0F+EBOGAyguGqq9geYuaHrxoMqEeg/7ubQ4YPEl
u0IuIUu4K7OjL0pDKfJ21a6wO1KMI4Xz0l6ipwB/I3h0tcggTURKZ8Xekid74skOhT7ENLjFq83F
H+eHBV9S6BUFjhkVGTHa4BsaFqSI2ixjI7NKlhm2TXZZHA4Dk3KS/ALwy91t9ez9tPvuh+Vx0u8h
efgcBIgBgfETyexeWOW4zv/lFet02Y3YyzBh3KlwQ/vzr8bcOecT0Kjrsd+GlvAscVjXkGNSt+6b
mg237EI/dYcYJxMsjSFogzQzORP2pVLjYkf3qqhcXlOQ5mRykX12kkLmw6TxWGclIlFIT9nmqgjx
HohEuXg5424JsglESlRav1Io/8Sl9/xb4czoxOfsU37nC7b843kqYllK8htlgLo2N8l0EGmmdx7X
9ry9zVlKZ3R8f5x9WHbmLEmQS9EpvEWchKg5nIq5LhahL5m3OIrAC8+XlPgUon1NcEWeb9xlphAN
4SbEbvuTolAEn605VgtDtHk+eCmlqgHNfZeJXIEUt1x5n3UUGv1FgzwOEyDz1EpXMRAsLsRtPLlU
uLAe6bWcIURM4C681cbZuqphdRH8hKMxV3NcHYoXDlZiN0+Q9hUepIFddpGFWmEaZ1mHIlBc3UiW
H1fbk7fG+ehJOgpLhWVR200+5DgwXvopTgZ4yye3YlKy1RV44Z8VIB4GcsIBEzPbDb4c9cn/YFj2
wVbbn+1m9ZF5S+ENoQymxugAqwgjVpuUIrQozTPnY3I+XpOyjau/A4p/yEFksGd4QDk5TsIE8+Cu
6FSxQpwtzqGCbUKK5DKu8lIIMmbv6/HRJd2fItCe57rNZQzOaCEvlKrAeOM6tHXJN7mb3qVIRag8
fzyDs8ucNlc8lZ+85b4gBzy00lgDtDbKGogv9eG2q2lZhvDZ+yxaPs8whXxS1MMP1UccC+Eco71K
iqfEfXo05B/0jnOKZj4g1eds9ItuDWqJRhvqjS0kMZ9S7otBpMHE/x/0hwpr9g2RkMNuvICoItg3
Gn4tg+wVQ8NKzG9d9wYkVIhz28A5VmV++6gLbbA9Ev5dK9/V9Q7LXxJ0veoPijQ0bCcdZ9uYqzOL
PW+mvKdkygimtb0h8D2n5kYfx+7d1OJz8WG2gEgxCZCw7GQB/55zToHzmkKaLJyvC/8PXTzw/Cgq
g+I0LfuzTc5VQt+R2MC7PVRLgvTtpr+K4RcLNKx5wJXRnfy71kjK9UktGjGqVKebtji7CXi0wq7k
x7nwSajLE8NgqgjtJUYE/rELnQ+8ecgI5+Uy5Cax0nZuqhdWe+bR2vKvlrmv4THtpyy79Zcb1WKn
rGl3V9ZNVURqHEDpIwVplu1S9rWwmoBXv68n1evjpikugK9Lb7n1pXAOkau0xY03GqrZvn3ntMsR
neeanF5sHmXhE0bWp/bd5Kl6PFbGQCmymPQJtOt2pgiBj+c2F2MnAi5pXlofYOSGAo5L+XSr7q+b
vsXhjKGC0lt1HwZHcgmoUsk5ZskMi/ym6okNXR2eZcypg/RAwNin477rxIGq+agkZKYk8ieQBwki
0T0C08+8eFbs52eq7i/u4BVVkczGVgY6wDqxWkIIa4n0HmZe9pdK7CGcf3RXvONxJ8XM0cXCUMpM
7gOEmZAsYJ3gcNanXDwpWDrobTcIfWWPCwLBQDK8kGhEgPGfuoLe+9TeTqw6uMxjrVCUtcOnDELr
cwYVfFc1g5E7fEgjiS7I5sbdJg5gJQLg6uuGHCYYI4LKqy0egGN3w9QLrphKTh80WbIvevZl8npb
ZdRU2f2aZwUk3KIKDgED9J5YB+LgcMVZNPwzkVav7nTrxgZX6Xaec371pPAwB4BYRILuIH7QBOkI
eWXPIfTi0PLEYhTLFR9WPdatWozGWXm9tANVby3Wwa8J35W2trHDCARx44sFl36QEPlVTElvsDRs
ctzFhafFGnstK/N2Js3r54IjfIDFzSAniv3PQckn1Mf47zrCPx7e5GaZLZrDEX/Mt9rQlKA66Zjv
gQskZjITYkmF/3uHlfCbYgah1p3Tq+jdn5Uz4zOhn5WGkLioQQi7JernS/6x1kCykiRHFt+s8OtZ
WLyhpyfYpiDXegqA3HGj3UMgTeuRd/JF+buWsHv3KffotTS7brVvwC44U5XvnoTUFVfcpwTtC5KO
Rv+0PM5IPL+xOygdrK/vOKoChLVeMjrjKrnm441ph5S0Ut0EUFSm8/nuYLyBzatov4ixN+gYYseI
qpdUOyGpxkoH27TLWobwwyAZ4x7uSATjWaC6lybwTn6/hgeJLPNetLZd49eK3gwR49HbTlz+Eabq
2hErFIYwm1LB7c3zjWNGkvEWnG9A8uzsQqNKCXZTCaEukBNuWstMHC3E49E3Mkn/OxSNDIwxB3cP
2ksWF7L2D1cR39yv4tk7o8CxwLmGRVZp2ChBoWGcRtWoh+316WZehWpTOrRjqVXCv50WYo5v+FzX
pKicql5P9FbvCC1l9NIZvVVlXwe5mrtD85YyGM4NGAig9Bb+oVg9mjQLwKjR0CmQnWEJpsC4WpCS
ZY3SMbou+cvCSBP0IBmw3bW7CFzWjqONttjuaEmATHbxxN2OVGdnwUST3yd4qugi4p4Q32K7EEMp
FDFXSbcjvifl6IOI9LW1pArG6VKdxhr6k23VkvLKljsc1IOC8t8CeaQ5tjPQbOdJS6TUfzcnwtAS
DiLcOxR6FIAA7kbM0kYEWa7Y8jXB6MMnqIGVrxlSoPT00wmlSFpyZMYUutLMowLiuF3Hsq+klvCm
x0sMK5yUHkqTod2LGIdMB4HF1RwRkQfy0u+WZpTZmosL8V+AuzzJGL+GBb66kkiNd5kcDG/m0+6B
YwYyUznWZUGTHYL02e1hfbrUiQtz4qJiAjVLO+JEE9SPwmJNvU4hDckIXyGgEjI2LSDsrlJ4WSlh
zhrnPnu1o6NdUkOIm3RCa047x4kIgXbL5qk1ygd5zAg77VXyMdYijCnGoBPkyCAXh5PSmd+aghH/
tjJHVr3nByuadz5ebLg4BRivMl931kg0TIiDLW2ZIdW+BpBpRUjBxyVkWqMjuAk+hPBE3gN0AYG1
7WSNmMVbFeZMEN/f6OKfmyB9Nskye9IuKGR80rD3SuRY2hzirwPLq+jtg+vwbbr2QoULVaK7jadW
W6zS3XhBW8PUkg+PJ8MDQUfA3Y8zEN6MBld8CcusKt12vXj+/X3yEBGpoEavTNmcB2nEEUKhHMii
EooRHIhaQKEe02m3pqhYMpk/4c0sFtdVAyf4PacCWiyiG0mVWmTtmz6C1VK1IvrrIdcaCbLcQqYU
m681yNh183Pg2MEBvnJE3JkwQtmaW/IIp+nfzSC6sfUGRQubvVQ1DXYbXNM/kR3yUtrgVf07cNCf
mQ69lkNiJPMgYlchcEd8PJ/YOVBWaxMQlF9cEgLeSd06U6Jlx2xpTwgUcxeARnrRiLuwDZeTqUxS
qivcFqel04ZI9YMTP4uixFRzOGOONFn6qbTF/x9mmLP3jQakNwW5zSV1lo3JRPuy4yOhNxWAKcVD
k11GVk28ufKf9ptmDQtBBY8YKnDRF4DcfccJk6wYb5bRdR6oX/9BZFBA8rW4eeaijVzzE7dVfeqx
3c6iowDL9vHqMc2SSCBuUIaqG/7tGBNPDJy3LJN4rvjwAiqR785k/R62VSThaWOEP3qLLIvCxOgv
cpw7NYqClWDu/c4x1443EcxXC8yPehSWPzfGxoMc4LnhCkdtuFCec46kk5QBfoHSVkxewC95/xOR
E4NaFWh9dR13QVdWDjt5KyYOxhx7qGTW9fUOGh/TRJc6lkaizd9E3vRt78/Bgipfvv5bNAVEK32x
ODXDhhmnAN+2Xu7xbB54mJLtuUDIO6WgbO0qFJN3bWIrrC1QMBy5jaheDTIlLktyfdAF5CkCtCCk
UiVXEJArc70Yuq6vtdWnvfWgR67MkuBebPw4nComWgV/OltZG5xBSchM9iiPvtN6yXm6WKL4/8gr
oTZxyzmVrQfoEudfS2F8eJc60iUBBzmaROhj4dc4QH2mASJRlwUEzZoMcynbf0HQ8tWJP3qpT9mX
vYddoue4oOay0+qiduE02HA3NmwXpfvhZoHjKidgRCRmbXcAFUYOjdaC1ALbHTmUzj++AIP1dFZT
0XLas/35GfRSHqHQBvpRiv7TYMtox+dsuj59/9ps09iCR5xgUAbCHAnHF4bdcVdieymaAo9tpgQO
hYJdsMEFk8YNFMmvb2GXasQkVHAkReNtQ/o6FioPVtkI7D8XGiMhO+n2O2glD3dJftKftWxaDtwK
FJr0SrC5X5oHDG3QjFPiehTMlQlmo9bagLEeHPddcEZsJb2MySTZK52UfpgC2o6LxfRRNRDm43wx
N+3e/dDhs42dlpVS6ja12cTWCU8JZEpzhXr8GE7v8xEsO8TTB4UgXiSW85Ru2PJJp3nZdyHKTr1y
PpcKsJBWT2VXpeHLI9XF48gTdADN3VlurGL6hf6dGq3mA/R4aeiaPDA/OQtN05gN/Uzp0lIVxAk8
KSREAXdJsWVQ1V64bgdPu598lpLav71haRC0qYUesgiD1HZVK5M1tZm4lbf1r6tQwowGGsLt98Es
CbLGCEN9M0XTDEEnPLHy4+yAThYuTo1/4EvqTv6DAqAhMtjC9gVWOimbxKlqpZunUo/ENCths7Pu
p14yEEmP9uwwPKimC8laJbCvW64RPcWTbs1D9n8ezLLDTvR1tmqdq+3K97nEVhaV6qMQNcOYAlV2
krGsQOCwv68Igm+aow3ozaLjS6DmNNoxhfwCKvxRFoG3nMSi6FaVWizGihtA70FpMZ1Nm9YW1JhM
bVTL0FpD1FCTgIQINBk9ORqrNNnKBWBWA9vao3KKfp08c6ZcztS/EtAE++etBcWzONvwpav7u5WK
mCes0QTeF9iXoh5xM6MY2f1iHFNvLjKt49ANzeEy8V9vrdYGp7/u4jeRsaBUg2iRQdJ6XKLib6tW
mxMJZmobY8b0Nf+ZeoVbkdRnSvA2PPaong8csuW86LtMKxKUjn61BAdIjIarFvlQhyl2OTPt8jQo
aud4B/+NGkxIzhLevS9VbYYlXNs259VdAZbNiIRZm0dB6wKuBV8LLcFpQON5dYYaMsjEhgCf5KzM
wiuZwiCOB+sm/+W9nZEOWDlbEk3GtMn9GttCgnQChUJA7pVL/OR87StuIOJCo/QW+0DH4gKVEYyO
al3I3cj/FBJn7asuemMLqmazmoAog9V14NLCnPeX7LYzPjzTUynlcs6KK3Yn8IOfOQcwfMGKajxZ
6X3nZ0byLvGKsZGB0j5IQkBn8a+RS7dtdp1NCEWJjgl/7yhac106loPAxQDAvX7ZbxrjhNdj8bEM
B96mvRJCG/Qqnc2PTHIFKm+D38YLBqIgOIDzs8PldGSwmWQRBOVWvgmeKuROH3rpd4bC39kKhqop
Cp1CaYKOzFuek/EILJuAhQexfyx4tKvyknnmfy823wxTMuuWpDo+qK5JhnCB7LDuE5JRWZxW3fEd
IF+xoFgMheZTnVxAt+UOcywRZCZCBoPHa64+nGuSbyjbl3QaiEEV+hpT4l8Q3a6GoXlgwS4ITBXU
25VF9tBt+IYP0CsPMrSlYtvZ+r2+69StTHJnRZLxx/cEFxt26h7uHpZt18fyV0zGasQwvGKIksi8
adGy+uZUOsYz/ozU8eYjr34yUjUEIwOihMEZE/e4zLhqY7DTAE707klair2zvweIkcEJoWeELQHV
bp4WYvjLMSf+qJNoV3rvN2Pzkcr7El98jIyLrJuyrXFCZJB2AfbWGIevl7spKJ2HbOPRwhiGDXzE
1QP13ztQcovnZamFY0ADOFHPNdjgCALmiuCdX/64Bx1ecGR0PohOF6Yv0ciQHIPxJe6t37vGgSAJ
+hEdPjXmJinXPiwosgSlDYlr/XAYFmD9KYnDH5Ujor95QRHGhp8EATw3QLU4+O1w2JD6Zf1GQ00S
0eiRae32cqD7V539kErpmx4N09qjpVNDw6PpeLpQvNd67XTLun1P8ZLAUU5QMMzLKZeuPYCzO5Hd
2l6tg35cM3u98CdX+lzcxFsyDPERd5Y+6nYG3KCcBKUZ8xbzdLilAbCG83xqrr+IX4+plYKHVZrX
IKMnb/Z8+QW7wFCiWcgyOS8Xe+/Ynmnm3KUSqgxDBjaVWmzDr85UCVM9zGdq6OytujNdQWsuKmh/
WkV7iHd+BQ1QWRBPNK67SlBAN6MIpInD1lLg1X8CIDrj3J+uZId3D82YVdcFGaGAfyNiNXHrJ45B
6DdQFGiTxXcpIbxo20cgg+b0+EniwOcUyLa5kGvMz/7Y+Cz31rrkpH7757Qfsgob9iYjD3Tcg+Zx
M/ulW6H/gsUW/mLDbbVR+ops6tpRk2U9V9vNaNERfJyqygbDKfTfLzxi82juSznSqZOg5sqvKZft
TQUwls1YadtCZksx9uHxQ+C5AT2AQ8FLrxRwrwnXeCWebVOJOLp+78GlzXSKiiTNkcI9QwtS+Lmn
SJahSAobDZXD3QDHG04iex3ryeibyDR7Kd+RcnAeeQ6FhgVoqX6bS2oRx7KOhldNgJu8x75bvrDL
bv1erzp6PEGqEBUdfkSxXnryt319V3NTRpjPoCRDpuKICJ19tCFCJg1Zv/nKJyezOXt+bOe0sP8y
lm8TAfaTdh5JEeAFDQ+shzoD9hapc8aG85Rj6ZJk44E1QU8vLGiZ+7afBeqUBIAwhF2ClenehrE5
Rj4dqlPBbDh0iu2Ig+Zqt4nr8P+Fh0jMIm93GEoO0lMV56ltE2vaoctdSiGjIoh4b/cxt5KipniK
jcMsEcCea33lQNRK+69eTP8T14kZVvD2cd3dBkgnasEfk6fOjm88cmOTzv1IN8t4/TkfCzI3bc4e
pbIfMtY/p+C0s3uCw3x5mMjvW5ubglHkwVN293kYtjRsX63NmIdOqPmOniu5v0H4SvKekaqQxIbp
jnHGLRthho4eLPnPN2cdDJQOJtSKNbayqoGo9l9PVar3VIlGiUBMjqqsEeCrNo0n8W3eAiv3/X6j
iP1WmB7mCTax2cNfSqU3Crfb10SSpiQgb/0likQzoILjA5KxtY5bFY4ntDEgMt9Ab4pZQ6Q1q84D
3oKqeRBHdWaAOHmlHu0ZEwRMufYrEPZdSr5HqVDuA6JilpK2uYnjvxus7psGh1HAiwZmNe56NqJl
wUE5X3U2Y/BTJSCIkTOy4goYLq3kiydbadwISZQEQqO8W+j+pUIUrcVAqwCr0ablrqQAIJUjXJKB
0QSMdlyrKP1ch+ViNcFMePk/7kgnWtXAoT9plLTAKg/5joTz8tWr8kSmma3hpLKYwt8ZQXCIxKFu
6NKA1lv6MuZCNommlvmaAJQPGn07jbVvTxkLtPeAw+bNilH2UjmeRHJSdp+3BiHRt0qQ3cjsaTy8
T3IKQm+l8/zgfD2MIzlqhOUf97GtneoSVn7MWiLOUKfZ2Zr9kyZviastK4HbVrBPSMnuhjdPsWH8
rxi4wa1UX8sfK4h6KfLRFHDdhqFFXSKv/cizxHwNDNhO0kMb8I1Vwp1ZJVsolJU/2kWTkQptLGQB
CngXZvsFDd0ULkl5G0qRnpdYO0RyjjpLIkrcgTeVt0jn2v9Z7wtbF1X2//ZLXNZEEpnUDHdYjLAP
Onhp+1DNH2h6tjnkDvrP2AoUnuSlYoTO3Qd+dKbi63V097B0aAfYMIl0m+xRhr+FLgmxJ+Z1aWDY
KhOCHwNIiQAvnhP/kRAzgcRWNAQbpK8a1g4RpF+F7fDbWCc+nyBlVB2AAxSDV2y7CC1sH3tE/Gm3
hbANFJyxs0T2cxq9tI5NDPrqNfFHFa+vQpo3nJTZVXiXcypb6n9M4iD6shfQdAehDb+ZsxHTdFPv
mfgTB+rzjo2xJ8JxqCyhCKt0FDn1CSceYxo6f1xLr1ECBKqMtLAeJnCIwyBOXjkKmpw1H2q/ePzJ
fI8onEG0JpmI8C9pOpLh7lF5zq1vng4ds2/7cRsmP4N9uWy9ObPff59a46mI6Tk2F7MRswRbwwee
VJsPqBRqfXPPZW3gmWJwS9/ufeGZkr5WKUKDm/RcS5gpWY6OfF0SpHvBbZ9/z2/Qu3RZd/H7k6tS
b5rfnNeMRx641mBUWrD0YQkaboTP5cIe+NB0RRpDI24wzcnbOiu75oDw4BKXYtyOhxYhdSkIpSaV
VEdzBjAAtTzk3enVA2VkSBSD6CRqhSipikViXTgIE9tjHZ+ucK4LBPvyxDOhrDrJW1teDbnhfwXj
8y7moohb5hPeC+9o2awF/LVF8Wiyyz+jMfyvjzXkF8fOLmFQAdPhaYdAlVdyTxZMvO0u+IBrcBjS
R4y+Uyj1p0Hc73SNH7J2i5hqrOOaCvZtXwFupjbDl8O6FyGpElgrpchgBzlxX5WDFSyHGw8nmSYl
ireHNAOaj8ItmFnKTFA2sP4QRvRU2s+ebXpfulpS5oS3z4h5xPQs0/++GbwOZOdq6ML1iyCWYe5Z
3ddJYxukt84kAFKeUrmtKSPoYtPyhcuUipMq6T8IOfU0e3qOfwDzBIT6n43USsFuwTqJ367UdH8E
H6cC9QCERp4cfRCffgjZ8v8wzfXZ6k7xaNqhCFj/uexLFry/31RQTnvUAaIQ/Gl3TZ7rlg0xn3ta
fWQe1e+f56XEIandALAHguYVKpTzZg2Gi5GFvCeD9yeqRlL7haLugPqZryFTnDz5gaMPggaqU6Ke
HJAz2/5nbaMthMf5gpZpc7WKkqV1U/w6oxRodonQ2tXCQ8SAWsw7tEBZbrCi0aNRNQLiWX47YhM/
M99D03lgVNCXRwVXj89SbtKOR8gq5k+nZG4F6kXBbUlQYqun10ZU8ZgUb61yIj+me/iQC5m+B2+f
YE26xcnlI9zcmt1zuahX8BL9lldKpilU/IUADRGWrk12OMSkisCgpA225SrTGMlbJtRgRPhw2wRs
Qcpt8icR0zK7Hzjfjf88TCsGb+W2WeyhoZksGEjio2KVBHGqm0vpywQBOcSdj210CzPm7C56YNw9
x6A1TwIfJCAWkIrfpHwvSrylf+gOcR4C+xhc8E6bR3LL5Rnqo/GtUKZh1PyzI8IJyXccZN1GBUC/
jd5x5yY/bEhm9kotUOMd7S4fh/TT1OFjO049MOi1ffuexb8YJwUXv2hpLfvmHkD3Qi6/2xrxReOT
JZR7YN7hQ7Y4aSCnInyozqof95W/l6iWOBiLg3Xe0t03L6VSfcvuW6T7xNATTEec2coTtc3NXgbW
jJnKu/uzU0bcqHwPxynDLz9SJMTZSGjSMSiWfHQG3TL86J+OAi1eDtiQ2vHK/QqN5gSpVJ3sslbW
EKDSwl3INVpVSb0HoQUml7zr1PR0tGzz47bHNl1gf6vbZuIPjq9Tz9LhlaJtBB2SWY9sF5WPncTw
9m9GkPjk7OBZyeC2PNSUp5PgeHgF8JpDYuixHui60Ul/7vcQRGAu8qkIUwZW71tfVALEC7N2b9kG
0sTzY19TVkNx7pWzxco7AfPSGPuYHOf26OdwOdK6GK5CqGh/bBTTNBU+aVAvrsMTXUDA6tcyx5vY
OF5awGgUUfTRKWFd4DsrOc7ablmudWRo+DG5G1XDnVoiaGMIPt6zoe2W+LVd29dp6dbvd7Q6gnmd
TJcIv6Ktpmrx+AxGjO5IjSf/G+JAts6pUwpjmJUhszRr67sOCwWPjEbNbktS2Tgwwj1tnYpF79J+
lipE7cLfovcX6qMRVcNXFKH26KeSGyEpld9BSEfZaOW5RkSrWcGo/sddk3NFRD5G7suZP1kGG+LX
pNfaiUIgWdBIldI//CRIX6FqjzW5BZZ48bodaJG94IeTknxT+H0kWHLaJEIHoFy12XaEWGnxnr6T
SYjonyA84TBiPUbvG11qWeJVJQn5DjMTksJqmpAPMNd04+lp9QIHKbsuMqI/HdPCaIkXcxdmyoFD
lUQwj7NExRcfFeLd2dvl8Id0zzR751rmj+zjOctaX+CvOGix+AmR3T1k9OjbDKam/u+dNAJjjPPx
Nnq4/GbFtlSf5fEVAAY/vOr/mYSJsPvt/im7+pZUfKuP7Zd76Cu54Jr8bfPs+org6hYo6pglrP2S
PzrH/LYYvDH2XRXaXoNwNb7TcAfIULnbYYcbaQbLCwqrZhFmGnRRPXTxnYQChCqzoI7vsgMMM1nG
PhUi+zivekCBuPVHcz8nEGvO4dzn+h9CLvsE5MliY7dpyKju6ShrjX8doqoS83POAJPnu7l/qTaa
7LqU31f4e0HsdMbIm+8FZJ/I+Ydygh00rNLwP1xnKetIR0nrEWgfCLrJXnHRETVnK9LrXOpeucjW
5Q2yupLRznZ2GkPTnwCDnJtkf7Zv5imUvv9osxFf1rPPqFGJkMNeYmp52qUDfbKXdl2MamU2fcAo
xJv9WDTaATP/97BdZahptHopHSQRJBNaXOYRf6hemyUKRColrmOBzH6Niot3gdy/lhZNL6Bg1/QH
xs62eZT/o/w7pWIab6jf585uuCoSz1zTQL4VDbgTSRAIU0TpmesPYCYqXsSzJ6zeKBWScSMD+4sF
8b+99OH0GDu6cKdj5mYj5jFE/IJNb6MG1/7+0tMtbs+1iIOGex4PW01johzN+CL4jOE87EwLOn+Y
/AYUIH8yVxIac2h1zFk37MQqgv5/knQoM2RCCMiR/M0gpVbyZFTo5dX5HP9hahnnBUhw4uRR/0GN
GVJV3OBIxL1jnuSyqI8O/HSZXDjjJiSU8MGnAjtHldO6GzpoTGVyHk4kGzXbrQQ0sO9EkK1MFCJZ
M+40P0VEVHKCyeNZa85MeBVuAiUZwciG8gq3QQxRTZydCfMhQJyLo0eQIEPfG1otU3NnKTBeZgXs
ZLDVapiaPnh8dW4X7+I3U7LuviAVFN6Y3XO3oGJIMWS6t7J0P1ZJADnXvSCz3HwkSXsih8F5wuSv
Y1p5eA9EkKL6l+p8US/0qB6ik2vULuNS53tRY4JDKDt30y7S5fch9v0W8oLWNen6Ms/siItMqrIe
A4/u44pF9liouE4svbF3l/FT8uLz9g/AaHOvHRynDxWXdfr9hm/tk/2udsITSr0YMdgSlzg+Nn5r
eY8B96qa59ctb+g2lE8Tl/AD5FLqlyde3hGkCoiZvWFMHvlV06HlV4HiPkzQdGAHGr3b22Gsnv+o
jQW9WmUHcJZrBVZDDPLwxdDdIm+/mWwDqwTG6+PmMMBKXIDBPB34NIhgVHuU8iw4Fgxt7kEpGo54
cM43ceWomKEz+yBeUeiQOlodz2wkYELK9anEAzvVHjZwIHYMvIj0bNzfWylyRh5c+A63uTzsSV3k
GxsNMKHBR1DQTYg/DXdtQLHwC7KJRLOTvPB16PLn2P+tD068W4rSgq/K+e72THb2Cql0JET6ODus
jwGkJVpQfpgh6WLml83qkE0XfP3abfsULc61F0QUkjBcVxmfYbqv+abeWs3cCGPMMNMm3Bgv2Twt
IVkiR4+g7a46EBOrFaq0PiabPGEM6nX6j2gfEaCNVZR4i9wCuTioNRngt7j2LRtPWrXUFv+3ZEYS
/XP38S46IU8jWOy/PVOGYjJo+FzlBuhbRB1IC3HLPxgfM6c3N+H7uRzLGw8A3G6lkmFcl3TKZ2Xc
c6hlhWNitHth2sm04Heze5VxrPwrtnblGwJETlIaFPnCXXS5IJzP8imtTMKXbTetQ+4lo7mIdcQK
YfspxTsSdR1uSYvPiPB19T1gMHw+DHZ1AkWjfPlUM4EEXJhd+LlcSiyZqN5e0oYNqXEisJzCa8bL
tXvZZd+q1NfEgZMVPfgyThNz2ncps4q8keeDcvwGsVCxfhDoaXDwWxdTwBmTW2Oi9YJIgsMDoJla
Cd6aDnsIaP4M8hsag9rwCJKu3J2LXe85/FhQzAiFhUiyh3r7/mEbeshQRjgko5mmpWUXl4Sx16VW
FwqG8e9/NA5DrWki1XqDj/Cw1X8TGQuhl2fZal9wPx5JDCIojCewg3EImqF5gUiK45p97InIscTo
8EthtH5gwLTbdTsF2irxySW2wUL5fVYqXPvf/fLihkI9YCuJep/X/LKyNCAWB78vDNsZl1qimUJ4
nzoEG7OREqTckoFAz4GMOpSo9Tqze30wsXFlxtp6dJWdDluXv2NIVpoFj02L8ppSlOf06aenbJzc
8r7WmiTowFa80DbMil2fEcDoEUonUGap9altvSqk61pLNoXhlhnULbM/yhSCSyDSdjUZ26qZQs5f
MjBrKAq+xvqqeCrzEcG4Jikta08SXs6zil65WJbJOfoYeC9jeBn8mLkumoxeeXPBYuTj+G5HVW0d
rQXxWo36oNFk95hOPt7FTDu4zqaWEq1IHGXuV7GQZzHBJu1nvbg0Vj3yIeLJgG7qaMG68BxkkR0M
PnBlVP6wLqysA2iiUTtNwuROb0ENvOu+W8eOJPTnITySjHfwLTh8aqNesZa6/ooH2QlyWv9ZTHqb
R1EgGkVrNGbBRzcfU1VHB9Fa119egq9pXBgnumt1t7NiO+64Qd6U/tli4AWl25lp+TaxHoIXhl2a
933lkqkCROiqrVtAdnjufQ9fIiMDKEZ34MbRHERhaa3Ld8YqnwNKQ29PwWxgehKlvWdo0FSN12je
/NaXveMQe0ACyps6jfZrkCJ08iZaadexDTdft2cTgm8s4agdUs/h4mULTRAQl1Zq44gSPFAZmNVa
qOw3FByFdg/JmSbLUxT3D1eiDX89QVRLaTeaHYAZHnXDUE1X1NZb7Qb5A+l367swUJhDSXFQD3m7
cb+wd8AXXZXCYBNdnKW5YKj3IAvnV3luka2wQFUaIzkppQExPzzyMztmkSjOzA++6ftT9vT6xKMj
YjRg6j3x520HIU4Ne/ju89tIqCKF5iKFZARdrlg76YMzvWBrwR82ew5kpPLK91dgf53Ei1m4wjI1
brj4I0oGR/5qtQ7Rytkxhilkmy/8TyxKixHpf/2cT3jxM2lb1Ke1LkfFizqw+E4RpkjPj1a6uC7X
YxAuKtT3MTmhqB0ZPnfPQTybjzI6LQ2Icusng7hvP/wBrUGAEUVV/ieJ7oRDKgKmOEqbka5g7G8C
EJxK9ipRPUELXJqu0FTi/+1kY2u2nR08Y+tTERrWWlQXXa50auQ59Fgmgr5Tv0FKePWn6GlBUYci
hJqJqoxvX2gqS2Z/OyiEs+fjn1tqu0y6xspBbGr8eFrVfKX6Hieny1+hy2pqbPrsBQMsYFS2LyF4
Gd53smcnFsNhO4yzjfAXs5APZVzItla/bC3yA9p/sR/CbWVRwRlmqAgFCM8DYvaLEYkJucZiz51/
pqqjDBpB+mx0KVc4JJSdxSFa8pgaaF87l/h942/9CxbNSn5HG4Iif4U/eLz5kYiUI0wknEnZXTGd
jES3iGQBddZuFiENv0qXLDWbjQVEC6IjU8IkCfEdD6GqBWSvxWw6d2bYMCc12Ff/Pz6/ijqpdxJg
tUCtnb3S/PmA9M/CqNc8b9e4JoVSlrQ7wqjI9sF70ihllE0didlE5OQRs7sAipGSwr1fWqazHokt
dBNltKBlqV4r2bNQC1MwTxUZIW+kUsxHIbS+E/f6xFq4e6HvYcxFWSEjjmR3PLoZfMeQOW+ZzVZj
sVH/BBMsmXS8ad0KhVmQU8XRvdnwVqmOZ54RgsfM227+G0YED42Eyb2YLMQ7VkdElNtmTdJ/GwZ5
TxbuO1QijrplWXJ1u1lZqA+9zjTFJS98RFH3X8az177kRrbBBd42qfL6SXuKiz+sHWeSNBz2TPWb
9PDqdYFknkt4RtMGhyUvB8wRJvunZS+DiNJ+kT+M2G0c0kmjJTDbUNRmetcT/YP1W9WYAQX/gz28
toPKsfrM2Cglg2WgOMVlfj2ZnxB4i5UJpPuoTwSDPygc7ix9UkRFGcB7UFYYPxdACQROVwCM6EDu
3JfswWE+RnPEoUP5tqXPI1XCN3ram4NljI1JW50YlM9zPa4pJVMbzs1LE/Sm+TNPfyiH+0iuG0Cd
nSsm4z5xor4d3pKC9/D+L1VW0+YT0xvjCjE15KXG8Uu0izVkyaZqHxIrnQJTGQpR7JlQo8eTNMY/
6a/QY909Fp0cOieXPBCuijWc0vnNzr9v9X77Qif1ANTj+a5lbFv7tlCGYolIgEIyPDpV2KR321SM
d1VfrjsFYjlwc2AK2LkiY1Wu24fLj24J10ZNuh0oXvA5tgdqvlYQGBJXW8RaDDQ3XdHxfuF69jKg
kjk5nqZqtDmWtysOavJvb2zfxSpvG0SbZuMYh2vUZut0PUXtdalAhKmGPpZc9XRYvbuEDVCgebhg
Q++MaAFqtZLINIgu8odkOafmojaSG6ylYrPi1orXAroGVqRCPxja8xMefXSGJUFcER2k68eJoM7G
9/QS8gJS99AJxSm3HDqVNw02L2EoKEpY30owH8iaEG7GWab5sKczmg/mgunjIoZEvGOixOwUfwbs
8eX3dE9b2MIDdPDaoGcFz3tMynAQG+yJV+VQkZE5phGgMMl8H2hlxoTBHDIZ7NOPFULYHp52UQI4
kJkKx+Sh/ZSYLvceaFoHq1cGePoBiyDZ66U9Gwvlmn/Og8zrNaqzfbSPk1VdKMhGuxboMPqazmBc
LamqZ+taxgYTeobpgT/0bZF4X4qnrqbwCwYZsLzjCzAN6tNgdm4Dqy3mCvhWXwS/vbzh6Uld2+eZ
+tlBYOPXF/dnIcGn9pea1wjKAfM1xchRfx0WN0R0QFDPf0Qa1g7/OIBtAKa402Y1+jGRNUjEch15
QEsv28jT4jWMl13F++//pGejGXli8zSuS3lRQhXeWMSvY9Q/WB1PyhUY8TSCYL6ffpQICnyW6Ekn
grXhLa6WtdzfrDZzQWj5CtWMg3gokOZNSQ5T0Gk/wEP7ulovSVNHJ8fYUNeAHuL0L3uROCVmGrs2
+OFjy91Sp4zLhZInWYzBo5Y8A9nzr1HXn1AzmIEhqL/Bpnn0msPLu7Drvhvn/XbpCbJtVDQ/vdYn
ZuAjpK3K4SlCPr0Bmgd4Qzhwy5n9pZHori/ACih1xtTg0BxgXduNRuDVBkfnUalztRyuy9B395dZ
XVp1GF2klABsBTTVArEG9ECW2+EY5f3QdtZmfAbBFBizD+W2c6ZPLo115l93Yvujw94fbSlIWxHH
beHauSgoMtMo3EPoZmYYY132DOksrUZqm+Wry0I9BvLzwEBSBlUiIj9lY0Y1ARLf9LX4g21a5whL
XaiTlsf4ImsVlFIBrfIJHN95RrU+F2zZgebQyLfPk0BAEHlVF2VvmkH67M1xs1aj/cI8xe1gt8UG
b8Q324PrUWTDTuqA8+/fIyEyXga1zs89So2TLm0hpB21VIUZbWGkHfk6C2Refm3fhbIop35lQ/nU
jHcO2qrMKQtBzzj6vUPqr9g6bUPQJ2BR9uGBMZtDIz5XUlyJ4+FIorDZG5Ay9PnuabWGYIQlUQa5
9cBbpsb4j8q3knY5Y1XW91mZHN2TFYq0k+CmBDKSHDm7v4byCEZLspWbZLsHvIk/sGmYtlHYVDrL
rVQ0nslBOdpzkYt1rzbkD878qLflIXNIMyDSGQSUhODSYUm4faaMGykrXmWn23LJihR7/eadqf8/
BAUbWyYZPrYtqrC4Skn53xRK+LQNcUX7vDOImeJMBKsHZHQMWTCBmwbTt+Ve8BvhuqsoocTF9Rxk
J0WppaXApD41RLdduGqf2J0jDIs8DWAFHgQBfHdaJ1li4Qth0btCUbY23NzeJpeoay994LNf5aXH
SuNPZWd64pTX+3nIxkxSgA5iqJSw1QOQsAXOF+6JRtjnGj4A7dzIXdUN1LGLftZxxgjMVX9sSPoI
ofy99OVnSsDHmv+n4xuDIUDj0HdP3YfcMJdlFpcqPCX1TexEw4pGukU9DdE1XlGBUPU+Qt4xVdlw
uKptBL74uhWe0IjhRZlNEMyHhPQpEg5HUo8UwyK96QzPkbewLLCe0gx0Lch7x7XpdJprBHuCNW9a
GUHDMo5MsrDHnj++3BwHY5KoPat/6SFsYYAd6UQo2xdk1KhuK+qm8DLFxb4kjn1n/RLxZ82M3SZC
198YCDSXOJKh4i7+IuQZqxqLjVx0N46ELfzvoKR8l4VO2+fxVx1WpHdzGOWzGnTP82UUHJZNYz7a
E+sbrxr7QaVdbfzOFKOthiWS+BOBwDqKs9OZqIKKlN0hp1xCFJlUfdr+NnopQlE4StUPGGy6LyzU
hiOwxjWzC9xUkrJAh+aW6j1nh403cG2hLENs2abHcSY7hxYU7E8deMlYE8FoxZcSAKQhVWSaDVWM
PkAF1H959B5c9mqPcfOQpawyBFp+tyCwtLekjADBHfxxx1UeFxk26/5mcTModSWj4qxF4R3ffWQo
sf6u0ZNEm4qBOqd9AtYkR8nynghCAC15Q9J2JjTejjtLaWjKhBPrBV69Gl1pjd62HZwop9hFmhjm
zMYbGXanCjtN6LFk40qGYKqOuCp/XtaLtnV854ogqIVYF7EysHXp6e7KXfMnnLMMASXtv7pm8C4U
V2vBGCBwTJVEGtOsOXWhoAnURSt4PxuOPxTgtGuBBq5/K0bNDG6VOatlH//doD9nb4+J/BuboUtr
FCWkyTvNrrESW5y4S/164iZiZXA9s0YybLczo4cTS0ZieYN5EqYFPB963eY5X8ZGqxgNUwQWTqht
TXPDQyWd6ChflKKy+pF3bxXRntvOwrHp7LX4T1x7aMepbg/Edr77tnYXmXC9EojparVrTLUzT9+O
aCHmVIwpWPn8pIEE1cZj9InddTNvpoaBpRwuilZePpRGyWKlVyjTX94l8lSCPYijU3uR1rJ8XGtX
NlhWH7ynzoA5bW6fKXihNwYuQOfBw69cN/ffnm1wI8zStOw2try84a6+P1+eZmfOwUqeLOjCq51/
r1hSprXgaBJG9fbecjdOeT5mX5SVj3Mc4ypzzA0lRpMFY9Y2+fPpq40ykxN8dC6qTZPtZHDTeoD4
DJ5WfqCAWcD5TGXRBZcvOEr6JGBst4OVAh5tHQQzsmjXfqhGWo7zxnKqSD8PNDq5A909iyTx3Wee
84nZHZF3AkTkkIxKULhSZ+SbFMIitb13q8lHBe82AAW/79cZ4pzqJt9VztAZqXCH04x72QlcEyly
gE4qfgUgQwt4g3qW9kGuebbGtuJXc7tcF/AAPiYXQvkCLBBJg6OZa9ajGFhEagYsC8Ofk2AcbFeh
YTXhRb79SBAjJxJOhwvJNf2Nx8MuE+EQoGL+q5+g3hNAxdAVyjHO+6kqds0ouEuTkSU1y7601K+/
s68FoYS+vCDsl3Sf0Fl0AFt4MLsHFdF32Y7MVWK+TVQi29P4UxdeFyL3BU+/IdYYr9LLR+uWo99m
VnyJPyhilZOn+xXPkRTm0WNVB6JQ6r9ndAJlthEfpnkeqaf6G/ucBfjqcBSZ9ox2uYjhPVrVjzZG
asWa/JXh6XZPPw4dic52vgpxzuk0tPUrk9u2Wg3Qj3egvSzI1/SzbhCUj/KnLOrKa6PRX4U417Bf
VumTsol0OiM2MlBe2eR/fUJASx70dx4QjiqPb96oArYGFJM9QFB9XcZBg9PYjiSw5tYrnLmlovCZ
VDMY1JdMcvCMeoha2c0E4WPMrJ7rKMOrjGlmqrylPmO+yGkBxaVYZOQfnUjw4MbyUB5rAqW6eoyC
PlU5rIH/1By7LNnVcw1kbsySRqHbWJUAIccd2WziFtocEFk0/qQ7kdXP8KKjd2OHDBm3LTnjUh70
b9yAPRWVYb386TcHESWpaDTds4QdgP+M2Jk1hbyL9+cD5f7lyYzmIHcLO9R1e5ZpP6TfvDPsrS9p
3U2ENhbU0q0WfUlWqEHiAVBuKlgq4sW2rnDfWJmOq8M1TCwzQLmEhGSQRZQhZCM4XNydNYDIRylw
J4tf4weyD+AvjO4qkTSzLQL9bgJPRlJaQTHlO0mkmkiDvAeKPBvODT/dQ2aCOLjzpPHCeKI0wE3o
7fLWHm6zqISEFeRQPo7oacqV/knjpVvz4mzQ1OKRE7cHXQu+w1ReFPLZ+bGhVIlU/GTMmnqSvmFP
BSSOkC7LJm4ZLMzX5oQf+W5o8iRKIfGngELXFaKfE2qOWg59vb8aLLH+XCYd6udcZKmvczapWW6t
RMIm85Q0mQxLWp0zKNT94ocRM2Qbz26tJUhyR8QZUnYnoxqHUkKvOtl1pifWEM7iEwgOmDk/YEKV
Sso1OEFuFaVrCv0/KoVq8i7HAAPITM7wbEYBnlal+egIPydFOH2d0FXmV3cgO0XO3921hRzuCx0H
wi/dX5/gDZ0kJIGUVBixfaYHjzs6vLqvHLw9tuIaCChmYblqsfFtlbyJGbj9s2ee1qBy7CzJGAio
fIQVX7X2414EHNz+Y8s6zdkbwutPjll8hh7fC38B2FN5oWq6a/xte3AxcUr8DXbw1TxrWv8jk9EU
HitUUHFZlhCSj1s75pm6Yztkk9ZygPZbt8vGMYJP/5ZpVIUvnyHIVhux3I556WZro10QvKA8D7m3
eGpvcDvvEoS/k21EawzluodiC74JYSgtxuu+X9UFVRfWBb43dd4fm40ZkxoZeiYc52yEMEbHYiwT
cGTCEeeqfIcwc/CVXPC3DCs4zOoiTMkw9gqK2jAAh+yIwHre1mVwuVIFhSzJ2AibMDwLkOJ5NkUe
Dp/VrZYNnnUbHpvbPfwfcDU++hAOmB5uGfd8qHxVcH4l/2B4Z5pQX5LwnFodCpGRaQB1Da/ix0Ic
r7Awz8DyrVi1PxrTh7CvLM6XaApz/dQtDXjtMvDKFuBTZQff6zrWpbXtfUTU/vERUFMQ56UTfZR5
AvpwgKBxtNgYG/Ra6BoV10nMTrI0UsWrYb5a4Y0/+r+tuUEwC+t+kKYUJmxB3W+IBeaweTFnikGa
5Ah3esj39+RINulju61nIYbdjVlz/j30PEx/ULiR1fUl8ywJtRDtXXpio0n855ES3I3TTMn/fm32
4Ed3aw+0BMXOYNvGg2bHJxK6gb6uYGg6guRdYiA/ESGvH6rcKZhzwvYksZ8xYER6Gy7g4pLwFs5k
skd8VT24PbrdaTv3h7Yn2oM5/qBaVN1pe7+l51VZsxO2j8f7Gpkcr58zACoxjQRNHmcPzXARYSpX
1XaCfPflz7CKxKQzvKVhfEGbkkixg8y1jTdz1bAj0Fw1k9DhaZA6uIcYkBsNSlx91gE5Jnntfbwo
GfoOfzgi+JljIsiNAAkUTmsc/7Ytjc+4oJzsnd7M92Z67VpkVaZfZQ67rHdrsF5JfBPPiizq/tt6
x1I1qoLLm/kBMZcWTgAXwd4mydlnjETq7mbJSLa6OrQTG0OWqWnx0khr8/4+Vhnw3nJ9lcttx+1Z
ifKXFahA3lZdPui5TfExbNXXIpZWkYA+eS/DmLspIp51mp+Wx/XV1yKh/Jr0CqOxinQQvxlw30Ob
f7g9LpwJgRIE0bnnBkrs+AKEBE+5ogH4DAYr88Y/zII7YKbU6hMLrKs0AsvQYj21EsBSuoki1AEp
CbA4MZu56iW2vf+Wdm6zRNKOQ3CL/qmrjB0GzcXCSGVgi93zPC1GTf9wzjQuuPTCxzH2H/3y5LNY
US3GvqllaAXp99qz4HqITm+tYWSVShkW8SFdfCWDIF6yUAzdh9QjbP0uOnZeXn9cGwFB2GfB+3uM
kQXAhrCQ1AeSz09AXI68KQV+377UXnoPbpsk2hbbE0o37kThf1zmLVCWhZ4nxDRoRQhlVHpNwzGg
WGPw+6JcAmBxq/ne8dC6m7/so4tv7tN4qzeKFZdygR3WxPPb0z5e0MdoTUAnu6MEDobPr+todSkR
EQeoo/Cp+nav3qsER1WydauJ+5EhRr3ZKVtRGw3w9IfIeqq2hbFcAqyTkAFz/iFJjHZ5i0Ny8UHW
jtVdtJ5QvQ5HO6OpJqpRj/avTE82H3rH6g57MvcSReBPyVQa2WGp7xVa++HB2Hkj4XU9U3mqKaX4
wBLXgEP38E9hyKknfTu0kb/exlIWdveZNNYZKtly3Y1iW1+sUTfQ2sNHZrE59Rk8s9gCEx/w4RuA
oif86fYIlEqNSJ8SPyrIuI3m5gR3+H0nl/KfRiQBwhMFhfWkONVCLKUmIvVuaeSEQZYReDlC4RD3
DFIXlTJg4w910EraVGTRjzXrZaDC4lGlo7jBSxIERMDp08/atmIhNyHMFah9TWIWdivLkLESx4oU
5/MkEFJxbRhM24zHsls1WvDqt0lfBvJV7I/5F2VBw97OTJe5xZ1szrrEYPPZa9nKBZBUvPZS+Zhh
neTuNFIeTczAeM2Aqm9xJRwFYKEDQ+cS4zMGb9n0fYK5BBhKE+oOSiUhwZdkRdCOuVVTgEBOmeE2
gqAKU6RQXTEx6/0wGLBHthvz+db2uZdgj5+NXJq6vl0M6gj7OO5nkfvVDLT7J25EuvpkCEUEoX5Z
JTq1hihMrsOdbdKMQEnr2rCkexoyr/0BMXBKg7+xJjvwxaYvb3To888X8Am8CbSDqLsjphFDHdlf
//CSGiGmL4VUDyDLTWsuc1vYnsmuQUTXiknS063Au57F/n6BjOds3jM2hVrqUGiboRzBiq8WApAw
sSZvUvK5cxtf08Hb6bsWuqC/LpTTxNQ6JnBoFq8dI9WQeQt3W8AoQsOxWy3pG6zj5hmJ6LUSBN6P
Rimyp7ZcGud9g7gE1MqML6Tvbtdq6YmpjpvEnfuKI+uDqnSgQq0UB0dN7zhLoTvTQG5U2mmw/oRk
H/Z7JPWumznUy2WXe4VgB3ZPdD6oAwrigjnWSrwH65gjpUF43NwyN/s6kX8yBsoWxn+If5A4iA0q
CKwplyZz4zAd12gRQ+T85g1IBWEjnRsv7OzojWXrvUJ8GRRHpxK0KNZeJBEsnzkZmkmfi3oDY89y
qECFHIHiWDmrORfTNA0GOrI0Gwv7Ldxh+x48Ip4O23bt4ZPKfYh3Z7Y3P57sg6kkD0CE6sa/VaGF
9J1DBYpa5SSyeICmMWluatpc6aBxYVbzYW9Z9W+GZyg7K8aYn9MjPZIa1pn1zVWFCHWIdkRsxpig
F6EoHzeH/DxGccGc/CLFBGP97wgswyED5RbWWFpJxMvsOBApsiBHvGcCdKlYSXRe2E8VfWmsLLty
Nnt0YUekcXQ7jUCkEbN2hewO/h9nq/R92vPeYlFcifkDjUkikE+VEO3uNGG0Yb8YujP1aREjcs9q
FEXgkxO3rROogaaLA2CW/XoRekJfdiWk7w4FfpgMpYbCutX5A+++08TfdhyokxazXoHBrb0AD6Cc
NbBctbLwozKfQw9ng1GsJ2y4/LctWHsX491c8VYhwCauDLQ5EC9BMz/bGCMiW5x+LaFqk4e1ZVCW
+pUt7jwda18gywlOKf/O7Cwo0zplIILCEzdxxhk8qmu56j1K4pcb4TdWXLYJDCxIFogZuXgarNPV
GPiac/b2gMYsM//M4njUXUhdWBFHRhpZ0EXElNh2UvGNNO/KzhrgkUwxms3wgQYdfSNG5rSwo4vR
G1xodhXazUKWSGPDKJ3ANH7qZW0FPEeSHpxAX0m1gjVMd5EOW2g7IVVMG5aYE9K7bVNGhWpljm1Y
81WwG6cf1f6HroA72iNao1haQ1RhNKnh8IrasrSTkQY02PolWKfaI5eie4QJh0Jc97vzVSw1Lln7
ByC8ZyxDPgVuhrF4movhSDxzB6w7Bkx0EBypA6JTksTXFHK312blv0pyP2lCcFaB586tP5+0WoWu
mF2F6/BuyChYMAqNyLNBNuRoW+HxpQKVhpt+bN3StG6Rl09OYvzKDp9lqQdMSbYaVz7XzkI6VMGq
l0WpF+v+8Z5dcHuY3+/Qi+XvuxmXANEYF4QP1kYOsoiDICmTUXrR05Njw7Qx/qayETPgVYQq/lRB
IObF+2c+vYm2WLe83bH6hpYUJ4aoLIOvcRAGeTN6r8E97qeE/s5QXsGWJ1qgTfxlaXRzC76vBaqO
O2LHv3mIT3o7f5ogcXth/yZG4GJe7z3lfxHPFVybX7AGTAtCBa2S/32ttVF4IAbVTk4oIpzCjPz7
TXJ27ioaC0+7i+VeJ3lUAqcbUfJMAl1xpxi6f9jlNyxis1UtcuGvE8of3K6aCQ+sw4jfbEUxqdef
ccQkxniz34gBVWL8t4UpKHb5qghn+FLied5tS/zBfPzzaYVCuQJUjZCavczjFp/Gk5RiVRiDJRNX
zb1ykODILzBFu5O8/4/dEk/CoZkYR03E4kEd+jIeYu4XNZEtZ9CSyL+BUCBV0P14fXYGtxIeXofq
I+d+dOK7kKgNtBJohTzvRzMpQeVu/llyAM9IUJUddfqJq4q+xjwAXbaeMJnmOwVuA6IMxlBQ5EJl
GF4KMdHb4B7nEyOzc9tZ8ltcGbuAN1M0KVLixnSdPvh2nHx9ayPHM5v4/0kTz065O/Qwb4g8Q2X0
CEwAAgTVnXwKvsfPB4Bx8YNM7HW7iwYfMFvRojP3SzTHZ9GuCHiYDRht12cTX622GuZ1tevtE0eM
Xti56QCeES1tkzlrntA7BIy+OeR5jzBQAJ3ucNKX3eIJNYo1RniGSq5/Wgnubu7WhBIkcL5ZLWpT
QJOpTrHY06Y+cQk3XeStohyRWuQUcPRZFvONCpv4U9EiMoQ4fgd3sxQYb+w2Sa9QuxO5YTrE+t3B
Zwadh2MA0e1bRoZGHHXyykMGyOzpVHnHMHNm8JcBCNUI8yURIphgzrV/VWT01GHxuDnB3AYkRWbI
onyJXDyyO6Ups9jte1a0LBgJbEXNlCoTqGDr60gmn1J9zwdpfTNRTUvg/XVG5xeCwQz8SVRh5Xzv
RJBM4I9gmABQvCs6d0EPRFqJC1ZEBrGw/nFiz3qNWt7ymqbXnhN+IiLvcPNprMevazm7alLdXJ+P
uX1JpR1yFSj0Mp7U8T8Ve2OCP3yFwdaYYu4OJeHlZOa5TkMSi4hvXeX8dsGD+OWDWJNHCROE0DXY
mKI8b7wC/bshvNSM6nh5uvjfwdzMU9uNctKWxn1taSo9f1kthW6XyNXGc884CIyzzof+UVGXaqH2
TEJHA+ArGtbFFqRm31+bAL+bRZaaK0w0hgBi6Ss4NVbpJVeodWcyk+BkJCaNVSQsNEP8FJvONHJP
Iuoc3Fm51VnddZvEA3WWjmYrWcOrBjisrYxI3dVxs+uIKydo+j/PI7tYzbpARp/3djGTdlYZ5/cx
1tvpBk2mx/pfuBJQRRyihwYD5+D3F64S9eQbdLtxnfOpx6PW0oyvalTkE/fMpHkv+aC++ohgAlE/
NOGbWDkvzjMYJqG/gW3h5FlBzZ0kI+gQjHzYY1Afcrp8wrX140jVzCpaVrUMXdmEVaKhPWSBf8a8
KdSC9IlGYHFWGFvaZFNEL5nLrgxUb2Zi+LVtgagmEZ7UiP7cMKX1m1tH0f5Doq7CkTabZno2vRnb
iDjISvtLX0EabJNYAnejQlCmltHAZNykdGdC93BuSNxMhND5lhKLLK4WQ9bptQiTZnQBtYyD80jq
GF+FDpr7tFpP/ZdxMuBRj1+N4RwwDOiIiXQdH3PebhNhV7j8dE3zmh/x8OYqSRMPeu/6t/ujoJQP
KHU8lc6wpXb2f7yUETUEhxNrkOKb1woh7QdIjz8JfBRMmX1LgFl0mBucqvuLxAkAVUh2gZ+IPHvI
ML6hqtSMz99ay2zDftaNKmNPZwgA32WbchoHwIq5BWXm2vZsVyyqLwVjfANBp9o4kbpv51O5VClH
Rola8mlXAIxCiQ2BPzoA4qvi97quOmyxW92HeIjTSmeRYcHUf3m+7PXeeFS/fBgnE5PY83ZLJcNM
Cf0Di4i9rIFLLq8lgDSljh2N9LALzQT896BEB1w31ifJk6PgsmzCKLeNWLzINlyAOtpl9SP6cYHD
9HwFCgPHxhwQKaTrgS1gLMjWOv2yCK9STSYxC41czP7cxXXfzmR0DmUb4z7ob3V5g4y4FYirFa8O
NR+ezC7SfZQIbByrDs9zfFpAhM6e/JIY4iT5y7fgYd0Fwhx7wJBmfJ2XUQa/AgGaXcXNxVAZpvwg
27gm5blIVtpNNWfDi55P+LiqK0UMF1+boxnomoKRn1o0RNG2vtxIGNFGCugp5XcG5kgM2EAPJdiL
LxtScVYZrA7joIQGKFek9kjlNO2g4Pmyu2Av8bc0QiJHDO2zXf7oBmQhtkqR3DPOU+vjtmb/3+X/
nuSbaSfXF4jjgcgefo7TIHuB7Tn2HT6yu23QhNC8/tYGqXWA4DlHj56mBwGBSXKbdtkXnp/Xoqk0
7meVT/3osyXDP+FGyIt5NTuyQG+IS7zpjIjSYW3oOOTUbh6csU03Dk2v/9RO4snQCoJNwpfiVDI3
4NH6m05aJqeySckT/6sfXhwK54cOW7P8L6Bjn3gBZe9rG4BpYeKN5MiHxVllfN2t+UexwIXF0ZMT
qLoQLrVClS4yN53NKm8zG88spRihh3uLVylidzMzQX+4K/hzAztUx55Sx1Yw6FhMp69V/dtBEW1i
b4cw95SljkdqdUBI1Q8PZo3jdOQhHhNKZOSRQ72hRcZKOKFTT1JzkPL6ljlHH85AcmvRURGG1uG3
Nd3+CrstIyB8JW+3RfqHvOKreIaI+zp7AYBg3nX7QDAbxHVEFdcujx27CSLY716WkLRpeQQ8+WWu
YDQWVJXkA8YPhPi45ovR3ceqUBCsth0QOZXQqvFgyXDddWNqAPvhf7A/VHxbJ8Bk81JJ+6aUzbsM
srTiP79c5FZYELhIJPM1FbaBhrMUMYdy3to0NP+TPrZPbHCan09ZY7iNPmo4ah0FRx1Gi6yjk2oI
j5UygPTodq1Ep87W5wsdGDhOx3rDA1ogOj6IuHMtSRcxBESalY3uHIFWpL+ERFZhFTsfvBc2Llat
iUTXXwoV3S7PnY8XJWSfuVq2QXxKIDWnHs+0TWfsjwQDUv+QZn+6uDP58oyrV6tO4gsbmUaaY+zb
mzgoNytEC2JmCLQc5HGlkzpOs2kGNrpmFXjGCzjZns2CVe+OxvPHZOGnab72Ma5fN4OEyCh7nu6A
bu84d3HKaPLmNUDf6x7zl97+nBtLe6v0MHWT4cMh+JSAtniEW1/61QJnaFc0NtsHEAWdqfyI+uP3
ovptEpUHOkh/R94oPuqXb6stjMpBt2BAiAv0ZHWhSZMHVo7xBv8RDSn/dL2O8ZZawkKvKPKyHGvA
NkXw4wFcS81ooEdJEJrmY/nnoEAPqc3IQYgpl/IK6UvlqLsV//fgu0Jvp31CZFvn+vfyWeS1lWvM
jXRlVXhU/7Zee5oricS+8aceeLBDHtHt5EVGajtYeUenL4HEhc/W4CUbXNZVNTrWFGpINw9IfqL1
4wVRJLXg9HMB4QdSGwSKZzNCE/ygN1Sd+rmJ5zRflrpxMKvrO+XxnoGpyyOl8DBWQiTmdCFeALgn
j/AEz7jGkLGoSBLexT1OiDoRrkEjBahZp8KOQJpx1fmj+8HIfSXTie6rvqdiNKvng6Y1kbxIlULV
EIrIY/fHnVgVkcStQRS+f8NNGgz2gOSbQJo8OXRVH3O7jDlLEEGqMRMIIXHXLPfn8WpXC3p/y7RM
msZloTXAGmCDCvVjuc0j80wHsXMPhrnsuO94r8waI+uvJgKFY7tRHjuFYeu78uSghESbuQx/aJvt
BxRbP/wg4WLUbJVkOEIEJ8hTyELmqTu+8MTJUPmHP/EMV1E3j1rzsZOLYrfG5RtuHgeOAg5YAOcy
Wc6CLHAxJ33iuSxetRXAzAI8FEDuKRkAcU1Ms4vVT1EGwOs4VLp/ZVc4YKiRCH7ecNU5nYqKzKUE
jLDrAyt5wnZHUj5UKt19NsRRw/BuMpJ+HYZodR9UdOa8Bsi5w5Zsb9sRuUv4D6GvZ0bLWCcrgxBY
Tf4ODtK/1XFtw6+1efPn9ki5pc0QrZWlT11y8hPTvn2b/owHS6tk0prp6d5Pc0q+bpaYrWMvJlSa
XP26RmuXgl2+T3Mz3QUTG6kjRR/Br/0TTc7auqDtB7vuEYuNWyY2bKAE5s6QYtrDZ/EmmLTAE7Z6
p8saKj87Ucy0MoBL/Rwz38oW3sFrqFr3sfS7FfcMp9ZpRLezQbhjoNVCHlqg0TDa0fF6J8zbzlY2
1KczkmkGYf4Olgt/VZQ54RHmdo7gA/4jBWNccb5pGfFWatstcZGgnjtCkKCfd212R4P49rLv71Me
FBXVyVI+lsKBP1RLdK/4sNLEpZSVZfyWwnTEEmJCtW8nJTdB2CKW5qQp/d5aUyaKTdT/YZJNRink
KUlHsj7hIdQlG+Tjhcf+vejMHn/34gpUzWgbduRwNxjMqZtqSAnuzQYlb3lWrRT1gEYLn7/g/COT
yhpJvntjEh+s6tvigxnk1L3G85ANgeC7+CH4M9q1OWfz//J6lZRJm//NKLSm9aHD53OVcHqCbIjF
E4p7voxrcSpmYjQRYoGbJq8qhfVeja3MDqJeyzNXpYmAC35V83iso+FE9EtCfOZ8xOoyU1T3he/a
TPD3oBmsoSZC+CRBhgzyWXpIWAQ0rtknBr6lhXR5+aNNvCuJeYwGkqNGuwJzoMyCq9+JCp+Sog18
MEkiHhu1sKpe0uz92uKNoJ56kiOiG/S1n7dMeAPfkLOjClE2SqP69xjmaS3rxMJ47Fe1GN1KImrk
jb+dnHUmOI49DnXtJctr3T5wcER9XBtiU3v2jLhdZ8jT1Qaj7QkQrhyyJbcFS5ttoPzXFVYif43P
GvTZ92yG8ZlOYxIbuOwRBWfgnorqwK3qsL0PfYmtDiDto4wwH6pomKZs89c/nEPnE77ha2bVJ/p+
Eh5gTgH8fPdNgUqMmd0d/biGgCb6j5oPuBsqpMxiRT9FLoud8YizYNGY+X19ZVWfaGZc0AT/eWEc
FkncpB92f7Z6U/5o5XU7FFHrchSASRYi5hHscxZ6jYngkAOyYdeWU6KtQ26h/B9drA1oZBthwON0
E3hXWLmd00Hx2RiLHvqZioPV1iKpIWR4It4Vi3mxsHiW+t39GyjCulj2pAvUYD0J2vVSWiWr96q2
rUewvbc9jZT1t5cC+vxm9ZDB1gxf+ZXEpfCrtgkU77oJJXir+S539AHxk2zqa0Z7C1b2+yoRt+Qy
6gnXm4ekBKFKObIgtmrBqxldVfgKMp4v9qJWW3elqZ5Xq81m/UuLhhZiw1i6pjsVcVIVAagU05R8
LR2p7psu6UGIdxD1QUGD1WcjizJY5EkD/pCwhSHa2tebXduGGG23/o+FjRE4eWyx1nV/ebnpGZjW
4MIpI5o78xSTxNoypX+PntxHju7rtNxuYG0ahRgF/YhyqWqIyJOYdQQIw5ueyAA5WxL+4cz07YhU
SgQhNQCXGuBXvgMrYmkAkcSPcbGdn3UACpk/Y+2aD+PANncVJWeIVMI8Sglx7uk37vD5xavdGyaO
PdHj9q8JCMkjmbSFtrqhRc07xOvxMKswaFdzwVMAFenS9lbco1PF+xhr/NdNseGE933sS8xvdidE
bvXgJU7FWfMTP2vqrvbgVINxKOSiehFbRBEjbzpX1DkCM85LXa+bBxecEHIxjAIkhZg0x4pQc0xN
iM1MIYcgV5BlKFKTLywR/9qoMbGlRqMDb58W8KnNOLFEaPMuxhow826rK26bNew37ILXnbY7Lg/2
GDAxkSN14O166Im9WSungYWmnm1pd8TzpBVHfZLen8m7+x2iQIoH/qC8Uhnk3HczLdV2OX3GOxCF
+p4tX+nmAHqfAZw65k6bja7GE6b4psevvtQvLFJf6L5gJGQcFI3jJjnK1M5ooVmm+acO4R7c0+jQ
d38YL3RoV1qcdcLfZoIPFew3C0HdJGVzflavdbQ/qdbEwjuBgrx/hb12fXbqZVoT+QD5UUuJmHNj
nh+vDKqOEs9hru0efhrOVZeaU7O/yX67H2miHxqITGudQhe9zrBbPqJfmR3IBpZmgCEMpkGaVg+A
ko8PydtDI+cigwlzFNi2bI2+J401Kj2iF7gwc8H8kXVuyVkowg8YRC9oDHcKZZORaRnol1tlYxMK
bXg9n0rKYbtVYJx1x1rWR0Ap1YaiAjKePqklSr4iaT6SuniZcmDQvPrlYkTwbELubps5U/kpMXcS
MuQhON4h8Fuo7r1xSKVyFL36tTfFcGuI6T8OXJ2A6kPW8ALXJM7s6HYnHLkV/9sXWdHeiCm6KsPW
x5F1eJWFMCOCYLkxypW9KQMsQ95qgL/Td9UhrAjwEVIM9dO48UvUODYMrjGjGv44USEjyrA0fWUe
DpyZbJdP/hhWf+PDERCSwRkK7tXwbLTBXE5nr/m3qKl4oWzii9hkiHoZh94ostF6yasdRiHuFFDU
/+1yvZ1DQfFhJxXkOM4v4TcedPXqKHWuu7LGfdCqjxgznd31DUyYm7ZN8EMlZ5iycjyFydouhpEg
IjSFLdq9rTikUaSB8DTu9l+IKcpjYaVYhv/JNpaZGgL/yAI1ElbBQkkhX+nkL6+k1r29qwJp28l1
ROwdMHJ+eL+rQoMn6f0Ab5NI4CnuD8JamySxhPkbxl8bzH0PlZ3il+5yQLMRKSjFY2YT42j45paZ
aoOMFULiAJU8UwMDkVJOMUOvxeq0fbG1wje9n9NsGeuyVtosy03Di3uRsd1UM1vNqvQM4NGYYY5x
dvWQ8FbYbEGAsehMjvBzXZ5iAJoqM23n+XAkaYLHRCPnkSl57E1Qyey9yPCNHCYrM3Gt7PnfBkTi
uRNXdeL3dQHNtSRMpi/OPmTVkncREes4D3SiPHothIl83BmHrbmjm010wqLg5COVz3B0xq8sVGFN
QdlkwfaTM9P1ypJbm4mB0uZGgQbfWH7vM2etZql9WoRD5+iHakevINRr6jhBqYVpuMvyGsipT085
nSoVbzCCY7M+jV/0/jSNiGn3hgMFJ4pzWjQQwlHoGqS/3bVWDveEU2iN+DsDaac+Z8KujxuOTGpA
kWqwEUevf0E0ijswQVc4rb25QWOey4Ot9EHvAZle1M+zu8Re7dP/vpAPpyXh54N863GKFajjqhyu
9QZfKKiEZOzStgwyG0Fj+GACeOHI5XObZcBcUWcLgwOQtOJMFhKQQBw/pN0nBzpoBkfJMasodIrj
P99mEwZi2ZasppU1NXNZafZ5fxfL85+KUmOu3cQEH6gApEqkLc1gbLKvUoLbdWDe55yb5KsZ84OV
I/eBAXmxEH4Mv30kUM4CrUAgiwK8MLgW0X+QXmXWA/mLYaMLDGEWgqc5hObfVFZ2ZDJf5hXquWkA
gswbVfcNCwkjDTMyeyO07xpSeGZVo1lr551sjtx7XHn/fKuztN78MRWyFZEwj1Az2HJvNwTv45CT
qyDIKGCkhQwHz2RSoasS5+pJY4eowpIvwHhzIbR76FhJozCVEYDW2TZ4WN6/N/pI/ax/tw+tDegf
OuDuCt8CcQ4xt3jk7aOJoF7q0h0DwoPEWB3H9jdkqEV+CI/IAhbsbMzpLU5sAdFTQntltnP/a90r
fMcEjf0pBIa0hmoF+bHZinBxgj5pEHzmFlIfZwgy0xrqFpP8zule0332dULnUEajsNPwvnp5jzGi
SKpxzBM2hyPwDhNIzkzIgwxd7XDSOW6tj0ft8UUMB2SUxkA2ClbW3nj0fv2e6A4RurtZSkUXJ3/n
9RHzyxM8k0eYg6+P1fNT9Y7SuERjYit3Su+LlmkyVfinlJcx4prGT1nUIq+3UowMXZRkd7XWE5KJ
I8rEhugLMa7jcti9RiFOZtX1iTXV2i0P7XFRBZ7IfMy0laA4KSomPnR4zu5Gon76HbIDsEOFETIz
4zFLhE9Fs9rT8gXgAeMjN+BkvVzj/LxlHGfXAX4gfSQ5lt+n743OD2J7oozFBsWzbk52MxWdrjGT
S734fi3FJtyrMhWUsTZp2OtJq/i4Kv9O2FdS4FcrMciH8xtb7sKcPX3jRWzevefhyK/Z+zS4nH5d
X+SuxwSKGs8xPEAcuJfzRuzozc78jtDfVibkv/CKyG83EB941QpOcqktp2ukG0it4zomlqOHQ3nH
bvS1wmW1GjdotlN456BZdctk/87nl87R8MyRt861PEHkxRLj8ysgpXd0AK6IWiHxOdekvvjJT+Rr
4oI8MSbTy6KqhDDNfHQTEx3+B4dJtvcdYn0PWToQccDq431KqgBnbu8pdWrI79Wst/1hqCG2lGDa
tUWzcetFij6RC/tIwuXP2MALYPf/pJIT4VU2YpJ/t+jeZXvpRFGtoinB1hB2zNDqTUeYqY2VRZzY
sVNBs5m+Q2VHh9rSCX0vMyKkwzMEYUepJJZSEloMuNzkME/PNs4u9+7TBtRfqmMBZXX0iunINjJN
2om+y3z4SRIC1S7kjYrPMrAqhQQfFYqRNEYvu7dmhO05808T2dCTWqHNWzuPEo+P8huwz6x466xe
C8zpZ/leZoYfQ2lzu9Iz//ZW6H8uL7U0+H48QvpCBH5FggFRh3KTGdIfB9B7P5MEU/54hor6X1Zc
ki9ollz9cL3MBlDgD3uiyqDgjTebObj/tnimYOM/B1Yj/kRjAv3YAwvmo0pzsIvSyXezfvmLVu8i
rnGAkwdSRn0951hWyHC5Jip5XL5Ba0dzP0dzbX9MsjibjaXrWfc9PPHbdTgbcWAeg7/rwf86qPzC
3+io6lm4VxYWE5eZU1FyEupwaYxT4q/JYnMatBq9AdJRSN7cV3Vk8rDq1lD1FpRWRQAA7jwkiJVy
LjxtayiFWtnfwrQeHDIfVNeuNzqriawcAeQ57RpPtiJFeQ8T6WG1LSdjAxnCPyZ7RqOFtct0T+kc
jLzT2kLJg/urSvFKJT2pM5BobO6761y5EuP0falubYhd1dB/pEAc7A0TG7lMxPDe7Gsd+Oruz1hX
XA1k10o7yhUVHuaY9hQaDBze19eMUok0w92YFFKf0wuu98Vr84Vyy1RJgT5rk2K2kqipH8B0vsaQ
TYGU3lnm3u8P+oHyW3yLXsTTIIPBHOpE4FdYXsu9Pcfql2B74L7BH6OuPDQk0hm3hc6n8nAz+5uH
kmFMo3cCOnpwbr/XY+eLnGJpkYx58gnzm/s4BFKIHt51sPe/KAhnnSayor5rHtmDFnzqaKnrwZbt
CyGcGXqfQ3Y9At92H7mwDfH4O3f974tgpUv6LenJexx8gsiFqlZR/eTyumIrcecWd51j8i7NQ8J9
Fc4MNrwvhWtbYuVCl4EVHAyIRAmKUK9KOk2z/ttAZr6Q9dByi97ShXawuRX4ZDG6mtadw6DCQRhN
9/Xk6r2NMsj2tcmoB6v7y9bC6QHG2AcCvlFY5gPBKf4i9kEjUFpYhIYTTYoyEsx0JeSXerdtHwim
R5tAzNhTtnj6TTboiiKX3QgP3MViUEOXlKg8CYbfHpL+KWthFDFD4kDzgcQfNcKQyAqq3CU3+jFv
3k3bC2Dm7GGccaprNZp5SuPYZK8Kl2rq5ieO6DTbGsP3sJB7ouYbx/3tOsPQgzAOxvmfqozUV3gX
bonir/4AeHkXjIt9Dnto1OJ40k8sOi00B6xuZqRgeZCP+bp3hDzi8e9Ep5Eu2MtWujSvBHnn2KND
PeY00rnTcA+Fbcx7qEOQAaHgHGsyBLCRZhYInwfk5pEonEtIGkGSGJQHr5ep8HNxi02OMfdyMeQ4
k6gRHM9+ZWS2VkRpA1W5paQDO2iGA3yhjY9RGw/nwkiCmhpoBCXR1sHYntVyDZX0cvOxtoiSCITp
jb44zu7trWPdck+mUVOnSWaB+PZwswqUlUqy66WiGVRPizCHm/ApbiYYhnc0dmjGoDrHZxSGiXlA
CZn98mAHZSHkem3E2aw7+QpCu7VV72kG2iUnBKI3tu9c7fNS8E327hCetyHZOgAl9BQVpsXjK2vr
H70HebIpLWUenlD/kGVKx90PwUoDUP+iqQx9lyCwKfIFlE8iYxwqye3I1P8+W1dj55c2BCdP+4/s
Pwh89nJdlFOEyvg6+9Cfy7I01mBE28ROrzeHjZ8aCN11btG8Xj971Sh+Ajqu07MeV2V3WncduE7H
6pPZIwTEq6tDOV2hyIl//izF/iUerGunLiVR4kNHGgebQasKtcx4bQu8dOTGHOe83QeBK6XW3rgn
FIvKdP6JVm8uCpaSVU+FjdcE7gyxJBGpGpJK3wTKyYncudmm/ulNzI+rYCZR27DscGCVb16y+lYz
RipH1rCaOYn8IOckbFtCTHUZvyY714aRQqz5DhkADTvFZeDSh23Vo0sx3WbH51QhjFZcuyVM6pS0
TjSCaYGMJqS7069W7dGJ7rLSKu5TBeWMZWB3CDoBBc/GHMjPlirZMX1UjURSOkkv/wZVhiLY1LS5
GetedqSr/JQLuxv6M4dYUM6VAYskXKlEtCur4h75AMsgFItdsxj9g02nErZ2U0PsLmTugSNu3SH9
zcGJMGIsRISlAbiPYSl0PmbRWl+/Gv5wUuf+K814PANWNZ1UI9jKbUjYLy0BFb/RWG2Chmr/yjFU
2EmYi6yDZeueA52o5TVJQ9Kj3lf5rttaxd/MFQnVOjYyTKYdMJaSqcW+H/jQn02IK+w3lISdVyOH
uJUVsh0fX3HWmnXkzQXkKJIyKxT/ICMa5AgD30fFwiG80AQfFvtfXnQEJT8GK+xW3VHtRXj66R6p
ruUdWmUAaCOg/me+t4v5kr8aZBWzi6sUD9pVfdIbVSdfRW6kLcjxz4qox/9WaoE2ciyd7rIpBD5H
PMex5OsW3K8GqnjKSvd+psOAkcLgiD3qbnRCstaffc7zGeD+K0Gjm6afjhdgv7q9gAP5cwTpzf+G
ht+BBWNAJoZK6iDiuXR229VqHNjLYCNLUuQHewJS1+TdeuJmy1KcN+Yd6X42l4L8UEtl+XnsiT22
agS/+L6uYuLSy2OnhkrNcI0UN51wCg+RFHguIacgVRl5XjRny4iOgNWRH+zJw4pnWpVuRiFXMQCV
cUjs24x4nJGprwnb/PT4FN8ahpK/eDs1MjfxjwPL4w74rxbe5GnESM4xDj3ErTF5bLEGFU5lUBFT
rWONoegMmjKnwhR+fGHuYIdxXrXE6tZGI1SAnCLNQGaQkpeznBSF8Uw8SnIsOLAIiN1DBtVPD4LD
41MoAaW6qaEAvaLzPPeTt+d4w+oeQxgMON5b3Pj5qt5fIYxCxlVNuctnZ/qUX10xx1Katw+Nsowh
qpQD2rByEpTc/Q/MxfnfF4XjYWMG0zVE9pjiWm5AhjTrAWEWEWCKrccSx6G9FbAFQoXIfGbAX4Jw
poSvaBNXJ+R7Ans1XFuIRJse68qlgWADg9Qcam0Ap7/7MFUVJqgr81QCjO9dXo4SbZuJAoZTnrGk
kzmavOmXuy2zr/slte6ZDA+mM6BqeeoZBsbe7LMNEwBO18FsmKskMBe4wnnxdPVBFEaWsAvvVN+c
WCCvammcT8aXUKrbbsT+WIL0WOzHqEQNRMWBNwJC5uaCjaYSxwjdXBorONtnEjn1Hm173vvLBR+g
txjde/po5culeGl5qucjwxeA6WUYPgaTlbnSJeTU2iJY/6TZDMt0mGa5Y2+kZUD4ggUdO0emXDpO
G9x2yg1PfoKeq4AmxUJ8b8RPzMnnUb0sZ70Zj8YeR4rsA54LLdsl1X3Fjgcn8vm7cLWby4S5yjUW
VneQlv8qYxUYUDMmiIX/QK/5dTiEZJlRAAaNkC+QXHp4Nsl3Wq6w/v8YEjgXwHNTu8JOT27deuT0
k5JAHumjhZzGQkcrEAJK797QD5APQpJA5rGiyPYltHHmW9GJSFjWBBDCwOizvpQV3nWsnzrLIS45
9l8FwGDBBy+s0loKL1HgX7QBD6Gx1WVCRucjLZnDSdbCohYefjAKg5Do8mZLx2mBx/pxoQJD7tSH
FH0wHulOT9tu31eoJVORRr2K28uirZX4AdHj7r96WA9ITS6MO/AdVgLy7mlpGamzDLYIrTDzThVr
v0g3Fp8NCMzMmbzqi271EtUyD5FX56mDtID9IJ38rrF4Ke5WH4ne6v8dlUb2lnFJcLB1az++K7Fn
TSc43IzQUWo4T3XdWoiwy9Zbgn7K/s8Pbg0LbKgAmTGvsyl5LHvEJOHAxPVFIJdw1OlM7LT3gRXQ
E26XyyLa/Qm3xtxhPStDZdDxzlpAponW1cNg2HMqSQ+wFcLoh6nDxKu3mysTmj+yydbD8qtzMWRR
Y0TtR+PfHP3g0rW0uT3TZAhD6pWRBZCDrbzyUoyOCgIYM6XOzcqUBv1l/f081xC95/WWvehCqR5G
gkmxhliHfUNL7UiDp61vwSXtFedDFCmjjclYflyg0uIJ/bQdfDdCZwbk5xtjELSe4HdhTxOpoBaO
Jqcxi4Le4ZksMLvD2zw1X2hh8VoLj+qY2N+Dh/mpcOQZoVHTjsmiWAy2UIYzbUloLwuam2iFkGYv
bX3khIxDWsPD3+P4Rpg07HF+KHixTzJGnBkYETLJu4zw4D+c1XT83xb6wcZSm7g3Ro8Pd1+P/09m
a2+rv91psS2lKO//f3um/RENqFMIHD6mNHK9NMmJlFsy8HNGZ8GH+NOIlkjlrARD7IxKsoHAUJ5k
5zeYk/YzWdh3+kfJweBsVVI6le/kiuxIBwxf6VR+RBGOYWAC6gZNeIWc/NXyT6hDwUe9a/EWoFGe
+ShGbWPjyPLvG3bBgvcoyPTHQW3hih3jt36m1qkAfiQwsEqTOpK/VbDTUhpYzP6zNK6y2yFUfPJ5
vVqWmHQzB2TyeCkVJ2fpLA3Tm4YZFo8KtzTP7Dbmk9NGH7ZeG7DwxScFIJqK57iGE6gN/5t1OYdg
VBBQgWkHpw1Au+aQs3qiMB1P+0gMqaV7XctD64KFF3Fj4lwedg28jutNPEnZh4xXp2HrQALeDXUB
OMfwFXgePcD4rcKrRGjEEPJzCa/NDpJYrVBoG/Q/GXn+IvMKR9388bcRcy3ZmHCTIVI78dabb2up
BcJ1Fujsta6x3iEkUgwYK9blmszhfH5cDqOC4nxgSRyf/SBeGqtKN4Gc8Qa6Sulw1vbaPbVsnUxl
hmhhticREgbYLfTZy5LVym1hDzI5AhpBWD3UzVwqzWxukkFF3eT31rhOzRzSH1+sjH2V6jolXP72
kFBWr3y2UcLryxANn3lFex2XhmHqgiuHjyS4BTuf7eaO3Ip3OYYCBk1HR8EtOvPc2uGFEzKaKAQE
y41uuOplrX8LKNJpH6l9FCixpymSm/y8AF7Z6Bw3nSxAPJ4U4/WyE70XenG6n+GzKHcUXsln2kxd
o6ZdSReXcduLJYN+HAplfnbd+DBoo2FSoSvWo459xNMR8mmOZeCCiOoKQXOHzsJU9vQ1qoKEmepZ
LR4O1AxFcK7GKmgpPQgBYoJR3FtkMH86+j2cWe0OejF6ngjuwJ4K0DMo/Gv4bXLdQ/QVLxhitfE5
+9dOyd8wgbKbktWG0anfg/ID1vt4URL1KVKedcsLzAAY2lownCyNnXUdRO7LkECG6fxiUA7JOU9E
OOElRnpx53EJKBmSrSuTJ9HdvoSnPcFtgjAGkabo5IVUgBkyEggrWq1gqNmKmyc5KDhi8U020B3m
cXWBd3ZgOggxC6fKVwOsA3kNrjJbDo7y8pRQwgfSzw2QugjPsmGvfcvn1ue17TgBBzl09/AT5fLn
x4TQo8BEgcHeZkUet5RkZbBc/4gTjIifLp95EaZyPAR6i429DqVI/C7l4L45G78rGkJyFWQPJf/C
IWRkkdFZdS9NVLSsBoZ7B7KjQBWviL20c1cGxT9L/FwSZUdO9nkwswbMdR80usdCHW8vXYE+aE8i
i0MZ+eZEGNmKLVZU/nfo8G2pwQrexSYXlrrNYlqLoHqnV4SPeUGQZ6sjJcUiOgW7ejITah5OsypW
96yvlIxYPjQpiO6tQ+Lv0MIthXnmMqWmBXyi5ErcAQnSGJrPX0H7hBZu2TOGMwmP83QJTrgwbNsu
U7DmA6ZCEG1nHjkhFgWD5rtla79TzsZIN0G/vVB0mZsVMywl9jSTh6SCQQG4nKgP+kbJN52HzJYl
RaMkfdJVMuVh3/02rql5FE5AvLomFN956+SkA8A61XiwCF694ZaidVp3L5jz54KgKi6nKGakCqJw
fY8YkpCy6X6fvC9xeFVE+9qWDZBMzRWo2RWNBhsY06tGO5Fz1d1uIUfcZhkt/lhGWsqYC8eLp+Sp
kTib97uwJgbZYoanQG5fzACaRT2xsZD++330UIm4fbMtqfpl/e9+Lv+jrIx/w4le5Hpl6Es24boG
m2Zsu47z1n3EMBzjrvvc86NNKbt+Sqrf1QJd9M39NmcZVF/zjKZUZK6kmx/RGEZovlVeEwoG4HvX
9gBPX5wdZXHowMcSD+6pmBq2vqxmvtV4uF/jM4iqMzMXDLlHtmj7Xb1rMArwqGoX97fKcdexmT13
YW748ZTbxm2d+ZcSwHc9ynDlnuWtJUgN5w0D/klJzYxRioVvdjeryZjc1OiQGgwv4PSmdfKAaI6j
IQX+zcriFG4jVtnL7FTXkl84xG6Cgs22sgXOKduMzaR7vKv8S3LAI7wNTfxlEIWORUxDonQZDq19
wmdaHHI1GcMW1k++gNO/CA5zluvEUmOEk1Phg2lTVpgPZQkJQFDJXnVWonmRdp0xIVVmiBrictLw
ciqQxy9Idq8zD89dDvsLg8S7h20g0QKbwMorK5BsAphgWQaU40E7DWkWoUWmb/PlArmb7YNOgjTM
FxejF76WVlZ4CwAwhYgTTHwsFMhyDhK8W1Fxl7nAk+CbP8zsIsqG7Rc6XF65pUQeFeesJ35lcPPK
TSxbslQxGiMGWJHC30YvcruzQR8LOhTVz7JnBgJqVOZszVNkkL4oMfOCN83Yh9SP/wBtGMjDPY6q
yrfMaiW9llIDUjrFC9uZOv+5JowfS7Xwpt1K2zq8J8S84i42ukTkfmtpzitsqtEGrSzz/qToNdF5
P2T723g0BvaWeWss5p+nkcfxNIqAW0uNfw0FdqI4PYS622n8fPKGHsrKhsQqWRLkvPAcXqA64oIt
6bgsqJwSxGGVNXC2BJOlMh1XU5I+u+fuHWs4QgdCidZ3bxaebXA92YBs/h6bwG8inlFVBdzb1SPO
kL0ZAtF3gNPA4W3wLSdtvaA0SkvLv5JXq7pNw/DEi35TjMm2Uyp9IDUFnbPr3vcKA9sTwLNQtECQ
pluZyNGXHNmfptZBlQOwhvNRHPB29TYOjg6T0BvTUuccLQDHct2Bt1NwgBblw5+HE3Oxdl9AjBnH
6O+YIhF9Ba0eDPnehFYN7wtv1yqqbJSe6AI9trAzAVP927PjSwwBpiCIPcC6cg9KcRZhzoPLEsUM
V22hv05idror2ZVuCLAr9gn16pwWLVtbe2uQJTA1ZmIgYXCJbwL1xmELDpjJ/7kQIBuKiY7BInk4
uBtjRv5rLhYwXOJc+IgHGTWGkHUAf9r6NgqTp/zzaQVVHgSA24EcpXrBKI1w+HTIUQ8zv0fIYTMp
3Zs6kZZFNJqg3DYvInUbnKgZYKft42oHTvqjUNoQ2oQMzfApEbVQjb/1xIC5WYjI6j3I5REz5/rU
BtFeJaYsSoD2VZT7/8zUDQQ/Gb47lfnFV7UkrN/CyDsXphGnKLKbq9RSieb6Usd68up1S8QDlllX
c76g3WVVHxbdrboWpFRfCKtTR7IB/G3Eti8Nl66D2w7jIRiBTUL2nBydqnFC3vwBEpYkerXZ5J9M
7eq50bQihkgHT+uwn9wJbqc8TOq/2WnA5QXSkcZ+TjiyMRq+/JyuftZZCetdmfIXHviIlDzWYXxC
PDwnKz+HicoH9cDo4KVsqO856GO4HLSe7YcZuNFj+J+y4nIy5rtikoZQcNRsQAlUN149yvnQothg
yy0nDQLTCfGCgiOOpuOXzjbPwSz65+0vnfZ2axfYrXYuiadeFq62qUuYxcdvO9z2W+hUgaqYOwsc
QrI+DT2iFO1AhAutJxevizKLSVgsdEOPYD2iknbooOMiZjYmF6a58+W2Fn7RDjYb0PzY6YWVK2dg
Z6iXsM1DTAknasV+UBmT00TmVyAIfpKsje80P2nmffg+LuW58UtRr55GGY3RQRXAfAfoZnF1jFHE
4sKVLHR3HLjp7FBs0gmoMAeh/2yXb44sS60xHdvl18d4YxAmkAvnNIm0IFG4qK+1NeFkjZkrfgOi
6kWJMqmjdXIkyPo6ZsN+3pqJg53/gobhkWIqx/WeqXr3hNbISMykEFj6z9EktCcWevEM7/Sbjeov
/IUyp7aeU85TFKogPP2GJyPeCkYij/6CHaXmPitKFRnu0mJMuDk8bswbsCZS+QSceVJwDGlwt4Nc
H65kBlluWOMn1UUHHhaMCCFMREMxFhmGytDYEcK5F2nvjBLk+kQ56yBV0CHZSwPxYIvmEE4K2hHG
ByYYGm3RCE1vpdNvnMSos/vO30bsknWrHHNoWZt4xi32c2YZaf6M1NKy5wHqX2PztNS6bChB1R8i
mjwEQgasRGFkqYy914MmlHWaxTOSdKIkDS8krVlZBdFsbAiYZbjGdOazY0c0h8b3pVs6bOVu0+zG
x5g1ACzjhMCdEr/l71/yy+iCfrMF1zU8KwpsYJvNkbKM5cg4DKUZ6/i+EKqGGqgnanpG48+TYi8z
M831ul9ouTFwh28umsPgbyAF25FvDFAPK/kAUZog4EhDN9fqPqNVl39DaMB5sP39YXEAcnaWre6h
bsScF4Oc4ztfQRAN0inL2ljluUVDGyjiA8NMOjEGsYMFUuiZCC0Hq1LMSFqXZQMpIo6ASsfdyUa5
9rqAsRJvffILUXN2T/y2yO82IkxX3QItB6Z4ZXGa+M5s3CnEwAE4tRmDnpsUWbgsOfz4EUPJzkeI
8AwJLYhUvGDFP01449EyQjnPMTfuR5+uZmNrbK/K+pp+fW6F9UlGRpZ2t5IFJmTn2YbzFpe1u64K
qI56QfDL4YF57+Rap/JBqSIgduIhIv8tF/9ggv3xJrWN9SfY5FgJ6B3MHQIGOjo9w+/BdKTj/ys7
4mwr742wsUjdDL5qa/aL3og8uNf2jG0Qk83nvstA8ttL/2J7kTNYZuLI8NJ2L44idUS8IaIoGJQJ
voX+indzSu3/QVin0jQ1AB2iWpmZUZ2j8HnuhFzgxfA0d89fu5ausKAIHN4+RQuZUJ9NDEQjrMB9
EWX15rHsq0rmG69/hVwKLx78dEpqfE+jqVOoyZW56umS3jv+lbqcx//0Yt8b2XktdVg6u1J87KsT
Xj8fKh57kGTfYsNvz0j1255Hg7ZWW63Bd18QavuI4Z9vfb8qT5YZGt/ttvFJZdV2kpuTTfdxk72v
QHcmTafPruATGpIv6tEayvJtOkY5JZdcu/rTSNqWyRHBu8QLt9M3pG8yGbrnnV1Xg8l4F2thWjGZ
Rb3gSurK6q545jZ84LukObte6y3IhnYemdxNAmVRYQUmDkB8OUpkLfkBGpi9iIHuI71SQThUOIQK
yXzpEg0RSTssbS/ld8TRIlbe1+Ix2yfK7eK0iDzfkkgqZzo62q8dsiOTl7lM0vresdArY31lZF3J
+9bBGmMcQoJKN0ZACC7wiQKyQg/Cyob6VgUV3LNwT+Nzh2l+HaWQi051dks5jd3UCDsSl1yfj8yQ
VsXXGBLoFa3nYT3TDXG58vNN8Db0j2H09JF3T7YQ0K67JFAuJl8V+GACD5XVr56ILm6eFCMNc+U2
qeLPQ7YLuKSICkm7bjWLpiQBm4ctN2knLcNUlXFG0nE5JPBgm7c2Y93kFP6K8OHaIHstSswuIKuv
4TnqdbUUZhVnKfkQOWpXlRXP7mx2iD0ozKZ2AVVpVb1ot7W/IZhLJGJ8UtRrB4m4uqocGmioCw+m
P/MhHT8+f3gX6zicwZaP0hIk64MzNVZntqjYBqhRR1fHihyNeFoYZ8X4BueY1lHYX532hLdZnEZv
3P4SmZxjZFuPsczZVh7gSSERftgXhR2dCXfBg/fjxoQGE8oR+YYWVxOUShvmMPdPOkj8XLYxNhe0
dAWoqyd4kQnpaicRz7SGUC1/U4OXdzr2sMdlI8zLSQFGrgSgZhY3LJx8ZLmTXKfLbSYodPM/Gcsg
jPz8fwy0dR89n4SHz/PRVDIAr1fghms1QT5te/VUjWcvcTldELcFWobS2mqvub9jJdCD5pRFPcUq
4eQFHngYg6LQHQact3CMi8lWdJwXfQIKS68V/DkpF9c/G5D+Jjx+oyfoYUkMPho7uY3F6SS2X2fG
g2zxGB2lhcpgY+yvxr+cbEQSRgo3JN9uJyEdGs1fITYSAY9iecBNd/rcy8LdModdvd63qSkdr5zU
vkncSg4AWDCUFjy0+w/l9ApwqTiQ+/2Iu/7508Er76FGZNKhnMRhg4xMKxsrky/KSdSZ+1zEtZy6
l/zvGclsWLjhxf24ltWXsTpwGPpECFu/5G7+1p0Y53QzYDqBBYPAQEQnsQ7Bo2tXxioE7KhWC4gp
+5tg7s6QVKHV+6lkGN7tiDRo+shVCKERAHoa6tKqovl9lrrOIdWp1AX6qd0AuSDqI87ELahfW5Yu
li41UIDn2si8ZnrUcuFB4BQ7hChQpzmA1uXqu3s11MsYWXA6jtawK7MvtarTIGdXV2x8QCXUVv1A
l2O889S+aM4pvkXPCU8V9dQmfzJ4zrzPQ4b/N2b9y8oAZiv5loKMtpd59RUQ2MPNK+KUDAOqNsAs
qy+/ij0pwplgtThvIg4j0qDe/NMPTIFTO46f5gKkSrnUv0PR2mJ0Jmg81GQX8G443kmgD7JA58QO
YDJkru9y3I+fQsF2ETIvbVEJ2c+dGHJTGAq3wsDpS/KKnOYRVwsqBj4AF+Mtc7gf0rejizph/vyw
8ps4sIAR7Tbn57qrzSD1PKNz4f5k6ThFQCse/B3HbbcC0XGliWh1Mk357WhbyMxUibdmJ3r7H2hZ
21gC5+AHT1+MavKKLkab1jBAJ443kW3vZxURqbeZ0bJZHwqnMdjjjE9Qac985CFKK6HDqUzRvxJ7
1VkUDVzlO3i1c3aXv/09oeva35Jcw6U3/PMeUKlGvXndiPTKioX+eBX8whFFJ8Z+Fh1GX8N+KcOH
/uM7qDNl4lS1lX0dVoW0RzGOl7oYYCE46O8KN3Q2AFdbxbkCGu9Jjsz+dd7XZmfXIws+8UxzW1WY
20DMy0oSNQzNzaWhw3xvdEw3AFgaKI+ZanbQflBR2e8jbhlC6c5R8r5r1sMHZDnE00kw4vwHo7FZ
TGHbd+UdERRnOnnsBsCM0zYGz4E3qWIQp+6BCVkl9/Sv1cXVma7XpDef7+/NaxKeFEXqSi3gKh/S
J/9vYYE+MHALEo176Lr5zH+xWT8OC0f95qW1T9tTx4gfRIDfL9BrMcJy38jy1AQHSu3cOCdGCB7i
uy0biPRe75aif3nwmhWz0pkAY/GTBcknqfhWZsC2V46/v368oA3z4vyq/lzIBRvgR89AyTbp+j9x
8sNll6HTRIAy6FX8giG1HYNA5iFVEzQH2/lOIhRO7ENBrcidY/bfIsiJ7xcchuSFeZO9GKmTwnzZ
/4frDpoxF7B/KUIPDvys25VLyZPOjhVLkoVkMZN2UhtGX9ejb90WeTtlKg118F5yKSO5xDWh5C1B
+M0ehN9z/MOOFxo6ZS1IPtIwDFZh9NVD2ggdsVEGZIpvciMFbX8kI+eBMFANe/nUn0KM126i7b+j
4sVIb4J8tBGAOcfGpkxTQKaZeqptqVC9x/pHwhJef1mbtHD6943WTeJ3CDn0o9sPGMJF9pt40MwH
40qfMKxnhDbvQT7aIjn7cbUYzkl8AnZtffWLnVySjIIRuvzL/La23fFKOcwA8Gb1UIhagKbSPw2O
9OBVjYHTewn+i8vm6f/jV88MvByrUc8VyGMXiNET29ggK+e6d06noHBq7a6JhTDFe7vSKURdeEeC
kWdRef0P+q8un3S5vwJQn+Cmiv6vOlSuhXD2XkE+q2rdBX8oxxJjSYfosCCD+2wnbuToS+A+qSZS
kUyJ4VYRIJswUjkvuaKcex9iFBtosz2X15AxOxyqIXB49FcZ5H2mP1npxQEdLuV6bdQOHN81c/EC
0GW+6b9Qzkz6iQ8qJhjhag3pTOQD3ccICxDn8ckjaaDOB5UrVqDVBQMlamtC5hvw+fYwTUvzbhdm
Xh6AYO0+np77Nd/kLC0Rr/eEJ4L+zfnwUlE8UGJNBzrkTPE6iZVkr3fvCAeLOU/TVc6zqr4K3ncw
4RPn47qT1IHCtLf8hVQgJJAL+0CiUJ+e4MFh2Fo1ammGbQ3JfqaLTV48qc84qX1JFnCr1zLQwIY/
C9/34E0Qyub7aeBOjDVO9yLyA3ZQe6zLA8mcvGPI6vJrf8mmm9guxI1C+MaxW7taWD1ybrZEzlql
M3wKZZh6ZgzxhWXnRWWBiC+S3bXFIJR/kgPvygz8eqUs71uAsKv/yBmCrYU9t2UTqgXeLuSEnqyk
ne5fTWfxhIVGwywPJ6bAYqDNcTe8R4tKoBDUPBXpnZG+MxJh6V3zaBLvQGKY2nwQBccPE6JN4P+T
vyncmO3bVcE3/TN2qDQwR+n6QM2Z+Ob3EDJy4LBRu54DFXRJFrdjYgCdO1xq2y4m9wFkhslRoljp
qk4qYM1xboeXN38aWuoXA+f8h+qYVR/Gf8HIwHKqCn3w/WyPTL2q6aWFghsgPoCOMNatwePDetYI
ZJsSAZr+O32UpiaUaGB5l0vTk/WueDDAwHvhP/4WkJRd/QrEGCUD7Z4E9iDbcODzW8Y3ern7EtUZ
FBAd9Pb/sSqVfB5BBh2ulPy7p9DvIgB8pgPd1WUjxkKknY747ofTPdaprL+rftutu5O4zg0u8Xda
3CymrHHXt94/KBd4X4n1QVRDHvVG3bRxYL2hlt72kCJMqZbUNrooE3FPGBR1ezK9Gk4A4qw9L+CD
vSZW2uuazayzx4XTU4YDnTBoQvjDbbNxCF3weC7fKzoOrXcUO81XROynTqGn9uNcocMkfQ9ZQObZ
uHdOW3DotyDMHKAXQ/MTGR/sdQhLm/ik7VfEqjYpcX9Qf8sWV+bmRjWv7PC8Ty/BlFK66TbF4g2h
daDzC4N8rEi851GAkixSCHtdM1ZWkO5uX6/F+TomETe6etv3o1AQH4NnxhyVNMAvO3OTQcqaL/Wx
7VbZyPmCFzlt/Jiy/uTMoeqlIWZOKTvfiwL3Q/YEl71HH7hwmRrt60/ftTvGFUD6BtPtkoyaLNtV
ApvW1lfdJHxTVTFrq8y44bMLcmbGi4JoaOfhb0+RXSKYTxv84O+FqhuRJ/HrveCzvm+JWM59IzSl
xqTniaCNJwftjTkkEZwLC77nl0kXFIlhlBMHiPy1emEnvO/WvQECy6Z9JZz2CheVzUsXCgLZLVaG
kEEKzsdhNVnQfLNJjNuF5wN/s0wqUyYGC+aZVUyndR2fINBleiLo7CraClbimEoEFGXmrEXzX2iD
rrAwAfl5qvbv2cAZrO5m1xNLl6arYP10q+GLLG87Ee8DYrTMQLBG/39wBIHD0v0LlrsFoA2k8doB
JRPzdoWsWBSZnOQvyMyJznn+SAcfk3qZpxI1U3xowEfz6/O/DRHSFFiLwWEUwX6ihsCJV3PS/cFx
BNv7ohbbd3GlWhR/iWIOs5JfWdAxdo5HH+RLf06raw8NA2eovkukQolZkVNHyuSuxWOxWC6OKiad
OjcjXc8gdWRUJpStwEHVZEI/OMpkDDob7wwgrTLuyvPV9g6paVk+i31MU8/zvka/8YrutDtVbRoT
OWv5giS0uzhheDImKgRPcmTYizxt88zB9y1qI0lMq5vQf4OPRzrjQOI9Ed8k99/mR3vNpWO88OmG
kHjoB1BInL4RqKuduKrJvQ4dKOLEmZJ7hM40LsURCyv+HCpxnd0MEMXlUJA78aLZz0IJ6QRDaEed
iqJlQyw+8nTBRgbWMgpNmiFGFJ8OQqWWewOrGvYFQG6Nd+IlBcf67N4UE/LPvLmDcMBm4k0d6hk9
/RoDGhYzwbqQiO2iCpjG74MKgCeKRr3OT95+nIlw3zoAQdReDfqwDWZkl+8YDtJmR3kWbpmaMGtS
TcjeNgDjPiLAqiAEBAdRwgjvcF/0ijvE8+cPntZPn6G/p9sIXYwVGaIsKMGeuYxG7liMkAvTviJR
5T+LV45NQgj2Jl/CzAmgdGtSNxYbGFkylahmRX5jFjXRaxk2u53W+Sn618SzG4oHidYzr6vXwUPE
rFLomTov5csljjzLN1HEnA21H5FhAIYnd/tfiEOM/JjQqP1CNOPYR6lzBhxZoWix4NpF8sLlFk2P
a16WEByB7IOuhycPgpvRUZqIjz+fMJYt08Z80bwJDqiQ8jyMhsTJL7q+uQ2v0DAOSOr3l2h3qqtC
1DPogdJ0Edks7rctuTKRXv6v5Xvwq3hP1gcdUPkg2irfWJ/Y8z5DcMibg3QDrI/xOaWuG5zd+BvR
PqsYdaLCgWfBhuWPmPRpvsJN/ZkmEjLvOkZii3Q1RBx2tnneQak/MZXzHaj8qtkj7xsAGetarkM/
GZxQK8d2yUvLZUfEVX6FSyfFR8Tg2VIvrmKIywE8tSQyYtjzujVDiV9Q/s7piAsPwGX2CRbl4m4o
aRwfJsO7MnfDw4Ngrbo+lwvFZQWECwH7uHa+CRx55WWhjtlxbeK8iviRa70QQw7Y2MKla3qvRzXj
9qGdRNlEK+dueAd4RGow8KXmzu/V0UYaGnsaS7AEpFJJuqQDdQYYnGaTgcPR4MzVXEZ4SaMFAlQk
Pd0S6eQM/Z/Y25uQaDlpFv7iYx+PNo9EmgTH+SNTOrDoRG5kzdjPJMFaynkWldqcHIlLWf/kHvaD
CpUNe5AmGO9YYVjgOeHa35mGuvjddCINdfzxDqR6qWd17xxhCh2+6paAH273lvfGjK8hnOFqhX4j
fr6Q0pvyq8o6YZ0x22slhwP8uxfhzlZb0/tIslO6ODRE8U4ifV6idfHWiASGFfnHRa3rRGD6mqqB
xmVtqMz5lULGH7LGlirTjZ4TdtCa1fRGhqvvM1FtZez8FLjqJ9jsV5pSSYCbqH2Murh/9x9DMJsI
pD5oOfAynJsHFcMQccj7Fnl/2m1V8W9f1hNtEOk+uvUoWy64f52gNqjVehhhf8dcSR+skvsrLTGv
vYT7lbqfkb13rYubcgoIcj9ZSyj39O854qHWLzE6mwPvHxAc0oaeIObgzatCdXwXDczePvTLpe2l
W8DJgeCUHmRSXEwvTY3Jlz/mt3GI8WA7gTj0yxBrm6zbTIHv4xAxH/g5bps2HGr7EXDgfA0rojbY
LI9DpGi5TnTs0GOB2rnxOqyw889y4xl2PCHkm64LSqIAF/iKG8OFKfqIUa/7gNX9K84UdjmFrIC4
wRl+ex8xlT6wQdFhGy2TsQoXP8vjPwXMBdmBwiPKLcusEvXmfCG0g6UMag9V8Jpg6GW+lLNShZgr
a1EkyxLHa1K74EkQdEWa5hJjMI4R61Dj87dnaA51VZh5IDiqUQqsAJB9pYWLeOjTrHhWMqMg4F9U
3+on30y1iH2GE3bTBoUHS8XRxkfqwdO6xRzzzbd28b6Crre6e6t4m/LSckqW1GHBurhhEYURtlpp
gAoxVP3mBET7/kRZRXCdjKj/lXr6mN492racY58Sg0bdiFVQxVG6OpsQ6dofGGLwLfEwhnKUIfWI
SwzOg7YS/wVXygfSColNqL1jF74OUnAWWFPRQAza0APXJ+itHaIdsZ8TaEDOn4zHDj6cLT5eXsk/
zPXQmciRPipMv6LRzsHirmGDZvwYz9NQmHMj6sFvPFrzP6PbK2ZlOazvkOaeuQg42r9bAJOaIEF9
oF0Ueu+NrhJVs1JwjGQHPor1AHTP2sMwPR6LayeeaObOqClI5O1T3O29OLlRP1J+VUgfuf6Zk+mb
08J73hOby83jLpm1umqJADeoK9jl45AI68gmGwQWBes1Pu4HvAHNUz9f1bckvMgR3omchfekqSeI
mQdifuf00di3jGhStPo2P3mtXuIumPA0OjamDJdNkSjqnidOsofrxIzixfKMp6a8i8XNnGVBBL1o
Wm0BCvXrzIDgWT4ciydqEElpC2ezW6rbKwhVRXeY3yKcN57FSnXcnmJNV9WBcMxuJhkW3xaKTGgb
wOb7rQCvwI4Wtao4mlzq/Z9NUdudGy7h9m8IjM66UngpjRzm2Do5ETsMbEY2EsW7wWfaebnhyhLa
0j3eIrtcX7UMXtc3V6HVTEw8vr3GBffk7sIU2iCdGupOhxgISvWexnPECZpcojRIHuVmvidDfthI
VwiqsxCpEECkR9zddd7PjBmrkNYl7rWheySjhkLncjEhZGLUtArGnoFhlLUr8fQ7j7/+RSFQXcgx
6t8b0tv998ePZw9MQy2w2uNRKwf07XWYAaqR/pQP2JJxiobYfNnZ+huOQkfvnQMIZYi5+TOoZ0/U
MxtJZr2yO3uUNxe7QWfpSYkLYE/zbEGlPafr+8oO4YfdtHjX1DWNPxJ20K2LO0T3BRbAXae7G6m9
GeqFFpms8n02jvbjfoEUgaeiwFO52bkml9NPEzdi7KDl6yvHIc1BgN6CTEQekyY+S7HWslOmnpwh
m+KSQaAfNC77jOyVrZ7XSjkOX15N4CKloKXHs+npJmYtqMbeuRIVELPD7nLEsaKE5Wvlea+iRfIq
bw3gMJ9qCs7kJyFO/K/Xe2P0wWHE/Y78u6/b962cmMA+x2FCED2XCIK9gMdxxTYrtQrNx9q0knPY
PlTwfOBJUfYm5V8N0rO+60gWBFvnsowdN/wbLQ9erD9B19Nx6q6W7q5mvHzZug+tGUuCLb8AvtUe
ykkJIdzkWyn9YC9p9LY1f3th2fmsdRLiu96RjR4iAOdeZX27n0Hc5ZSRSBs4Yu5IUBp1ZsxJhR7L
thf3An+ht+bdY+e6kYd2wLTPr8n7864fxHblzmBVjTEH3QHvmKOR1tLfBXGmgCz9da/tLxIVROEG
+TaAmNtUkD1F5ZY41YXIzsgEHix+NCArLpiOA0WspCkox/ATem7LuAeT2C1SOQ4LjUNqlEyWZsG8
SquLoKgZ7o9/yXMbYKFf0+C3XuyCBMviMEsAU4NaKmBhAj+i7pOrOSc3D8E4J+dx8273IMPMYnf0
Q+7i5odzlWQsfHyY8G23PYrGmVpRmsJWafyibmGhJQei+flitcei8eXknaLfi6yYlVKhyH58EJfG
dpG985DT38vw9fn+XxGjrLxn2D5WCdOuBerBvGIBBkO+qW5Gwo3XnulMrlAaVAcvyWGFDWEBIzOd
h0uEhz6TjQIP3uQfEydAfcs7l+bPMMwZS4Yf4Fe0LEOIeBPfU8DKvvSNShItpQpHCe9BMfJ1DsOi
xZZPg1U8+6lwevtQQtxeUSeFEsAizSBJuEyqOy8X3hs8s9BUIxncCZU4JzKbWWkWBGxC2eYqwNv9
cvwRdx/6Th6Z3XW14QJdXIcEUmBGZ2djLieQRWGeIvO6eZ3k78a7t4LKx8BEUSZ9IYYvuF9Jkqx5
2FI9TD9n78g6ECSzRUFM9Cn+EHcx1hltnODVtAwffRr1z+Qp5iI1I5CKt8dwhg85soo25Zyzr5A/
00Fe0bYcnxEGbqshswt9stABvwa8mV9BoDCJRwbEJW7Hwl8c+J78MajujIXzOB3PG05b7W+eYsUh
rN60sb9OVmEHYODVySGJxAGE2FquxfHG5fdVgFEdzGA+A044iM8Y0yPDdDtc5xMhTAHvNHKxKR1P
gUaKSKAZ/1PijJouYoBkqXbkHUHQAaU/BmAbjTtzNmXtxZC/iFSSH+JxWVW2RvrkRbA+A/7WUeeo
9EJslufTYeS9n6niM8DT4R4JHH84srjLmdTGIQfDU9Uek6FIxjMlpFZCMNVvi8MiUPMK46+hJzHn
tur8oOHTi1GA46QR0uc1vAAfAkpfvQ/tbL8zMEPJhlZmfZ3oGVtgiLAp8EDvsssw5YMKax6O/ZUZ
mTugk/8gu5reat6q5Q/4nbP4+kvIcUEtato1tqxJxHufqC8j2lB+GX7zLluOMW/1V7Jd7rCWzZwI
nhlwvzAi+U+Sm8RTYq3sZbUi6HssnxkBJUxxsL/zIee1l87YOzThrxDmeoH8YMbDRuIrNro17I1e
6hYe8i1Br6wAYcc0WLOnHWvxrh4uSI+HFOwuFm3aOLb3/vQTQGDJDde1P2G+7rtPnnHyTwYxW2hj
lxL0tdyG343jwlvoxWzsX+rE3Y2jcUCZl8tIHLxmdV4zBBNmUnImUrfjo7nZTLZMhGO3XUDzz1GH
giWa7uFYSykFo23cDHsPtu2ooFivYHxDTp1JJW8PK5/Xm/+yAMxnI8bGSgzoq5Op17cz9g4XnrwB
Sy9hS7gnDXey8sQXIENgwtNQu6Kh0j4YGrSg1xGiJ5+GWZhmIqJgP6zAJj1D1h5Q3xO9Vd6cID5E
SCfu/4iQKyz23YTFdgidA1JmKXEjSBsjn/7CQ0eQhCZo2TgPXM13BicQqn1U747TbK0wrsDaCl7w
92UJDiw1otrQuV3EkgkynsmAdAjCT8KyRqOqZsax8htnutL9D8pzmCWOw8yhPXFvHcUG8hIi4q3O
yqwoh9KccsNqWxlJanXh2Z8byl65uq4NZf8uLT/EiAbe1PSrFTe163/kQE8777123la9j4ayeg29
9EqOoyOV4dHvYJ07J45MO9OEVAUopjj2Td77EiUu6a4tLxNX3NgihSWCaxOtHCSHjUiMW6z3YslC
TVNnYIRvS+0qFshHwBL2kjzGqHXVQIiDmbEm5Yn/tO5K5NnrMW5q+lJNg5MA8gOiRQcxoI64EbN7
2lrYsKqc4+S0d4k+e2XpkVEPQavyMERmG1ED5SrmCTxwcVZuy64EyAiU0Kd4JjqntKsL/vnZOjk1
1qsiX6rdYKKMPAPgHPGJ2BQXc3c3n6bYvxtBtsGgVCjjw5gLzKGNaSJCHeBL9Llae9vfPxdVeS1a
gKqHLmuTYI4w8ZP50MSW7dnEI6YZwdF1k+zZn6/8/b6YgeZtuZyM/L+UmkunVbEpwdKlJ12JgB3P
ZAzGxMV0yCC2SLJPNN5xsdOWRvzXNKfHa3unNln0XAbmGO3WDt5zEUjA+P/tsDmmSq9urOIgL8kR
a/uqoV4qWYPSRBKoADlnYnUt+APQNU1BF43+Jxl6avSibGAm3PgX+hvcd1lmrEPF1PS5pqDaXVzM
MlICaPLl7tVijvmQGztn18KKjauX7LdddPkoMOQvsDawHaMiPwUdyx+LmvnTseoq+hzEbbhzLQ1m
xX0ZJiAkyHdri5BZRJuWRbS/+OaqHmNKYSbZrIG6xxnB2anvczUBPVGTcWOTYzAsFB+r6ThNd/uI
vYskSr0FRhlnseoAr5R/TNIjQTAt40Ou/k/0IojVjmuYwiHK6C4bi1DcgTsVPBAD+ysXlsR3XESr
7qBZwcFLklkvNqmRo/MPurxe0bytum3lYGSo5dyUdjk5QaYuymdP/svHSobf2IG2zcy86qf+IyGl
xcAqIXHhmF0TF/p5l1UKjRcvfty0/gXp1dl5iaddS6SrhsUPSNR6KSse7LDZykIz5emzeR4xYENi
hAZDEsLQk4JcaWdfeNsvcm54+6Wl8aCdn2VNbWhUWVl68Gf6T/q2l3hhUgFu1ixI4649IdCtAYH2
f+yEr3rV9Q25JpTCsxZlqVb5LnNVJct6olY8A6ZsjKGeFqZvsSkzbRccHMBl09RS+6JE34BrPF1X
Ps6G6ix9gDl3unfEFu/OywbFyPouSKO1FjUrG35i6q2YzLNjCuxv3AGcnWkkK0ir820Rr4i2Q6ym
VL5L+A0BMGgj1CIYZhmdQMvVcswmL4KN+9Dpo7gcpXDNc5wHdLFKrehrymX7SKL7HQjDStzcES19
JOOv/jSPH57tcLOrsvTQYwAJXEkTYK2pZwsuATfIIQCki1Eev4vYAajQWfnylRZeAiUXXqi/oYhC
5HC8X9QXNztjn+B92yzP0TZpyEWDKRs1QmUBy5no0C+Fq+ucOPlC/HvnORVVfQhGYtsCGCQYSChz
wmJ1rdWMSOLB/OkiYIXOHv0y2CfOPTbbnJtsAMAzuXJ9GxbUe/a9zcrCmH1aiYLaJ8+cdcxJ7M7y
VzGIEervi1wy3rJPK41WkzmW7y1G6LJdjQICkJxax7Jk8t6vrBf27CDRm9XUGN0uAscppJTOfD6u
j5DctQ9xYATTtLKOXipsrFpD/Tdt00X+oXuw3easz8Meh5yO8RMQBG+Fsts2sXjXMgAm716+kYF8
cwnof2zHrWQhy0fqglW1RFNM4S06RmGN7ss+H+l+85rpATYWLOvYdmRMQn6671InZO7AHaAfiiLb
qzbTNFe/oBPKGS/VkR8UTDvL166VIKccUOVuzxJs6WJCzpOwnTAd0cRpk6ihf4uiy5VJq4GGNhq+
fFW0OcoPGdumN+O3CWYI+PkupeCB2ND663dewwcunkUQpGfIPwvMZjeXWiCJLq5KAHzKFzRmv2gQ
lsCVh3SHVtJ0BVWf0iIAsZNFFwRO9elp0hsSyVNyMrY8c7SYrvtNFwAgePgTsQK/urjOBNhj8uPI
qig2GlkiLbzi+l1aqmXzgiCEW57QPpCmtpOCfqSvSSsGKlj9ecUeDe1JN0ekktNa7vm6rUINA9qM
VSLeudzm0r4iM48RSTDV6S5XV7OQJnrX7oiypgEYuJs7ZuwdY7ODr7v6TbasB0u5ima80FkZjfU5
5REEVZZS6zu2dSpZ0fB8hQArF4e1iwa/TBXSYqynArKATjjVUclvInJjopvx/mzK0f95BkCrzW8k
HpQYsWOv0KlJ47c7cj2Iq0Cp3jXalyrlErynaQ4vqve4N8Ycdmmb9aXYTByufAtSe4jZ1d0jDVcz
HY4OPrjXIsgzc+v7chSDuFoqWCetuLP/g70pxBEeV6ihNDiq5S/BtZbURpaLiVb8qfQGvENxeIil
qbL+4ufw4KwjNhKLsXJbR5ZbFllDKuyMVoRucshops34DL0C7zWVIqxvuxrskjvrAYOraL68jy3z
LaPfDgle06zfT3A6+eA/UIbhs5e50jIOqM8PeXyMi7d2rA14hgit8V8akD0VJ0EfeHViH705l6Hu
OCO2xsEX1Nlb5AaEjmxjw7hFcVwzpzTdwjJZb1IR9LScflOqAu2MWlGGOHaaaJjr+AGc28wBb3qs
DlNNvFUOh2BIKV6CgizI2UgJdKCwN+7M+2BIO4aFU8kOT2Nnss4Ot9E7s/+7IfMTSpEXtmbNwOcV
b+g3/Os8PyW/b6oB4t5pXLT0b928N7aGC5XEIfPEeA6eHKXvvhblS5a0weARxTybehITkP7Tu/CR
i0NY01fe8KCla9xZMYO66cCz4EqRD6Dll7XB5ZuDmslzeze29fn3I0XxBgN4vivufDEkh1AsjP7J
HdaXNbgtrGPJo5mAPLMB15EyIXzkHxb798octefWEsKhhrAls0pLqgIoNGXy0jfrOC2ZDJ32SuBl
uWBcGq3pJWaJf6F5wRkKm/wvOaCrev/a7Kj6EY+X8+UgJd88yXi42+Ixa7hrz9TEc68Q+lpOLp0k
E76w3W+uyWnJZ7UY5X2kX2PlUkEREJ8MEKjwnOZUlp9Kzd53Czo9mUO37jOwdhkHLDecmY+vLynl
ugnCVcLvC+gY9TVo54xjbgjFqorYKkGHst562YYXJvQ8R5ZeJHIxB/frlpLXd+XG9wlL0cGadOfn
FYnFlb0f458zo2Mv/c433+tYzX5PF6aPIrBJbOyFZkMaiA/6G3Lqjz4tRgEM/o66fxf6hyicn9Un
VAsCOMw2PJLt8jpIDl5hkPymUZy3+0eecoFNozBWnapQ7NrE5Kc1cD5paIugoWH5zmyf5U/Vp/D9
ICKfZtConKbz4Yp22105S32PTYIISeMHNNAHnA7XTDCYm8VgT53Ev0mOGKicbuvPD8tgq4uvvpWI
X0Un2KL92CwAZO28XdDof02Y4iguF0lb4K15ILa7ExlBbf9xlgfHNAJRiYtC6Oo/YegXIowTH0dW
3CGwzP5qH71PyFTO6YL1WbYHvxVSBa/QjMiGzmGo9eflaRjhmy3d2kqNZUEY4brcI4l2ywL8CgQX
SumXeFT77jbF7fS31iKfY4E66hTMZWEZMkBbnJ+dVRCNcvUJhqZP0QYl+5PRk1qQviYx4WXf+6VZ
3wL37/15IHb6cYpnUBQ4VzCnWqbNlxEWLX7X9utAqoH2qSUzEW8PyIebB7BrLxAyoxOLu8827xji
IOvhlfMXDG30XS5i0K9aBoo1AVD97tlpzmVjwCZnpBVbGe4+AZ4PZqGsGw0WZPCrWAoRLW3Zdqpa
40buvOBJPLoNv188arKVz3Mci4mCBaMDSY9Tf7+m5gZXeAkE7Do9Wtb/I/WR4nHKDmolDith6lM/
rJTWuJP+36YaWI14muXpyf8Gq87fEmHrFgjp+AQuE3r8Gx+O1L8KpznHiGhSVeWKyhUTwTGw35TI
Xy5hbzpVzxaXqWCjAt2rCyNisZpTSyFkjaLTtPy1qhNHFLcFNdF0xnU5jRAJ11PPuO9i+UXCrids
p02LQA4aBuHrYDwkfenPH9xnGl3wG3h08wPgysOrMNvTPGMbteL/igmWkT8lSe3tO29e/KJ3nr1r
/hGuyqMh4bEqecZuWBNAUmgy9i2bXqqjhNG05DTi1ysljzK1UyyLe4PEv9uu/CE8WiiUkExdRf1G
kA0OADqm/IWSZdaMNe1CZ75jHHZsd2N0N1SDdanqit0sp50XOoqBBGLq7rHXGgg9xolkYkMi+BNs
74O2ASYH5xzP5oF2IYDuDeF/WzuPC523fKaICuGqeNbvMOzOMmwzWe15U1meY6Gir4PbhcAMWqOY
PWnoFdVMIG8Ua/c8Vh9Std7e4aLCqwoaqq0Kg7kkot38d8RYCSSqUBuuQjd+kCh7d9HfVPXVc+RX
7dvpgSqGkYKFntKD2rSoABpIcBiViZYGUrNJaggkZPOrpAz+eEL+G1tG9WTDiPtJK0qLLXCX++Aq
AuKyBNvHMUazr394B2B83Gun2WZpcCqflkfuU8xOCrZ8jsbDzQ5BwuL9zJBAk/DdCL3fmMizn3eF
gLMnz193IAeL4OEmdnMMIVaeJoml8q0uFDx747buAs2pXGbmB/Sd+m1fMvEiNLDKDwbAzMhXH4Kb
yGGB431NFGU5boJ6oXcqK6Wi52r+TdmVyWiurTa8E3/QnpimH0BG+S7GIwXbI4bWqXaX7ewKMpGo
Cgvo0y5vtGxIgSYrEmyTWb1gcSP+mEqQB8iFw8kRN09/OSrFGDAVUoi5prewJvZRc4Ik9MKVPn8E
s1n9rRvCRfs7u3ok2yiTq8wdtiYcGdbhgppUUgz9N1XlBuC35SmZ2xvtl+j9nqezDXeE8uG7fv7S
XaDQmLx3YuGHNSPRjmXejef8GukM6G7lCuU2gjMIdITXkulChGJNMFhgdq1F7uyomQd2H/pt81re
VljAYd4f8fA6BDAqKtNDu0tyNAenr3qaRuYEtLdYarY0IKyg6RtOnJU3xQK183sNxGYaIaVz35YT
J4OD1wvf/ebDmxbXaSOGpLJfNVudeF+xGRyFg8xR67vnHwnBYqhURm+34tB0HqzGTNJ0vSZ2zu9X
boYBTGFPFA7DD2O40g6ENn1PRV0QcdHfq74VpvZ867K8WQjpTR2FixsErCV8rgyt5Kg6AOm8Vy8r
fGvI5fbV8tFa2shm4N1Kcm9EWaOB6IspFXisds/ZR9CPR+xQSn5AxWeIRS1QlYEz2NKkfx9cIl3n
7kDLxVBQv0QE6cZkNzVztPbmv9hsT+en27/UKx02xTbK83JQm1JnsYNWb8C7tQjptsGr6D5KoRSU
KNAxVYLdNvRMTTD9Ceae2NwhEn1oXKVG7g8qjJA7k83EYPhNKXoEcaGReuBQXeTnFsCv6P6rnoAA
swCFlSoxOlE6grejlB55AIDrrxtx6rV672FoLH0k/g1QrdaRQT9mCZ+JS8FXcUqh9KkMxD7BHKuH
neplQB+RGh4wgt8Zp4A/iTbb+jeqt+SiMt6KQ0aLKxwi9AmK7xPFMXV+4FMcBJbCCb6eFk6RHuNV
UAfsi6+rCuFYAYaMAJiNcMUZLPT7CGrz6TrM/1Dzwm7EoyyRY7Ya23yKq2o1BM8/VtDf2iqJp7Am
bVCfL8iGumXilJJHOb3RkLuo6GEWG4FcKggFqSxt6gCpnDlewQ/gvDtFVF+jlo1vv4hFtx6n0s19
9cy+DOFfv2FI26CGIL4Q/sDeAYIQ5FPxZYPsmfmEL1zNwXbH3Fug0KqjriXVESQGVs6Ey22PzQFn
cr8k5xRfAadktttOGWNyW7BP1cLUWyVP3vH2W7pMmYUz+ZDcuXjMsB8EtPldEO+uKcDjjopRQb9s
6tZfkaBQKDZMQcdtZHgXZ1hSdUq4eYkmeBbA6EfDoCfcRFp9nKIb/QMgk4SBNYHE8IqfG7UCUMGq
sOisiCmMMH/FEd3EMW4F4Q/0B8n2N89kd7jtNg/t/XOJ3in+dtY23aXcPuxDQA8G1mlTCYhbBL4t
FMHP79mTW7DBiNnNZnDiwvViZyVATkV1dran0RSiBQTDmiPJfW/5RX/Zt/cfk86dhXIvYoqXh/A6
y+dvz3v7TuttAdFfFoT3v/I3H3FyAs2/ixeUmk5Km6epRJXRL2VtWzlvaa2s+U73TkpeVSgTRJ6+
MFDiNrCP6Z/i7EE4UB149AE40Q0Xkd8EVuNqn9iwCQIXi3fp/UOVDH3fJ/DVnrIEGivp+0rU7Ujj
W7DRUhhUF56o7S3H6ehb69fYXjmRGHbLh3TRPQUd8wtjhwQegc9c6N82bt5s0eQT1AjUsnMvpP5z
eZQ+6jD0x9WVqwTQc1sRuqQt4NfvRknD0DJaP38AJVGYIrDfHvXQEmhedAQXDGwv8hkEfF0hBELU
POY0GStEp8+pCXN7F2gCGh8p+vTOfrYUt/VStyT2taDhdQ/EuiJKGwM7dVbY7hQUrE91b/PlCVZq
dmeCxboZ+Iu/f8FIxO5ocBgrfpYQO+nF6xt9fyKefsUhgMAS51/7HBun2jcVE/srexCh0c2CV/+a
IFkztQcygkL7qAeKbqHohOnmSlium3fqfpR6daaL436fs8JbmnLG4tHkGZPvmfoEQQeHYdbm1ILR
l1Wbj7jF98X+5l3Imm5qo5vQXBk/OjQ6DxzLJ1HcxfS5idqdof8yMMtzIdvhCQDQ4yxgIkpI31Lj
pvO3olbiwSsmKwYmqQyoRM1EuCZlNLFIEarF/DtTf/xMB7ALhe34dY503AyDfULOdc4VZoDB1zqV
J9k578oMekr5MqRIBfR2huvk8CoY+yfQc8UMrZiR5jsHDgJaKohN3TUUk0dmOXokQ4SVMIlVYq1N
Xsm+AsgSJ1xnJpNrBqRtA7A9hsUVZemgSlZI51YyRE5ZNJCcWfzD2vKNGLXpJ9TxkR/1U246TGwD
Jn1n4gTJcVP0uDxkJ6+n5DYvv0KOaHdJUlwRScdYMht4pWKulzRECk5kiai7IJM4NI9TkxXEFjNR
KE+YHUFuQc+n6U217lNGlOewQzEqP2ZP3lE3Cl76cSmxwdGyfUNl3UujhvS0RTgqm+5wTOegHQ2g
A7hdetYav1I2FjndjvJLjLQ2gzK89oYGorvsWUOMcD6Q0EoTI7HPB4q+ZFS9m4i4A9MZwOvNhqg9
W7VED5imOuUzEk8giK2X5TEqlSkDke3mTqMN/AlD9Cu2ViklCyIBrL2+EmJl5i7bM2Xyr72+OBft
qjXxJv9Ls2KIUOXiXZZ2udAs40/4y8Ap1yWKLiCUU84iVUtIeIhbm+2wfWddkeTPXFPDkZ2EMn6H
WZno97cdHmXUAA4O+s0TGf82yMb9z1n9fQxKtiF/Vf44MRqfjrdSMCjy2W1BciEQ9ext1vf0/8OR
jD0Z08W1HzVGBn/fLEAWHkGg/72fZIX+Kw7o3dnavv6ARAISBAbhpbqZdileCwozF/XeQGeLsYpB
Ue0g1Q0FAM3PZX0ijPw8WJ9kG88GW6d2CzhpqSrzDN0ye2vMcz58vJflza/oXbjwSTDIuStD7Dsb
Sx+iSXQ8ZujTT8pPXjNWZ5NDdesBYcoFx3/THPES9QPLvu8ggyn4aE7lkd4abyZHiXpNcfdRmPNM
/XlbKoncRC95FpVlA3eswxz4hQn/ON0TtcICiULEF1d+0gi+JJSrhZpON/fA/sFyUxPglwRkH7D9
fnOleMSkgFNFiySi5ucIcV6WEczGpDzxhHYYY7Xom0oFA09DH84+6uMqxg7XGv/2PrKkidayvCJq
Sbu46Ft0bD+rpHqDdRPeWkkS7CoNenXXaCMgHGcooX5GCdFeUuovQlkysjpfK4286ZN/x6Xhc4QN
yRccekTHlgvJMdokv4JRlGZP/L1rIPKgJm7NA2C48OcDmlewru7E3SkqTxRdRYC7XWfBnmYh58t6
pLsskh/oKoga5TeKcQ6TVs4kkLvegH9Lu109IFYdbnkHH6HbuGV79J9eSkpnQRiJ+GSNNNZp6L21
vQHaQnEo0ybWQPlImoSgsHkfKqbr2V6+MDhmCoZI49vdJVDKKg3FcD7ZZy0vsD1/UauDDjxjVQLe
Ao+VViX+emWpuNiAkjTHeqipqcZcqpAhXhCwWBVlEz0+qBbF3J4MpT6gBkK0KKfT5qZoK2fDtHta
PmROAx9z0YiomXHwGJZpl8gNj3TGnLq4dKzv3ey3F+4CG5rylfzKtPkffyMpawKLOoTFAFX3SdwI
8bhSZeGFm+L058u4EBoMmjS1Yk6hyyQqdOnFXNChEc9OXEk5bdloT5DAVR0Jh74zw0/tUnglSAuP
10p2ozIcySrmHOm42SJUIKrl8a507QxSVpvqm7pjS3EqXVPElqxRWOdnH+Bgr+0fWTIu0DdOIDkv
rlbNSF/1WNoRJCESApGtrYfzBrPgiSbN6wSBk4NHBM55Y+sqX1gTNwWohn3CiyWB5cHaBpBM25Ic
j2fCOq6sdK1xp0KGtU6Ij8mSkqzzWqM/jx+MNwlYTIVYfxAaKsQBLPMGiAz09JWd/rjbjm8uVsKb
0+kAlEDHQ0RIiqZUQBv+tsju40J0FzlPa1lY5oam+YRTSOmcHPQzLXmMWTsHXTxnZ5t2fF1sgF3+
wR1DLkhLaeWzAHxfsnxerOCw1EGEthGdNdunjq55KcE4QOVo98GLiTlUVHbVfxfyBSBv1IQBo8Dn
tyGIDhwpVQjVWEtbu7XSbW6E3VTQSGtMwBwyWeuqaiCXGHqsHwf3LnA2YtQluJZ4qVGvz+3CH8rJ
HG1Uot39eoKXvllUaNh9ig+kQ6uaV6+eqv9LM2V4vBbzX0yuWG/sjNFX2KhSbsHAxy/yiTWpXJKu
PT1Ecc4y+eXU1n9Gj/SFbZQg7sRDT7v553qaHyJsIhKV9fEjmLQm//g0WUkDvoekx4VHqDONnYLP
4KXrWXKeL7RFZKZMZzOt6zkdT2UkE+EGZbQNWxnt07vY1Pf1n0w+Tb6CqvE0/RqVqNR9Unk3SgSZ
jJtu+dWtBu3Y1JeYXC+5tz9NVDTiGa+NKguMjd/aYV7XwOtf8LUObsBZCMgboztPvmaNyopwXi4+
oq4xjnbBkhN2UaitgXypUc0YRd5k7irevDERs3+X4wM1YYXJsUNrxnTQrba6VjFZ2n3iClLyaAwc
+fqqLoh3XVO7m8mpL8dhmNYiVWONeHpdVAIrmQagGFWa5WqahoySTZKcznTvekXqKMQKIzIbIPxg
LmFGGdK/PLhoHmrrG+GyyKYviDFljvQk3J5I874q1OGlxUq31n/1mCDVmAtar/pmYDIv/n0BdOAp
5knqSd5moHHNjGVXHw6G63vw5EviRQpBTd8AhrkbpuPg2UHjzUWHRLnRoRBVNwmUN2sOOAl04PdE
Eb1PnOLVlNf3+7nxztD1lvQeCqQ9ISVhlQODE+4xS5BWDMTkpdMrLv/4Tod/ocOG8HakggnPfFAo
2e+bM5VAwgnLx2ga0w1EF2WBuZ5Yv8HbvIlzaQucQqKtMoQv/TKTq4zCEfYHjNIV5pZ1RGtoQdg+
Rj3P7ja8UVtJ+UfgBvtYErTlDub4fDtPNHrbzMN/MAav0GGyoynmEPpm4Wea8mXtBkW1DqlhAEq9
mOt0UGIRQxcO/V/G+SVr6voKSCxTtk46mJ2V+5S0iVmPjZvBGyXyZiKkrlEO3QZAJ0jSrSMlcxs9
CYS1QXrA8ohOycy9h0uF9JI04/cSNEORRGnQpdyGbiEzJdfWcgzrwzm4fmaXZAYIBZ9uUEOxHERJ
7mRzGKybjKqyJlsIsToyxzslQ1XNs3GAkQR1L6hxk3dedZY3veIycIOhtSBH0vIjabCsfcALHO+i
eI2bNdsZcMNbYI/I2J8c8gGMUaymRPdPdPmzJdRq83aztwB3Nj7jlFqXhRByXik0YFaw1OStI9wW
TG3k7VVudyKzWySaJB3MshuHr7Z4G+uSc//nExOAYkJGz5TuTNcK0UENf0kbzS6FnVRfSjzmogob
rY6zUJNPhELk98hBQ0B98yXwER0/KL9z/mGhd/Y96v0N3oSyHUcrJRjwodIbhaRy3C+mXQHlAWHV
HRsJyzCXSNUJVK6wQ53L8dtQxJ+S+tGB2K9m+UHFmxSBxZah8uW1qWLkLbGH7MaK/6/wp0RUlNlb
sB4moJxBL9aMggGxeOwViXcDaqg40JQkzqsOlXRwvjPIu6Kln53G6FXExa5HCniM8rwPC7HZNZbs
+RIG3Vs5s/EKZ4qNR0tXNYMC7laxnxzIfmmoOKngp6ibG7isUx7S3bYoNGeqG/UevdUgXQwxCWUP
6CWfRlHKVQzVJiNjOzqNhGTZJdfxDCvbPhfSUcDJfI29Fdzi1i6+CDd3kEXDitJUhgo4HZuLIUFE
k4xB7vxHki0UXyBUMDnBmoaw/U3OSPUYC11GXYYbDOXgMMVmgw9JgAjv4sXuXExYer7KLoqGIej0
meExoqbM5Z6NZIcf/GXxlerUSucOw0sYTq4yjfBkT5yq+o0VENFdt9/3KZFrMKoy2J9v556SI3pW
GrqoiPXa5FmTiB71+dYsSKnSLnaAhTFBFpZsxZ2V/5hAXdhtzFxsxuZ+Mk2uxtebELu8hFq+mzuu
ZteJBXCkPkIa8lgPeVGiT+Yol8Uqtsmf8EqdJ8Dsw9gBOUg442hx3WEmMGPzdl1sukP6/qPMn87/
g0byjTP7K2RqyukDDrGxZN3nCk7YYtHlsNnprLCTKTBYYwcXaamVPp49qs1/AG6x6iRlBBQ3l44F
19VV20oh9evZa8YGmUuLXDscHkc8mrY5EMYiReURKA/mHR7j6gFxz4nmm9/cqf/RMHk/5Qn5h+M1
ekS5qQndcODXjwjkKdJ5a6xHug6fL2kUQwIwuztWy/Pg51pXhR/8+Q9jNYVp2WwWkYu4Ba2lCMTT
6lyvUwa3iGY5T0YBF8Nr7hNkptJpuQ6ZeV66VYVjAnIrmeIZ3oAMKg5ChHcNiUOcNobJAZKa/O1i
T4l5crIX3vF8HQAQyRsgXF1CPPIxTMV7KtIsYsYoL3lUIi/p7Bq6PR+Pl51mW0hh+VEumN+QXHbR
VGtjbSrPnIh1z6VmvKsIP1qkPuzBJcbiAcFihY6Wmc/bf74cqCiyNjsgO3+IlDXj4oM6Ty6BwQRl
yGYx0S6U4gP432hcwmhhBioehWLkzufxs7kRTrRuNNV+X9+vSd6xDjMGIBR1oECENZHDCUcKfrPG
JWijbZ8GMEWnvXKc8uDRJ98Pa5eezl18ibc7NcdzXPPQNETghBA5w5mDKy8afY2w4FbNW7XCdcDK
nhLqMZWM7hqy6zzvBBawaLomJM0LAWtHjc7X6wtw1qR8jdw3ScBfMDXQrriAgvCcE/R9MDu6gBa8
isCctucrCZ2a5fVCgpn9BGyn3DoxP4wp777lM0un9ZzUTZsk9ecLCvLxOxOxBGuAxjd7fKtiVVLQ
eVZmoVEo3fozc1m2KZJkOtcVaL69cQo1XuaqkMVd6EX5dsIxJUiLGz7HKYbsL72kXtmPpCVlwHeq
5h/+QrUm9EvTFjzNY90cQdycSsdb6R0EVmPEz/q+Zqyqm3KxErBw4nJ3lHiOKp2bEGDnBpXasHJC
7MKGZgkqzgUfQ19DNln6SSAlrMHQ8XTfbe0/ojIAgK9cU2weFoGg9RMFrq02DJ6QolAy49cyuvnP
I1aqPXosXmCNsBLbd6I/Z4jwBipzsnZDH+yF/1TMLHZDnmI9utkdIexNksttJ/CVLrCE2ngdCeKO
ozgvMlOueC8a1nQ1KjTT6jys+68+w1sDeYXg8Btt2JIQrIwZ2lktUxMmOIQNQd5WnuVpT9fQpzUY
rIbkXj3nasVFpWlmyCkzo/WTp36O3Z5vSk8MTnqnX1SbIt88djnFFnq3ZiOYWzaUm7HSDOm5Sci0
3UJgR9CWpt+r5oHmMGdodZOImkPw+GS0e+WQnJ1xqy9vfZAED6pELyOUyU6Wf26dzJsPrFIOJ3Qb
T95w3pfIaner0gn+ecl188LYpZbvaWzjaTjUJwUkjw3ZqBX9ZeZOvEOoq9xQIlXfRq573QBetqUR
aBBnIacc0yzgD9vk6hMnpUGMVO9OWThI0pcJDFho/MCR/qYSpp3evzeS9KEJVHmEVkyl7Trtu32q
uGOFBQqzUsAePDpNmlZwwBKne7C7ON8JYmeBjj2ue9JALde8KQmnrv158Wpwp4uxn1mOhgy2TW8u
ShSPmno9eNNkpCiglwp4YeP+zi/jnrGQXuEIifBNgoFpSijHOx+XNg7ZBy77tC56FdSmKyYTsRy8
qJ8DyorQqxbRoy1skTlfXzTQYmtRTkIUif0lwBhREWKYjqTh/piDCUor0X/P6WnRt6m2Jyw2qp8q
TRE5MxiQ2GRJXwYLqbgwpEwif0anjgaiLSERT6GyAmRim3JngcHwwZMVn22eLH1TfitQo/F8Y51P
WT55jwkpih26SVxrNpn4jd2eYdtJMWyusb+cfDm4i07+h2BmKm4Z5j91WsoFRdT3WTZHauAyAT48
ow36CNL4ObsljxMkR9gU+oEPN1luDAl9+DywikbsUccGzITrziMqB3CeVl/XWp+LmzJ0dcO/TWcO
10xOM1tMNQgP3gNFIyWJJzX+wo8k/jvMuWSyY8OUumY6uaglPL36xhIbGZiwvTlgZhBYSY/69J1h
f2hZL0arQWffu2V2GhwKitxJnrFkeTJvIeDlBJko7jIVrj+XCIeeNSuvYt5TuCAtuIoO6Gpb3p3n
4XOK1tPUwxsXUf3aVTuOKjCfKmu6iZH9XLB14Mm4rTL/vGroW3iQMvFJTVrOZjK+wNnegFuTe3HB
WTu2kdABrhXwhHb0Z2XzP4N6H1GMmTf7ZnIPnL/EfWZzx6vE2qW0zQ0aN8GwkRshAZ65AW0rPnRb
azt1QV/hIugpwobfyPKMNqwDRpZlcKd9E1RorvE4aBKi+ihht1O+WH7SvfVOU5T8blPPM3/3Jc3p
Qq1iVLOA0sWbQIcnMZI7ke28JzBHMUTbydzQP0ADGvWPAigVOLrwaY+kqD5hSc9p7Jy1J6dfB4PD
oLU5srlnapPEEkDmPh1MPm1ngfE4IOvNzINH5OouKNM8zUKT63B3I1UtlwcRLh2dL44rDHEA/xir
xhKKa041RUSYP44YZQx64FnwbK1ERYK130Tvv8bDYEqKDsweQrm1mpYMdHc0jML6bzeorTDFMoPL
2fge0xp6Apa68F1Wku+LLOH3P0L0Sa6eNhTBmAktAne8zlRxn5k6nmWDQlppxLZSNLGlC1vC9fAy
D7Gsdt9DQxAxOV1OG1UFiX/rmjXbvctjGp4Kw+YsvzYYKCr92dy4ENwUg58AOoBqoh79pPfKjKtD
sTt2qTKQV/l6W/R3VW/AMwrnLIHTjpKc0arBBEnDj3/1vInrLKyXryWS8tk5PvdMWdfSZE5ETvQ/
vb+//D9SiaToGk1Hq7zhiht1T0o4GCsFV/Kf9lSy1NvXtG4U4W4OT/259yIt6LayMI+55YIBBaGq
w+7ul/84zf2OmP/0xoTmaCnN5H7AlG2zjmFYytSzOscDVlzewp4aqiyLYLaihUFw4aq9Q2WTw1QK
YF6Sa9sRhbwf6HKBY8CDBJWgTy8M9NXoUi492dfM6p5l8d3raaEgDLDZ2DeFLCL+EdWknQvLb7Ex
OfZFE+W21DCmNb6gIdLr7gFQP5nUjCesFTu48aa8y4O2zOxff0zkBZ7PElqvTBWpb3ekzwVObmsx
DfGrhB4QWuq+JLllRhhC9OabssPeOBk4I2Ko8IVOKbebdxqr8yVPbdlA5rvjH7aP8Gd5aV+UB57O
c7yfCiiBDjzO8+jvAY3jJat39e7I5N5ti94EBC9hNp14oGn66wcLSOD0cO0PPQeph679b1LxGVU2
KQY4Gkcfc8yRqk4ngkDyjpqmN/Xd1UAKZe7Vw5SBtPk88kWtblSndk06vcVv8fs9U5pnLhpB9fGr
hTbwvW8cBSU/In2sNvneWEffKC1DZIhqJeFnw0TQKBJOCMdLNZOJLZ0Qh2PhANBbVWVvrJ6kpsbN
xxPyLouSiCgClvpthgSQtqhdx3F3sbW3weROp5Vy+on5OoWKMmyxYYhmofifDpoPRryiBvLi1Eba
AzCOT9g4SgDSOgdYEXEwsAMKgiMD4qvhkcsvQYof8PYvI94wXPCfyTto+OT2CKasK0aO337LPMXg
zS+MSBzNvFMcxRdAVPy071e7B4ydUxCjVCW0SLEnioXk9gC/8BpO8zslCJnL4GZ37+QKLZgFEIJT
23W5ElkkzQcMN+vFGGzl3wY/zJjBAJ/Aahb8zi1xcCACFbWhGLCu/TerbvHHPeyRt/wsHDW40RFy
Nj28KmiH61ual76Dubk3RsweNYIUDH4a34sYani4R5xfPXoqdWwORRCPWOna0NWaj5KaFepQEcEe
n1wP6n27XUaLTOqydaH1d4/JKBeTKJUj3Kl18E13vefP7i0P+55DBwJDkLxwqdS8dadCRi4p7QLN
by81Joe3uUGGegX2TH7sLQkJB0rOEnT49snVDzphzVNu0ghMDys9vNxnskCQ8eOVDChM19EKnaUz
ePl42O19Nt0nNh9mb5wHbBm161FCR28/I7RYcVu8hEYR603ZFTklIM+UgJMN16VThNf2SUvNarHp
ctxc9lZLTmUUQLdZ54btgRrtKue/kFVhqLcUtRCSP9vRM04Vx7+MHsxYlGDxlrWIFOyHekRnqyWh
RIhjg9MI7DoTzN7xQ2rNuWKwK3G7TKLUzrFa0Iub70xq87uCVC3QEAF4bs4GDJe2rAYRsxkn/CLT
VNyR0x0qbu4jjpb9RjudcPVOCT3O1ccb8GTnFMAaw9LHzluiDFiR0wUTrvSKfwjuvDnpdClROZtk
5V3FQpwlZuRLrGxpG/K+iUIY27wJyMdsQ0lsrX4VyXmM+bOV8Q7Jtq0VbaBszQ9sPFooh+yWHCJG
+6KkriXB4jvtH3dCQ/pfvBrUlGJlpNyiqpDbL2+4QYPIafgebBigckQtU79HOBJeli5umrIFelKU
xyzINftACpW/2yTZlx3cMv6peNo2NrLvscArQWoGRJcrb46QcOTROp66E0DxCm88rSIMAEo41M+L
HKuxM3zydCtHmognlmKxak+DkJQgIqw7JKpEdGRY2BT7VL9asbR3ghN3W0qM8fib8sbeKIFhNGmp
bzrPcMeyuTxzgXpjsfSCtsXIWP75IgcDIJNIBi5Qy32bBWIr3hS9NdiA2nkENVFvfRcpFME65+uZ
Qe80xTRtlO69VcCiFw+8YgNaysi9QhmRLAkj1W9PXTflDywiO78LnVP21whqwgyABIkhwrdlPmH5
/11nzvW8l8MpXAQrnht8QAu/XWSk45KRpWItIetQTCVDgD4ZqH1iAE7sq457R+11ru4gwyr1xmbp
RxFn0kmBAPwQNOm0micwyJzynLLThKjtNn9j2WrLZOO6br1+PCXZmFzxIEzt7iEx9EnGkxdWLmA1
b91uzKoDJWwOQe/JwNK0b7DwYEZxocCyCt7gqHEVYuN2UfNCxBtlzXYVKZjOnNwLQdf31LUv4qri
DMrdIlrUAjCXR/4UXt1QKR+p2i434bcnBlZncybglE7Q1wEcmE5Q9+UU47R8SfIvVUJJC7bsU4GR
ntgqlNZR2WUx33pUjZoVw39OclHlOuMGOnxwgqqhqhDrf1IJStuBKigte4lD1Yc4dih3r3FG0Lpi
QvPgp5yWk3LXM1nqiYrSvlO5TYLyFFMcoudbuh5IG2PvU/Cm2Dzs39O0Vz9WwBWa9bORCDyiAaKC
5RhxxuzWmgfQ9Vy7IqfUrZO5QvuImLxD/bICH+aW5HiAbjLkxGErlUIQ0cgX/6ZhZDaA5T9SaOfH
XhtDSrKzO83HYybLPflR4wFuUQBm5rYaVaGptDg9u4DKphPDuJwwN6ZlJSProxvd3UvaqPHY4MZT
1uYorsLgZjwquH1BKMrdx5WzIU6NbIphFIn//q1H65vS190cNmoeg33gDbo7WYgqatBsXW6ZPThT
JeNAQEAb31tpzCCXpYlGNocuo3122FKvGHPGLDonXLqXyqRiHJGYJ8moOHCHOGxveI0bXvTw3BQQ
UsdUMjiC2nEtT0tOgcgx3tYTlvzfXvw23ygfuYbYvaGligpeWfsKJxn3RT9tdGgVSI/F++9ZkU5X
uidS2WjVwW/S4mTH2ttpzDsx6XZBoAIT/0EuBGMOO9BVN76MKnQo0y14mPlpEq+jmkbNw5cyx6GZ
H7uKQa6/nnSy1xjZwi+8WJEN/rU7wLC4OxF4ENPOt1QVS3fjZHGggIRRGzamw/n01cICHlagjT2K
dAZHKhA/mfETC0zVVwMVNa6Az0l4b0TtwrdbKNyD99BSKGUvPKhdGAL2oF4b6AnJGOwO0LhHiWCF
wA9TDPjXRIC5IYJbMim04SSkob1pSq1cIhoGy22MH+drZSHp+2ffuf/AzxIikw/0tEvxzlXlJ7uV
3Z36Z8hlhCnqV0KTgvAo/x6Ar2EfZQ6yMBRHOPtWYKqAoWvRb/R7d3lHz86yiI9Qlouyjswoh9g9
DprUCXzRdncsOavKS2jxZDoEoVBwJC1hWUgIe4KkG8moR/EM8TqmeyhS1/m6cvDpWC+Sn0RDgVOm
55kULixcO+HM0NfesBRY7YnGdm5S/UA+pkbobAT55UoOVHWJkLSRy+fzTmZg1tcMaC5JOWajtGHc
+2gEkAMdhztgDs60RB76+LvHXQeWQf8L2YuQF2pvbHx30IyPSWLKQBBJnvDiddz4ZvPmzERb47+N
Zzu87YqRoGreTvMck0D3CEaoNIiUYRdXrGSojTnIP8Ob/jtxXvF5JbDwKQiVxnHQ7ni+JI6cfsu0
YNm3X30Irf8IjQQGrFrgh0R/0NOpY/zS5jnI9XBgI1ozYxeZFXnWsV3jHu184Nh23YwFDjlgs7+D
+XZJDt0DeA0Roi6oHIMzaMZOSvF5+4jhExqkMZ1FG1QlwtRA0dChscRszuAzTG2YjdNplYDJRWpx
8WijNYEZPJ6MhIUXaiEeY5HayIEGbx177m6e72fmj0aBdBVT1X4oXlhxzqsIU6jN01vuoAeU2tVl
LjXqQNJwhyExMjTGe5ZLvWnp1YW5SQguroWZlJnNPAbzCib8H7s4MKY6TmHxupTDS0TFUjrtURKq
h//F+626ZEpTjcm9bc3ZGvrcrSiDx6ognicjkWQVmd779Cr/dHLmwpFklggA2yv2I0qd4OMAsdx9
ftLnUCKNFhlxFsDb67FRTXEtnkM2V8/q3/yBBQEeEB5jFaE/z+0RP4UdfgKYgfiDRUSMiaq6Od3E
ECRBoWcoHGF1tuT9Z0Jiy8VQB+6KiTkvrsBHCDot5yVhzu9/sjGSkRlI0LpoQ6Sip3EeeqG6b6Ee
pYk9fc432/6uicdOx6uG2U5XSerT8Tuzx9sVsRJjdAcpqrYcMPupifIThGsfGfLBI1CMDWRLE/w+
GW9b7ckG70CfJPjOE5CQ7rNJnhnRzR+vEv4neHBsFifs6w/zR04J8JlDQvl5GC3jLEnoO1GZ/bo2
YBsG3WghDDIUzapdfFwO/GrdqyzuSrWBTnjYqf+44ALA/sgX53WX6E9af7gptWtnWXIS6J4o7ENb
B+9VSH11IatARQZxM85zVaJwVl+SvYHgOobY1UzqKvd/onVlKISrfq91LbOkSEZgiGb1Kjf0/5Dq
XgAlVWuhTuXXNcz6I3a5RVh+Z3IRN3n2Ho1bxFv69QE9CiRWjCXVtvKTCCmRwO8BCCVU7iC1zb/H
SSHCLwqVJ6itmAyWdRWuCR1GN678tn5Bbgi4jfmtTWfufbteHECTWUQEctqgCqKZLk5NnLXIfEBa
4WVC1anw/yg/lAto8VTn7TDNjxsZ5ziVB4Sg/GDeSrqc1ULjJOASe30WEEPP1ygfZ5mYUK3adBQu
3Ye2Grn9GDtxhkBYvQ75AkgqvWTeB3KzSHk+bLq8bSYqe0BqW22KVKvLSQozBzuHka+1xAMIZZP9
d2XY9MT19zWzxWzWMo7xFgfKozvZMDpxJiiZgpy/pfS8YkesLJMo9Beyh1M1S5N/0ZDnfgu/6Uge
GuldF+acT2N74xvD/z096kq+XEfr2dl4kRa+yrdEZf4tcnClQH2hFTWrEkPjVCmk5xRqQnZoRiXk
8sWg5tJTqTOPc/XvcJ8g1jeHZg2RnOsCpAbBZKfLltjqh9FMnDaqaRBC959uMsxSGi7FDvMi9G1u
CPO3aHGQenzmA24byBKj7HQWi4n1ddV7GJO6Rqj3sZFrrbiLZ23urg7zV4vNjAM+tWpRrdm04GbK
YdABhbG8R5TMcLvyqBXSAUz+v9FoBFJMBejUijR/GAsfzAZq61R2ITL01pf1AkRpb4oAePN/S56g
wAVMEYJz5MEPRj0m9F5sZxB7u7E3+NbvHAZ/sGtF/7VjfhVxKdckh57L8vJtrsICnfsiDX1XsxJL
2axUV/3R4HACrIrUZiOW+P+EgTbmEWNfsnN4ByHH9wmm2A4O0qpefdeGMQlco9LMTwsEOjITEpyQ
UwLiBqaWNgZe3luhgqAJjvS49X2NS08cKq0jrmWAs9DwMUZ8NiQJ+PRQ3TKguTqxY8gjry0zaKju
XmFtRSOrwa4C+qKhdow5zTh99Ug9CMqZ2Pz+4cH1l3Clxwf4/uWeUaUeq6czAdTdjzjAlPriWidC
1AdZZge5G4PhrKxnd3HWnHCKEiK/hJlv1c+7pw/5djbignBw//cyQzNVZqcLdjp9D9YyXAITiO1B
NQpDq7FVM1gHF8j8yTWCXhjyMrrZNO++k5CQ+uoRNxgslVzdxhC412HlIsfPF2MLEgk1kHeGlaXc
aerQKWEBSsKkTUQur9Ag/ECObr/nqOlj+oYr9lU9RlGEJZ93o9dD2CaZp2wGM9SjBugiprs68MxG
/RP5NWgGrdrVfOGthc/pQe5vvLqok7+UhpqW1X7caofu3I/a1QKfNJvexOrR2pxwBcMMEJFgj/BX
1KOHnapUW55GoeTEPxjEwrfvKYFMNKng8wDGhin1iunjjYX+v3ZZmkl59G5eukcmlxTzkkkCJ69P
My1LF6voVLYDj6khYw+jgBNI8d4DPBw/3eZ6BC6UPyE79EpJ2TdiQzvwhAHldEcvej/W0nypspx8
N04gL1C+vAslksfT9UgYehlVgFQP3qbySZgDz5MJNKgAMqzeGA0XcoY/s79DUDia5lZXA43hsrXt
RVKXpCm+lCVg4/7SZdlufkhDRkv7IbuGc7krka9J+O4nts3bimJvvfoXofd04+74fH0kSjK5rH1K
EdFsLV1sgKeImGLUeakNu5Xx1ysiC8RyRxdH5Fdbf2S8kvEL/0R87U6wZ/e16TqEbK8TVkYB1sb/
hztdO1SlxOd7Q1wR+m4RCgaonErZlWZtFFVi446TD0wnKTLmtHlPipGjl/wqLM5CgppSKW297jtA
HZliAuDdBXhzQ+8O5HyL/38NmQqRKKp1ESqfWHdAqQhwnDdwGZ42jasJcCww0e3Cj4ZhL7MYEA6u
Do/qHINxMuQVeKG/seqWzQYdBOWnSo+OB6hBLSPd47zGIWrsHR8HmJHMBI30N5Bcu50kO3aWPihN
t9ilQjPJzQoucKmlyr4Dquu3Oo4gzNcbek9viLxxjwB6oeAQEncOmorzZWX15TRZU/gM+7biM+G1
2MHI7KN2gb3gghSijZr/8bb4sNDSJN4f79uWK7czT4Z4/2vLiUQtlV4fzr8dL9Ke4hKZvK+5HR+Y
TsOykqvojahEu4dAeJChtKhAJtfOf1X0I098aDXHkW7huOKHDRZJkQnEqQEJpCiOLMdEuoxCZHx7
aTtzwk6dYY+km5v5m4P3DXCVHWqVuVoEdzIKh91MGNDcenwLHA/VAgMSsOCMwrOSEuudNiTay8yv
nnSjbYRSFGSnocOnShSW3tr14BNXNnOLKCvzEJdwMWC0yOaZgOfDbbKU+WiLqR1HGipDaUkgicAi
/UwrBam18cpWM0OD529aqUOf2Jp6rT4OXA7wgNzj6EBqCzyHJL/fELalnb/9XpCWrwc7dat4fTMl
9e9ZStcHA4GmgApnd7DYeq8+UH721E/mDkTXrNLktpiTV1x+rBFFcMwSFJst7ymzNstkKszqFKCn
anIKvy/Rw0WBXQox7vRkEuDBufprsyUwKNZDg/nI3pqxcm9Sml8L4C36oOkaNGoqrHnOahdtxxJL
HHBBlCAHEmCSV3OleqjSUvB3eEJHM4ZsFxTaSc1/zr+a8wYq9qmkxnb+noUsW9uJ6bVwMvDAB6QS
f5TceUE+4l+rYHVcZtvXKKGgZfcqsN5HTHeP/d9zeG+zkZ9zip+gGxCAAXwZejuOParP7qhSQsh8
klmHk6f6NLoKNRNPPO1S7tXooxDetqTPyGr08RZzDOK5YS+OzMj3o/fGFrqrV0hCl3x5jdJZAt4E
AufrTTNhhev4FA7lRqi9H7oEmC9g0sNRuYBNmvJJlVf+JLciENzJURlVpL+K0QQypsK1DwPLCJ2a
O07aBYZsJEEWPRvGZ0LM2aBskEjE31i2zoQuEgCMFW8Icb9j8eRe0opvgya3nCeMWTLTL+perqhf
ou4P4bhc6fRGkjZ71op1tcjoIKu6vUBAVNP3NhtTwt9/+Znv5f5VABN0sRD1QC4GySd8kTbBZZTN
ViKEwgOjHiH+pyiE56glh7aQO2XFyiUdPm0ARWI07nAzgg/N/s1zyaE0F6IVrvilsp7B4/oMWurA
UU5XppZsFXDxmmNGVzKEyZIlqv2OSPOUDyaOv73qbzxeUfd6VCGLfbcnnsSMFKT5DBdHOusYnK21
ByIotDVKmwVsHUvgg8zKAR2uQoZqpWaGjJso5HPUbWdRIjEsIiUTLTuF471tmdIesmsOnKg8blj0
IyVyUT5NN0QqlyLeDhQ7X5mMfun04dwTx2Cl7ax8QuvEEb56QrEG5lc9kkVaA62Cm6VaIPMk4tbD
z8NIDQwaBD2MRsayXfCmdWA9E55YFLrtl0E6v/jKV4qrl9LsW67cbXZixTp9SlRIBO0oB5ZtRYIN
G0FoH3/VQGsMcdpARg2Is20RYZv85rssBFhiLv6K+IkZdq6ml/EO8LKMMkZTw9B0LUFG426qc/jh
dwlGKWn1Ip8wOmRmxF5hTlwU3jULxDUl9jNZyTsgaBf1PiPxgbke8wsc5emml7Iw9AK6vl0/xWMa
glSbRlCQkP1ZOMeOiOUXIcLz0QF/1ipAeci0ilp3cAFOmGbcfz6UTZoFAb0idd6dpnupAdc7O8mn
yzonREv3M0e2X7cW/UOeMR2J8H3EELWZGry5WQpLKqJX52AqtFrYAudB7l6W8/uVLPg9bynVVFIL
T60vsKXpbyWy5CAaKhDS55ImMpMkzQYSYdHKovAL6sWg4I6l3gDu4EKqYOGFmjDK3c2ZEpT6/NNX
DIjeWxHjYcOMox8LPKoX8xVr9xL8uhB0Umr3o9kiq97tjftbvAavGDFwAkSpegUrnUEaHB8u9grk
M2JzmBK1pSztUHyGkfcJfmwFVDbPquc0IEci6J7vwwLYNENglpElV7AlteJjte5Euer/Y7UAcZzs
5wMiQR4uwzcWzkI6VzWIG/reJNzDh3gwf9jZU3PxEMK8S/tJBrLGjO/9RggYVs7dGc8h8VDdL4MC
x1UT1jySUbx7wpkTIW5wbkJ1VCERHI4hst61iXN8QmDVT9biwenVH9OoUsUSY8o6XNFq1lhJ6Vgz
JohD+HtDtttENXQuZoug4b8DvW60CcdBXNN8dKcoa2j9Ek/Hq86a4sxS97zVm1QCNiS4natjL9hv
602taPXqGbmRTRYeCncUED+P6dZ2xZL37/Sd5EOLa4QiVZ7zLePa1vgReWGTLR4d2Lal3zvLIdvX
uAMwHgLYGIwl4O9NAgQGtwXgL7Q4g3HF4/kzKc2fmvvtZL0F8gg2dwl3Qj6Qw5vfqA+Fm06T41jO
X86fH71KTultyje+S8ECu6c6oN9jpv8BkHG6ALFk1i83NbltR0dPSo4X1dWzBMayMrNGURKTI4n3
BBkvJ/X5nhQ1pgeyZUEBdI2f8SmQgxT/u9wtRoX43I1C00YL0tFYQNJj00Y5Xr/1Dkq5uJgPkTEZ
yIJuEtx0O8Ui3+0DQXAQ0a9vUSAbzRdkClABNrgZiiwS3agwn+ocqSUf4v8pRbOzNJNooYdXxPkZ
NIqM3LCXKTpRvCvGnuDOQYxpR7roP7oh/tvBBzacQ5n5vvTwlZDyBZZehR8Ussq00XzjyG1JXkqM
0xppHbi6RSjQdJ/3gF9OlK9a0nYlPbqWOZDLmThsiAJgIZsDQj1WXCD0YQwy6SChgjjtn1g7mKgA
5zyv+brcbW548d4T4rUnE6a5hT3P/XnnXFyXjfOY0LAiTdqfuMy/B4NEIy/hZUUr4izWemKlsNUR
4W3aKwYp3rsQK9TV4QM8Wa/zE2MGBv/OzRmq44F88JUw6ywb7r8g9BGqPyTISWtDjY6QcMjDWvmI
6FYKD2plvJYaRqjvq+I9ruVIKCa2HHNZkMCwRwh9LJJOvYwAjI42cuAxHqsgILISQvn672W1EQYM
AtCpC0Syi2G5M6A3F8LiCygYA8OkSr4Y50YEkCTccve8S94jQwQC8HnfxLs3Q9vUSKciXbevmXDm
+yZWtFjL7drViytkHdFVqgYYFOPaQV1y9p+XKZk3JZSk/nPDC2alV7sUs2QkTw9hFkWblVSBBKHd
6+FVTy5SVPGiVHI7x7FndM/MPK4iYHMKZEQ9SUruxgt0P96xM0Vxp0Bxp694aVALPtMbpbqVcwMa
Pn6ClZ3JOJcqBNZrmn/zaUmRa3nYzHfaACw4zGuXVoy+NF+cxVQazJU0XO5k3dswUrrocknfVaDJ
MlybmVeYxQ7ReAZzP72lD6DFIdwRIGNCUI+CtxjoevGZDBEst4O01d/qeRiQpvJQnc9uUo+Lz8lS
6gUL0ARMCmmETS2ZTq54vwj01tsVTeklQ7UIY3ENC59ZA8LM95Dk59lNff5fpRmR/aoZAIEr14FL
xwwfG2Jr+6zj7ZoEPdpnMR+bZZ3Ddxf8t+sm5Zjg6HJC/PsChLJ6iTOgN7KJdkNnF8lC60aRPuQL
OgcIx4S/ARqc03oETGYtG7keIgiPsmPRRA0t22CAc4tEebKiImbEyqJOtZaIYjURERu5Ws/Ej46M
jv+RSn4gAZdakAE1gMW1/iLE+GqC4VMfJfODZDezzQuQNNVp4Vwd0HlNIzk2rrdQVu1hkpTI5+jP
R+YbEaXykk1lRhKDpRHs3jhLf8e23B1N6W6x8Rqu63YsrhkY3IyoXhv0nkfh67IeBDHiGUs/Rr2W
f/uzTrXpOHmum59MoUf6ThYBSIQnw1i6HBmUWVvsOQc3anNdD9XC31F12wOWwkoKZTmBQERQec2o
R1HYoOgYrYTJJP0stODZjMjtRA/kmYFXlw6+sa+ounOUUzdpiEdSSYVqO9+6fhXpjX9VA9LEido9
zy+HtZNkOzhSVe1pA+eJwZviqLIugfFRNJeGv7HbgYY47MNQltPgpJEJdbdhoCLFWhi51uHWugkY
ffV9rRBYeZ/jXoszyF0Cp0AR4H+cO+EgtE7aJFvYgTxqIrTq15GtqCcX7W/SdmCGXXt2D4N72rrt
YmDeeLRsVaSlSioIKQcZxJx5AtfgqqnN5UTrl8cgTRHjW4Xd376MSzmbmS4NVvdzOHw7ijAx3o5r
JDklqIkNjX5pRJbUirJG1BJSALFARau+8sB91g8NTukYlvrj1Y1gtSI2SFMhB4tJJ9Ig2gDB1K/H
tx7kKbGb0jSBIpwSZWdvftwxSsluTQclc1lp89QeIbHqg+5ceR6Vrv3QnAGs792g3nUK8zse7dMl
bXIaEVP+o3wd89qTbecYNUmoavKoafEhjvW3meVLJubquPpF3h9Yn+pp+iUkJQPwWmWplyRzZsyx
0Z5v7VyFRWUmUXl40j3oXEfxLp58m03hnbtGLgIk/sKWM0yncl1H+6HL2Bm8Qj5VcPE4AMcxHne6
xBDbWgaQXUAYsVoL0+KjFWcZNhkdEXkb+GWlRE+erD1/kTyDXNZQSbIWZDs+N6c0kvx+95pRohN3
yMplhs8rX4F8k+Be+mjWxBcHpB6unZzEuB0HVCPs1t7Y2pbqQQRCR9nEuZAA4kmR4rmXTTGCnWFe
k+DtTCNzdAiDZR5ZFtKqzQlJPTQLOJqYDd82IiF6ga1mvVKJe4dktzh54Xm2K9+pAIN5yW5iipml
wbY/8i81m0EQ4fn3WfckMan4EJTkd0nkkvvWphNn8l7wGB2fwn2IBmEm4a6T3TQRIdSptU52dEYP
neKAEaCAfEaJrGCmzLdXnMMR6PU+Zl1zj96CugXYRwoDaTxY9pE54htSgMxyBnxAhJQNP9dDVQgm
9YKVDh0BIB9QHc12Q+bscSW/6vWUQ7kvQWRt9PLaMMTSfWR/6/jrL856WKeWvqtQF0RuuMqQpaSa
WFDRRSeBjLKsrxxFQgTvHubhPk4YmnAWT1DLGknXM0PJcMvBqTDWo/kKgI7WC6ACRXzOggwHzkEb
Td+Ch3DHvzB8T+gVzM6AJ3XtWUAdnlbXBOVeXV0e1ehTEf/OT9jvQB7iJs2l9HNU1nNHoYhX8Sod
8k1mBhhqdrGl0405eBxAUcsLj79x6hNIGmERnN1Thcjn1vTLh/Pd4ij7tA1ewwzslauiHzQ6Aumm
37UU2Wmen7ad/ShgOgBSO4xiNohkedQUlil5SF3aSj6Dzt9NkmwWgMBUCv8deu49SiwuGPmhv2go
eP80slLos9hGHIiY+xLbQ1xVIN3MbNkUvymJTTcI5+TIA8bPyFCotJfrZl8FkyGt1kCW4Pi56G8g
Oyu0LpnTrl7v5bvs0gvlxHxN+EtTFVmfzQZTnCvvi3d5eJRN9ByEWn9tX8NnS8HdkeMU4TdO/3JP
/PeC+TqOfD6pBKjfubWOSqlSHMesaIK/lSikQP8XxUbN8og7hYiR4XaRIYEuEYLX4hcBuJW9S3EK
kKAaCxFRKPN299T2XXN+JnJB5JGLSm0FjL9oVJdRA4Jw3jNhuHid43ay8ylhEO9FsKhqNOvQLUHK
iCNRkwUyrcmuoNdwr/ossHjb7Cv85SDb0nktWsAY9WplPdBBIZrXxjRQmt/J0iTnsbJ9PZ+26Fy2
YZlIUBJNCSKUcm//UVBCG8DiSyF7O4aitNDv6Ho8zfqObVA6PgXm5svif7r7fwA4o7H7PYwN2jnh
Hjx3/Gz9C4KV8VbS7kGhxr9svwWHU1Rv09OghjBHLgMSJeS/a1MldFHoIhopwk/I8cY8isazUSwy
AWUrsA3iu0fUcU8fahLzYimP1L5O6qtx6tQW6pYz/PZTnr+riLqZJI/lnnw2sFpoj6yECv7aTZpG
Tehx1/g5E3bispoGy00VntninXPcRMeie3LKVyFiqW49337CYxc7UQYjj8BILAJBmoajRP6mvrpJ
pNFM/8Qg36kiYRrtNGa4nVVBLqguQ2fX09FKUxwaiGu49zNhZFpPuYYV/FIBtEh1MhUdyBqd0XCh
TSBcRbCIzQE25/5T6aMHcuesO9hWCyoVCFUGVd9OSPBfLykENH2HsqHyA3ftHJwEpL2hihoHKNLA
6iHMgdB2XtHrMkik/kpNiZMi+i8SjWZFmt++ZFxHLTA/9ANLggqFLLcjkPkcS2u3x+DWFjlCBJB7
kNcmxxMLYLFjTaaAhe13tqhL3GMpuxbb8poW8y6+2HWge3Ug8GJR4tbDYKsu1ajDZ/akqIjzJ9kH
TIWU9R2aLuETwZ8u5nk8MUoMjfsH3YLkQyoRzxu1iFrPX95y9Hb6GVGeQHLOvdmo1aENI38tahho
rmDk+kCM5oyLcQUs0ePG0XE4xqjlRvJbI1jJM5sAx/GOikHwqZ7D2TzZKT5QBjLI9N8tyca0glv0
3BSikQDcRPH6073luXak71Rh3qQ4pJU7krqI1XS/kK3XfltASJQkMUK7u0vw2uTERBrv12cQjIxF
ttggdn2HJrHbgljB5cE9cfNwvHI+SsnMEszBCgIsJa94QA5YnNd5yvl45Xf0sfoq1orWEMgRW0Mg
afRonzTH69uFsHhZc9PTSKWqwJ8uEoRlRoFECaeSOhFO5USen2Py+wqsexPJoxHwSShIL0o79vXL
BaJrTtOlX0lwZv2PLwSle/Ikz12bs9KOY/D/YKJ/7JmXhOizdBcgI5P2x9cPMJZKVxcfLOrhoZMx
644KzS3cuaC4vZSCX6a7tGpjhPFn5jXJLZG52+toU37/5P7m+LsQZcjVbBNkQRl9sMq8L26r8fTe
ZEleIqFF6CmdHiP/b+pBfX2nGbTXFyifY5G5YcxMSu2Ms4Dp4vlYLHhtDJDeyNKFtOUvjEMEWBfg
k7N5N/Xf3ypBXjTilzuCAmN4DeBz5E466jUzsObWAzkAEKWvHbrnBw6g0/BK0a1vX/T0bDDmkNaF
mrjvHTJ5zJWeUAoz3uifwHb8qEZjp7PsrZlGomwL6WoLxaW9MUwAXBa1Q0FtioLD5fO9rR57CllH
K2MLs7UANSkBj+mGNL5R/sooV1dzDCPrVmw4rGZx9dm3m23FSMHe+1gDnnMs42RiMrwvTpjfeuqH
k/vRVb2VHBFh5kBo0zq1k0v6+ZJNTXuV0K1b9EOoZiioetZR65foKjEk117i5vHlNAXbolhQoLU9
rda4S93qTMrK0nyxT93Prh9VJU/2mz6MiCtl+jfOwoakDmPKY5srzaOUIiF9XszieUfE4xhGRQGo
kt2CChXwDcpFy1I3EdQ1s2G9+MDj5nSDqwo/mYYImMudAoqM6qrAKb1SpVgLsmANcfnWjznUvxaJ
hgIpWf8hC4ZT3TV9hgGQuSHsFDHOLJ8nb8k8stfB1oiJmAm4C8TGAmvA8S6v0Wz6Gkpp9zwv0Ekc
685K53MwqC/kRH28X8TQ6Lv4aHPE7F3R0wCh8gX/wkPXD6Rta4x+rQD1TxkwSf6vyTggQb7pP6Ha
KJCG62zsbDMAwEgI1jz0hFFNtWV7uhZXaj+PP0r+bHS6ePFAtAlVQy9iOqZBNdsdfH81YSeN4W1X
sos1zF1FL69C1S9ahrl57+j28PsijJUng3HFEHjAariIKxY3rpAfF2tb6KiNdqnNmqOcuqK+bkzF
xWXFcbxTxd05SqQYuRFtdRPJ2BM1IlZWpqpu47nPrPAlpPv5Ar746LpKw6jEBZp9AHyfiW9iTebA
grYF+WJLK6SKzFwZ1Qo8JBnsBKoNixEny/SurUom7N6esAIeyEX5ubKfaeDEhVmfgaPV4pblmRtj
rP4UPGrqwaDbNt+lskkDwS2mcs9r1FE6S5PRlmqk5btRWDWqAhWic1GGyZdf7FqNjGcVFQgvyQNw
ABcaTKVfsI+QEIEPb//9qi2wuvwsvIBVmU89MuRv4o/jWiQtYWfSf+gtvUu1oaR6CzkeC1tGncku
6iKXzn0Q44sReO6fhlvKc5MmAS9po5MhtB7w4C9dCtQIzP3CAEiMJdzBkc0ePmJgvV0AoL1rKB7U
rPikVW/Pr8czpvbHHXkqYVXhqwA1ArZ72i03SM2idlyCMvV0OkvdWMVIP97AUhnsSaIiCsRSUzKX
ij1+LbGenw3LVA4BVuvXOEMGewplWZSrTW49nmm1DOgz03hUGG+BOYj/AC3kCZ1TLUh1pV1PebJN
esstdfkQLGNLxQ2In24aY8fr0p87z0J0Y6sxIjNhQKgH9tXt/oa3o3lVOc7A4j0gFM8Lg4OHxI6w
7g6YszF5kCtatyxadorPa0trArFQDN1SpW+PMs6LTlmk0yXAcEqnTQo3OKLMg21PSC0qXRqr93VB
5xKYyFc8HPGbfCNyNAWaGU4H5AdTrKasIVeTsdagzWHNAHKnnFJ632H7Ch1uhG/QFXwf8LcU8eL5
0IO6nYgngw/K/ajnn93cCdD37xtmI41A9zlToPivOPVNCxC0fMtrN4a3/S3g+eAfaEgKQ37lIdfD
NlGhVPegGbMcA2xGSD9Wu+blXu5w4Cnul/IG5CwH6ZAGjE72N5U/4nFAh8OF1D3UI4rk30jrrQZM
P8tlwIzQKISER1jp4mV3TSFp6SOqtIFZ8X0QnjOGcBxZQFF88yRFwASibGuNPUz4ehumMub126SM
nGFZ15qApitjqcDd6f3F4HNfXr6FtggPq+RZ4j8H0doXdnploiDoHzgMYTCpEJdf7yKWNjxHTdpE
OP/xgS61YFy/M6rb5irTALj0G3FBmeoV38oqiVCoEu6nj5GDuEkN7IVuIbLYYkFisQYZbKew+tBh
Gc/HNiGAURkcjcx7mhnusK6CL4g36BBaRB8eUihnwuJ/tJBQqHCnvLawbCiB2TNEhQuZjCY14dbj
3CK91Avc9YWyt7XnIm6RI/5qRD6yJQwrgrJgi2qG9u3i0FRolox7/3CWpl0Ue3hCSd3UnhabmEDt
GDfmZYgjpmyFQO3/Zum44UCXoumj4GkMxx19vnzkGM+zgLg95ZeJ1CQPipLd9CSqi7EGYJS/hqWY
S0Xb2PdkwIvG+3UyoMSVPCojV8BeFP6bggJvZDkmvCmd1iNJpfOGJC152hP5W1vlgkP//didXEsS
C4uwN8oWov1a4MPk3buuLlbCHaSi4TqgEYdPJa9yBp65Wz2frT/OfLdoJ3yN21FGNqIf3AD9E7c6
HjVr3wyPK7wU3HGmgJSL609juCXuejHILEKRKxlVn5jJk7SksPhNm6mIXFCD1cOf33X3jNYSGwO/
RqxTxzQFR7HQWQrGNmi26vl4robsnv8qphLONha5R+P4rQmx7x1VIm+MKJMLdppkCzfhqGaAsiUM
dIIAHVo/JrlkdR7AKv07TxjcpKulvVl3GpWnaA7S4N006iEfouVB/5tG9c1yZmO0GUeaFRB8FOHk
HWREASS7lpaT39iAVYNXnVoDMaXb9BO5kTriGztY2wey3/waHLxnMtk649JC7iArnJ0gppGYGVQg
IuQ7ohU3GNt6guMAF8viRbitoJNH9l4oLALy6sL9Xb7Ksg/MPi9DBbVo0Nszg9bOEbhCoUsm0t9/
2xQUzaUao+E+9JKiDYS0ip6hP8mKm78PplqFyoYq+RixBMTfdJX1My6ss6aZVMuyIbKEhwEoFLQ/
aqx+brXaMvzXL307LgbYfNxK57vGeNa8x9faSW5mtmnne+AFcdL4nbsX5VlS9p03rQC+zqz67KKT
gIyCquXwqsbpFeKccUmwrQzuxwXuQZIfGmz9O0Tn/YpO+LHjbEQi2AlJ+0c3j5YTrKPYax8ntk0x
j4Jk1mpGIdAq4T2peAw7H76L/FbsTaxMdkooHjMWT6j+y8PWUo/mp4NQoKemDXg5VOs6gqvb8Uek
zIXI7sSQvOdITuYUYrVZz0q3zuS4QpdmAylB7sbJUSW0210T0XALcig5lbydacJiB/GTzxOcJw4z
tvVYQfw2tGrzeZwt5B/dIxbNxZK46qggPERO1+JjCEgEi5kAKJev7LBkkeuYEoLVLaemgoO2X7v+
PvrQF8Qa5egYNm8YHOVUGyVIS21Ujq5smIIMs/0GWYf9sSQAHo6Yy+Ku3y2U4m3b9zvt7sYyWXBp
1LD+w/wJE4Id8kubzYK2+TKOArgCDRB1gWEn1ZT2l0AKS63ACOaDI4odCywubAHx7QI77CXm2k2/
cezDTwACAXkrKYWDZLUbZ5ddIn13BToUwXu5ZJjtTi6+VYG72Y3fOKNKSbGl57t5pfEzlJHdQQFr
L5pCX2wkRNgCGxKl8O97lw66hxZQFM6apVfeOJM8nxP0J2HrAwP6kEQqbufubedckAdiS+LtH/hr
5FGT4X89R87GKzRpwvjN9QyzegK34LjussA+bvR76kavj25+GixPqFIgwbwr9RGZx3/UhJz1kxLB
PJ0vKwszERThpwbaCZvNU9YVHphfuU/X39zFZg8z7db/Y4ffuHsMUogdTCJ7Zl6djvvTnw8YuE8Y
rZ2njTPBrnOrC9h+SEYQ0FeB3XCTclFE00Vy9tUtMZnQ7ZRBRm7IrvxZOaiidar9qlDxUj1K7p5q
UepbsVSbmQyK18iOFM3qzY4MutCfiTnhOp6c1YkiqKx85y4nJqqhdl+Ueyv5jXVBifXQExDfYOX/
3EAPkcJC01c2OtnB/ZzQbNAr/cxE/09GvQkMQcHLeGoC57uxo4x2FHrGUHPvYS9KixHAsLNEfHkC
NglIruQySKOfB5IYXRLMFEP4py0RkRBFzk09xZDrVyPrx+mIC9LCIvlo+AtE5WSXPJxspvVpR31y
++UaQsn1YKkc7TKxofoD62DPbj9ckgL/zVBLg61QzmwmW9FirtRipqyt+MYidQHb6T1AW8R/Bh6P
NQ8fy93MdAc8HwTtdJL5d/2ZVdBtm7ry/nKxv2nMb+TAtK0fLdPs/EsUpXFUy1A9TdTwFMUMQZdO
A4JPtjmzWvwxHeh6XgN9lhoRKFtdRATDN9PSwoXW+4ytJqxmBvVDIuxK+YEYb4GK0qYCs1CFAMvs
Gxp5a7OUZkO/hXpcbtscovcryDiZkHa7nWIImmJnbEzd7/WcKxgfGbUaYjunmGQ3Iq9PsJyzFAxC
MIsHDGQ6O2VxIE9udCWyj0iEcdwunAKVkXLTHGKZtB98uHg5CyI6dGJfGRBNQMUdad9AW+/TWrhu
BK3ugiWH38SAOHETL49GbKjAPnsYkADx9pN/tTvBGHuoGjG3usfG4OLEeWWE0Yew55yNDjUrrLbC
PBibJtzXbp4GoW5IuWjgYjkuFZVYxxfP6C35l4/nnfjRC81cA1gW0MNIWdiIHjsFETkFqIe4BNeP
98oycDrg2hOjrROZjaZDlYuNeJPBseZ4sabQaUZQZiOMY2GOhSkmmGlLa6QY4aUl/8YocK1uor/t
iyuJNE30Ng4QxryUCR/ya2hRxg+51bhKXwzbKBMAUzdSOmdmZBMao0m6XRsZyXR/kvDzXKsTxH46
cr0ZhE0NnOlvopI8Ene7TOOGKWhWVzWTelOOHPvQP2nJUJCfViThPo4fnxUkFYGxu46vlnuRgVEp
URVLIwx5Gi5l3mVd0zbL20ExGD9CrnaVV3tEYO9C4j+kpuwUIE9ZHCxKrVCLVLNUvxZ1YXz+2zrk
SJG0DB/twBggdgxps4rS9VdeqVn4KcdR+hXLAxnbGAmyC/ZgapGPrwvP1nw7tzQNgQW2RVHQlvOH
MmoIzW3th/K0UTDhnlx0DqYp/wfxVSmNZQafozNpMhJt09EHRClEMZEZVKaqSMQDYrp8Zd7QlfJ5
1Odqc9pvIU9o4tae5pYmzDyfety8VkwnyXxrZ0Ikur2G2R3mULOtb9IZ9pNgeQBNkuG2kE7LuF73
B0sfR7eWpgSuE42fd6fnPMy4sFvlscPiU90wVcYoJkh9xt7PGOWaDCp3R1wLZSe9ba0WNiphnf1B
sRDGeRS5T87wK1ZUnD8KmmYII0gePAqgllkYPNkNyP1Jmd6Ym1ySc1NDZNPAEIDUcGHEBrHnt/H4
0dqigo7gZPIC2iE6ofnmRFzmqTO4dAqxPsP8mIqTnwbJ4phPDN32KZt4kfSVKfZyAhqLX8bw/mMN
udMgXNxsOMV49/hXIwI/b4ypMKfmSlMqH0O1U/UJA52/VIECqRs+Gkzh8ofYmbPjAyvXlw5CpzfP
5N1+oKB6kkwqTG0hjLWrmpgQN0pzdlXUDZ5TLknw8sjVnk/JcJ639+nbyAn1zgeXMJH3v/t2DDtJ
JeUvcC4WNrvHq+0fUz9ULMRXgOi+2imDxDte8trMAbsAqXsNN6K8KyG7nYJG9moAcLqMUO0Bi6mF
Q72W694+3FQd0KWes2d4UysWK4qOmMjcGA2j1xA46PzkQjPRrZi6tjZVz5ZhOa4ZONglk00du3xD
FRVDs9f241Gp3F5mIAhQZhJtJMbWfWVgh0xv1dCoOR53jCnQhU9eZD3TKOfmBUPISq99rkgjNOy0
ZthdoDb8dpaazYG8sSnsP8tX53VJ8bVKOYTqPkNmy7F9/GX2SOpKr1X8XPBZfsVioYzfVwc00/lW
10zHo4kNtpS0CrggCFf7Km/z1mo4/QYT0kAIHjOMRAqyzZCZkG+ZutxBtLzKFZYaHZKahWXlddKM
y0pKmB24npEk6UBNjS4FU2LPVrhIaSKZlsNbjcIuJ8eHmmKemPT8kMxj4/IxCvMk8HSNG+SAHlbr
D/BHeUOmRFH4usZ/dkpIoDG33/CdFRdzuk7xQfjYyRDZ43PBvqeI+7vC5GYHw09u3FXi5S6/vcze
MdCsDiPZYIrgQsUk7VHy+J46SldvOP81zgiUk6+FB+oDLJeyUybm78PUuq4DTYiK+J3j2IA9ldUF
PPe2cu787SwVQIFJ4RekafO567wvN4KoyBv/eqT5V0BKZ7j5xci5T/wxHz1pP86/753Haamj4/Ku
RYNq4AAdXaSDdBHhUQrEw9RT84FjLkZx2ClDhexkfPDz6Wq5KyNJ6NxntdzibVHuLZIDYrJsLAXS
tGUWEHCCfckPiXincFx2KC1ezLthQJ1+IUGb9GHAfyv8uI9tFwBK0RXthNjgYR8Gsp7zmjfTD1JW
iCaWpJJXNB3h6470G2wyqyVwYcLkYLpNR9dNZbQLYqsusA9oHnmCve4Oj6d8NGEr21VRJ6NJnyPU
55euMLX1/vklGklCsxGJfUoEIIlGBw4/Uwc2GyT2dOI6UAoDY17hsKMuLUQ2WRGB/MBdXB41DkiX
8YXCuo2NxRaEmWbU4+ICeqjM3mPRsRRSzHtnLtKq/bl/vYKB8gbThzIsKJFvDP48fVutKQh31bmn
Rde2ToLxhTXl5VUBTOGggN2F+yOKZqNl3+xS4NRrwOMqeqdAPqJQHg8X+qtzM3hoi5qY/V1uVl1Q
dcV7PAMt1IjEBVDTOZyJwbFHJhqOXQ8GvwJv690/l3FiskyzdyHgsMx7fV9rHCap1p7eVXEgi3+g
PwDguHPw8ewY5qVpJVBqT7y4kh6gVWXN10rkIhCpQoVrw23XA94icYQna8bfP/1FS2plpre/3uCz
k2QrSyE/G9wDhhQ77V+aUpMk96O9OIMzk/ehUKTpbvf7501boXc9W2yrAjAEzvaQB6pOYrg5nL4O
4Qitv9aSQhPapemf4PeqPPcBDPeZHbGp9d6rupQJ8nPeb6ZXTEASbq1l+qnqgxDGWQRKhwz2WvlW
XBAXwJ48VPFtcpx9sy9kMsS3l6VFflAOaRj2r4K7/MjeAVO1ApfeZPTicmNekutAfQXD6UEDeG5p
bNs8WnPXWFrwmm6DSIdKoA1KRThyPAiWcPSgsI5OyrxoJCF5tiLM6z/ha7jGSjMnLjK0n4VIggKO
vv8GX1joPPQRNVJCZ4hFsf2mmAv+/3xh1WjYNNRnLLvEDhD61UZWieheH1vgzwStNU8CPRp0pOth
In9RUuazHQrLCIKDX5O/nw5djAAw3+USIvKKrmt4mj7fj9lthS+9bz54endwScGk11g+UIaDLuyi
cK2vUK4crgHJXua8W2GDE1JAbI0lk8yA8k69zkTHv4aypfh5VurhnLZgv4mNGiW172v/KSpjCj7G
VE9UMqIqUWc0YstZrjBLFNK60ZcGLqhgDl5rwGVqDEn4v0Hyzn4LaMmqyYNEqT1ykh+E0glsLvNM
V9zUc83m1bkqDkjZ33/Boh+YxaeeDC3kRGhWmZFG5CPqCK7jnJiu2FpV33OscdYFtVhOp0DV6A5Y
WKmgcT6fzREIiC42TCBtuRwaP+HTXVyXNo2gvG20nLAtsijabPd8EWAkBYZagkwBn05gYGF3NutZ
PmoIOyRkaQGIYBsX7mHaErGswyBte/I33JjB+ATxjputJ1QRic73enLFs0kyU5Taq6z841eONyQT
7JkXejUpqLZ0EXIuM8A2f12PVlxyYHNB/hilTThoj8a2wyDtjWg3I1aDayQO4k3sDmOoZFDgVpGT
8YiuCs+ap53/TJCSBZZ8caMENXBy+gPNqersG2zDmWYtHQTiqz2BPPRpbjlb2ufprq/8P2zSlxBl
oiN2oiHVemaizLyQ5FtmpxK8TWx1HY/vg08T+Q1b+V+3NPuZl+FhoDxlGuNm8wgfAEHsqsWU+yeY
qYJGBOsLq0NM0K3hSkZNzjmB9GzvT16E82lVpj2oSTEKJbQGuy42VHte/XTWMnCaes89Yz44s3xt
MEZqtbZfSFxvx+K4YqZ35cSxtYfaEY8xeT9uiYNiN5iMrDnDwAyeoraR94aC/CG4S8q81jk5AVFg
TnshsPiRT1GdeiBJbwPV/jO08VFy8aPCjsT2euMqbKTYHyY+obOy2Yyk3GvrDpJI2bDpAdaXCgI4
XckP89a8RinUoZQkavqDcsElY/iEQr5UWLav+UHDuGu3NfSgix5aWnOtNvxiTPNpBEYCsEoIc+gZ
zF67UE21iwtgLcZrkJxKCKD5mqGNHzyNSxVC+45kd7CPTR5TGHKlsv4/b5vO8ZnCSO+WukLdhiUN
GjHC/j422D0Ejo8NnOWmoOWyC5kpHNMB5GjZRHzWBfb6+N1ueaTVcId4fsYVMsATv8nhNmeIX5Dn
vhNDt2jKy5RE+BrBg65lvkG/N+7WSANZ5+Xqrkyivn/BvLKT6FTaM/UAbjlaaf0d1dOhYd/nmNtV
FpEyLuj/+xnWsH+xG1wUkZ8LK6KRvlrIT26jnCo8gu5j99SpBGanu0jB5R9cESjaOqA76SHhDAro
TaV5nQLY5M5ctF6l/WrTjCDvR7fOuwpW4TFnHrpM4vM6GRH3eSGoslcLLn+IzMUpRoiYgLFgoU9P
Xat5EcaUQ2V/iUE0jwh+71unUfqnWo83nPET7Xn7eOd8sG21kLfgpFl2h1D/Y+4TJgT1Z4Kt2E61
OSX4LN/w/x4RIsfoUuwHQdayP1jstNgP34ezmckMVqyvnaKQlCkSkglI38xVt5YglyeC9qYAJ/Yd
AiRZXQnMCgYe5NexY/epENe6dFZG1LpiPhx0RqBF9O+85DgTVFJttF6SdqpQQnVPx+rQRrhXeGCm
cWamavkDUraGLxLQ5R68cYnwio3ys8TLSQs4WbbRkP6h6saybVBf7taTSye8JDHTtoO7eSFP/DLW
/S58WhLQ8ynI/TwXD679JpifXh/l5LKeSi5Lrm+K0DtLiibD6PeoH3ZtzYtuelKjG3QNGNV4kVox
AvzvbGBjx+M8frMY5Aeec0DRh4Uldl2wc3ZCNNDjyvP4cRB6sr8yU0HQzRUTUf6bgGH8a73ptxm7
hlwJFwGtg8tsZF+GAAPUDmdIScfNy9Y4KRJfzYEKHl9G4ua13NsWmSiYh91Tt0CH62omP86RU98W
bfwLEdEOjYyLEdiPeT590phaxMKTFP9mZxPkcyIHLRKqpHC23p7SL43r+ykdWEg+WdziAndJSNuM
bZtlNbcbB9jwdG5f76DyGuVYzK+V0NuDqN/C3kXMX40VXN/rZcDy872LN+I6Mxy7RznsMzticGQb
RCj3cgUfKK5YTR9HcJ6qxXzP8Rlr7JMnJnHT5hnqq1ymR6GBSwrmgPyqGGu4TFyaM/Y/kfDqU/Rp
VNnAFLAYwNn79SmErk4viblCgoakLV+o17am8NcFb3s2+kyvlJ6OQIoJb1/KZFFAzzukh2Jd/q9v
28glGPYhHKm7ur/DKn26Qd5COgQ4VARJqzH2qDy8Ag5zzprKz89vQd2LIc5SpH86Q40hRj2MfDt4
Bu8GZ5OniWXew5tjGeKCYo+bCCiIigVmb/MZsgewrAr6TP79Ty5dupKkLJNR3rAncJhtozLqX4nY
4mnqLrcvGMlxy9nWzVo/pgDy8wexQHJ//WDT7zuqb8qlWlW1J+GOyAZi+DsexNSqE4mUJCYlUdbI
PB3RgJKTWXrwjcC/i4F01+Y67ax6ghIiEo9RqbjoTxDWRc1ScvqVKz4xfQwVKSsOTbwKIya4GD0w
+klUkViBA+3hx5tAo9EtHUarcEyk8uj1QEJMZ7II3HkF0d/skaQTsZA3q3hhNXqN7zvnkFG5snAW
03RBjZ8sbScApnKQrmjciG406/hfcHctlL0MD4fTfNB41pSxJG7sqYLl0C+LkqczNgHjsHciH3Gz
Xn7m/TDljMg2y50vowutYDB7sEqY7blsISAyVwKjISQbY7MVJxZyJTr8FIXeocEyBvoWdWMsuTLw
Sf/ZoHn/PUTJIND7qRkQNedEWcHqTtel6Fpe0lWpwhKZd0pFKwLLEg7MWfsCIAi9mTtQMUiQ2YFP
skzLIFL927Roc0xor0Tx0ZU4Z0m9nnxS/vfTNz8frEMMH8zaxc2v4BE1R9rYmAOquyiIp2PaI9xR
6/m9L3Q0X3zaWwoRUxJMNcBek6WanPYzk2v40RcydZkEQamoKOi8A+y0o8c3sO1qCoSVZ0+f7gL4
wSKBweJZhSGw+wnrsNO2BtWCB/XjXYKCl/CpgZ1289tv0ZYspohPjRfvhO0BEdJaG/7U4RTCvBky
fxkglq7ZeNJ2O/CYQoA+30xGfVsaQqtm+QKQhS5HvOcr9XcN1UZ5gQTfZr2/Mp20SkJWe5y8uYl3
2d7C2gtmyQ7joLVOD2h87mN4q2w1EYIO04nFXVBRsFFp3u29sAnqLAFk7EdMRrzXOo9PbWls6Qea
A+MGLv1Fshyss7AfLqCRp+3qXnIvT7IjsOJ7dJ5iqPeZFj/RUisXyY2JkRaryDyc4FNrf4ixCajO
hgoD/3tGz/7b5lh3cC6arT2qaczwuCfyNo6fexODyn4seoc77RNVVh45K/nIDFRh53RoMjwHQNMe
9E8abBSmt4X2hp8d0OOc7rAzJLLQZzB+wyzihQ3d/CnC1n+zeVdvHsVKpEnKPXEf/Qsk/rl5qvuK
YcOs9wklTwfiR8mAy+vuV6JNGWDogph7lomM4iC1TD+tiENv5V8gJucb6L7GavNIZo5pBkunwNRo
ZyqScUIVXJ6Zw3MhVTs/ZjXfyOn09XbKpfH2oXqSU7LyLLEfjBZhotElVZ3XLwjme7X548pXl+8p
6Xf9BaPuVbXfXOUE1PDyiNGDIXVXPvuv/vhWqbLrfsrYA8e8R1GfbS2XBR3ZnUmrP3lm7WeCcqRq
cd/wb1EVuiEjfMYnSXfa/AMOPr4Bm4GkwOm7zMFavcCZzPpvszA6l4X9hUBf5AjBKIJ8ZXlaNbnX
KzMdijWZ8Y2ZufFNNiaoRLULDoZq2QrBbpCTXipfohoIww45jyP/oquW/VQULClhPlsHedP2XHF0
wvnZ/TeSk+y+ojdof1bp0F8HBNL3+/4NbDyKVsbiW4QTfrsecjkfU6ZwqVL4XAU9KEQyShcg2Uma
Zeiwe56xfsqdcqbtjtbempQFVshhokLHwf21aYmv18eTardI5VLjXY64OkQqKmWvwsHnBtnZG1+n
EFNtXdVyPQI9AH3jG2hSH4ScO9hUDAH+cx6TBw9luKYLTklWJZepl4aE/yxx63Jdc6ZEkmac1zix
1Zjy9yBNS4+XDcznBHjocX0RQY3KttLikBWPpUEBHgASL46yyG2t44Y+qfd7spffyRWo+e7jaXKt
e5tLP9OyWEts3HOL5EFvaLKy2gHT7G6J0k7sebgbhDNlpCDFqCTbqFGGeE2MPQMsRkw+1FEKmxMN
U2/yHs/znuHDxChFj6ipZ9CdG0smB0DxP1bHVN5aGNMRsa4Vz4PbolOTbMY8/vEcCz5mnS+rWNoC
o2l8zntKBwJA0nwWI0TzaQqC9i0jKjgSvNBIWZPtgrahlX1PBx29mibU25n/Foc2Agnt8Oshz6gl
vsPoXLCzlDgjUc/qlypwqQm4VpxYZ67xQMCmp1kNaUDLSpt63wFadEBlNkwtH+7IMUuZDyJfwsEG
h80lkpDRs5417Py6n2/rSN0gCUJlj3ZGSExe83iBjQspm7S8CejHz2A9ZBl2H91ZLlP7KxtfWJxw
VjqbF63rxspC7ecpt6McRmDuZtj4BHjoz6D0BeOQ6FjNAPVeIX5Timh5jtW9fvk6k7auSRTLW58k
Jgdpy609kEucc3QpmNDlZ7JezX0+CAgY4oOqkbA36S3g94OjRqiYaOT2FoznxT1zYsaCFFgak2HJ
goubYnScl+OnMKpCh6xdflgcmK9rHxyYgGFK9klyLXbmWg3/XsUu0tNEXKjCUSCmgcTeuQT9jfd9
TKfgTZTdcZMwgfUrI7qUdl59CTkDmEinTyrLMsJVOs7OxOSD1r0nOaCh/mUJwUEnkaZOnbJ2r4DG
Y7Yj3mFTFsoVvDYDUCstn1ZvwQrjUYoSlgJH0YyrlQt9/sAjj2WrThshpLJ/DwI/NbxZzzXHU9HM
z995+LDUGgHPWdW7gPfoIU5nJ9DWQbv5HwNajVFRvIrZf+Uz1mHpkbue4iA2L3EigtSB/VO7Cy2J
kBJG/5Zuh5jpcKwPkaQwqvh5+geGPZujR58NMvCbvzddJCFowkdtRcLTNZnkyMeSGWPSj3+MWjkz
aML5B4WwWaAnTuRw8cgKhJi0/rjbf6lRYUQ48ccJJ0qeF4Vz8+8SePXdStgDrh+Z46kFRzXsxm0k
dhc3oCOnmDgQJc2O9DTLTaZNbBqHvw9J0h+QW1jsRtQKOA41GRJ14KN3Yhs4onf49yTdVMAtnodC
V/ooK6+8ED8zgGh3jp84CMpuTYwHnHi6tsPKQqB4Z/FS/a+Tt0MMYJO2TTiiysLSBNHqcnGE1sIf
8q13mU0LoIn/hTq+jMmzTB51wFaLTtnSe2zVrFrNUGZzwD0oKsqD9bOprq0O26Wxc40qsCyYXtzV
LeYKGhOslMfce7D9n4qBFuw9ppM2/evF18p5+SCVKop3ptE8pFGZWrnzuLZuap5NzoLv6CA2jikm
jAGOzVKr12QAtiy2hutTjTg3W+Ns+vM/nwKiI0LQisqp1e75iISG6H70JxxhAzN8cdK1EtEZUNjf
0CE6uUZ4Ldt4LoG40B3Njmx55iUjy3/ajIqUgM5fd89Hs8oLkB9kdKXUKAq9LhsuvhEgHmo0Hkzv
zJk8vQ8Rm+t79yRcIXK2KJlAtLZk5+ZjpT5itfKUTz4XCVrEcqzZP0YJgLO5TA9DPesuc2fXh/5w
oi+QlkPPQkOyqCCh9iSoO0s3E7gPQ3BE3n9vgPfkf1FSoYF0Dm4xHQxAgMrfv4OnTgge8sLbJ5Mf
1TAUs/nHqt8vnS73dgPotlwQ+t9o6/w8gcu+LISXqNcycxfC/m35yS6uhH276OgxC6FVr/Kc8Ne8
T4ISOxPvxca4DWgIG9ojYrf+tHSoEuOIjl/Mzwlafb438vlFKP7URYXd3rEbYveeaO1tRws8AZUM
4JK0BtI8ldNVNMUF2ulZlMAS78u6ORvN929UQSC8DCUD/DZ0ZpgbMdfVrXRCnyCWeyaST22UOyG4
fUA+xFgIVGs0pEqMQiiJwuZM2uFOcC/V7/YlETM6kiKmpnZkoyVcfDV93gjosbskkXY1PFQg3Cuz
3ynLrB3EVeIRh7So9uBh1XNT4hGFESbVcrhP9C2wgq+7HTLwxRCSOJ2ezU+Xl4vU6Nog+LdUc8JX
004OQ8yyS51ohETRw2nPV7XKE5mpx5t/H19+nX4o8h46Whp7SOVCrWNgdnP50hbD3cxQRFyh4bat
d1JoEQ7iJUeXSmvS7ZdTxBuLMRhP00StgWeOThAatJGZ7SLrItf2s1PNGTerUs1+9Uhor9lKQWFv
My+upw2eynJOlnWnvO2wHfrJJDODqcs50ZBI68ZH4yYi8XvggPyPqoYHIUqWFjN76QlxfRLfkt2D
jPAdroJZxQR1FNwVOXv+XKEO3/GS2wZVd2Djvej1/1PnHd5i+kFq5JfHdQN/96H1KMHbQH31ESek
hoeFlep7cZitfC3dW03+CLWlPZpO2TiStZfaOFrCY1YD9OscZ9IKHe/RzebC7uOlc2VggY9Kagec
eYJbUwe1MXNTXT5JcvUxG7kRuF4Kn5SwnDlEk1XAxZAxJiPMU7+JJi7U+lqcWiB9gW3FqMcxS4xg
UTPFoeG1vPpZB7FBmmutC/j/LCC9DwC+EhljurJ66b5IrrJXSbnAkzZ099hy9KIusrzzF099u9XO
JRA5WNiXv7AJ6YuCbadIzzNcK5H21xfonZsv9VlDSYidsk+GidAaXE7Z+TmsurbGE4YGdDLR2Eeu
E2Y+UWNzPl4fECROiXLlWRFb8sXlng9zRLmlCozaggNUFOysh/XJVXiNFjHd+540JechqibM3+HU
GWWbT9gClBmc7g4lxqsq4VuzMfSAdLTUzWZTAo1PhprmT7Z+VVpEgUSrSzd0usVrdq2qUBpWp4I4
sHxgRp/rpTphdjshhpsFRs/sOVYK1cNnnoKWjCcnkXmNe2itYeBch+LJJd+VevCQbIoppSwwhu3/
C/xPDlnYEJgFc3WodfqvgrJC8VPoNr4o2pl9Uho86DthLufphyExB81eR+yjaszVbKlq9wcooP0i
caCvoEbKE7/cHqAINP8TUXEUWql+AFpwfIaohGKGji6Go9mUPL4C5UisH/NppKJCknuygs+664v7
FzfanP+GOb2r4mSZNi1BRIE54YBoUYFCL6jhszGazKhx2Pme5OudtCrFZ/8CycDLZGNe38EVwQh4
DtFHFLhfwAWtWXIWAvWV+YZkpKFDGNnJsjm+CtqR+y11uLYGgRlQxBY8/JiIQgxhLOfQM+o6mjpb
DVS49suvCQchjJ/t75qG5sZ/Ko5jBViLBTwJWoTmk0IpgWXzjbbqu/CspeTONmFLywLOMP9og7uE
xCofxJNwlTmZZSSGYi2+GyoHEd0YRUy2jVnBYOj1RFkrf3To+R+Biw+rH/WQ/t3jIRGl9p8KRo5b
JZ61NnXoMtoS5U3G6SA3YTFBpE5sOND81CkVwetg4jqL+ycHduBaIsSah/WKosc6ox/ZCUkTMWoh
eiqG6TMtGkdp3NylPTzqmFcLjgsCPnHkNFqddvjml6Un52t+hYFNG70047B2l6l9TJYNuvNO/Maw
3SACFT4gUcafCTFsHKAPNzh/8/VMhcO2nNsIWK0HQXDu7VhOg7NBDmPhXrwxNaQgyoyPk9CUn10V
uzkMujAcJe2OdBMQFVb79THD76UUHhCsk+/MecjjcpYqoF8FyIEWm0c1kgqpuYfaigDSBw7AVV6B
0hTV0wF6NY6D6D72yA45h2++o2JGgHQQElczuQMtIZfsVPB4EWiNyN4kw9+CciyNNf51YqTA+nXl
qswwt2hwqcseJHhLoAGWxmSePfA2RcrIxWjWONJPzZPcXoIc5Wbzeh+AsryjINiWFBqr9EXp4S0N
lYbPFblHwmZP0/9HwyRt8/RrR0SZqvNCeivT8wNlF2/DNB85T4rLTKdwjyJqBv+fsr7LEbk+jbDd
apqkHvRsj1fcDPhQjRiVGcO7gnGwt9Mxf1mPRoMk3pRb2hSgoXUbctu4kQ1dQRElULRXgRIucjRu
vGnAIoTWD0bI15kAv83C4/ZJXuypsFRL85oDOZuby+OLaN/ydxjt9r+T9AW78Z2VaLZhEYNMbjlh
rmfIht4GjuLD6+IWBh/LiiPuvCpEnsgE3QhCVXVtfUncshcwWsaWdFSiIh0oh1OuvSpPGhvuCCJ/
j2TnCJFpajupDe9zpois1mrIlr4XhQXUHB9/mXPU4K+37tWemaw5Z2exCUGzFLdxeFJUVjZwZUMK
fdgcbWjzdhFE3VsbdJ6DLO+WDDl/ey8rZJH104emKdTNCqGzYl+6rBsEgI2f5Oa4WUqg5B4OlTvR
HEYgpuqlEwCtCGjq2hlRTvIUnPzBtb190VGShGbh7Ki/+ZzI17M8cjjDuReM1IyT1BjOXASOBIcI
THGqSOTtfcwnENzjp/g1ujsQXr3YRJvOlmJls0tkqWN5dYR8f58zkoC4/4o3UhKlVOQ2tgHLtbJT
xCZnlwd/L/H4V5UEIv3TCuB3Rb1DkCKNsAK94jYsAr6rny5Xa7FSC7B6Rtbw153xZQA3YKfBM+Xy
5114iQZfwksPCEyZnDP5GZvAzQsnbipPKCdWDUjnKemV1Vo5pOia6ZD9o0ECEBW8RDo4HEk5XoQ8
raRA/Hj7iTdBQ21l84oEZAVLblLvOAAlZDvptCWXOcNQE9r8NRw66W/A5+aMnGFtTHPPi8S29F1T
YZ4Pzf/OLgAmaw7oP4A4e660ydY+PAXYPyTWgIbcWXF5T4/6UHpzt1tXk6VwgmMUqYhmOgPwiRQH
ybnmZO8qJPmFZ2cFuUr6TrfKZDaarvZg9roR7gailbrJglCr7cM9epTzTcPVl9k50D1Qe7/cHY2L
SKMsEtqfRBbFZYPxn/vAvasLIgua4TzATS/YIZ6XJ1NcGnI1Xf6aeQ2wYBubxqPsw6EvwP4QYUig
nmjMVeNOeQpyh7BWVLrwjgbG999moje9i4dI8CLURjUHVKKATpdR/JxqplTOp4dZLYh6b32zFO15
rMviQvHy1qeivItprMNbxQT8O1EO2TjBUJuBoWla6dS/vasZwaY/RYD5rLxOGxVVPvXC0wp7KFUb
YEKdkfPdZIdSicxY571mT7+cLPQKG295JT2NhhmZJ3MNdVoQ+jODEI6CX2FeB4ZDnysjxZrrNjbN
r8NXdSsoSfkKFR4ORGkdCXzCYpCIAYGQjQ/HkMhMX3roqIPXsmZdRv7TF111ULUQ/pKA3qRTViYu
c/0x/9gZJr5rGUE2WF/kmPSENHNsQRWMyACd2w/rE7EizHqCkA8JQerUlxkXmOwSFFAdDbTiEQvc
+5izZhyA+BnBMnt6TiiMoON6fOLgl+7JqCTiO+kxfWuy7is/Hxl9grTvYn9tn/mkJ26Ty8d/SiLc
MA7bnYdJL9lDqWdR49AC5Sw3CZ5dtrUqj2oRgZ0Hz9JHJM7JN5HCs7BCsfSC5STz/9pOGcf0CSW4
4RO4D3cUiPMeZnqHz7rYBqR6voR9n8ze0xFsrIZ+vkSPvFzhA8XJZM33ubv9L6eu5pJyuBEMdwXW
aGbOEgvMwrpvE4+cMaDst6WGKzgoRu/CYfcI/N2DqOeSb7u/qyqyhxqny9v1MypZmgvThAqYd4t1
bpMVXv6Uesh6xUMjWNIV6slIAuDWR6A9CKZyVUMIjUz6KVkMZFHyr39c0RDQuSCpuKyRbtH7oXc0
yoAaQvrXBmtBWwdSh2VQW5IjnmfuITTdhMceR09btQ3x2oQ5lnnGnB4Ca8+C1vPm4EaPrsfJ7c8Z
M4s94KOcVnb1PMPUvlNp2lLLc3YbXgJJvVbHPKnaSq+oTSWgP1ZprazGng9lM3HrkMgGOZEhuAuB
T0OEVMMI1BslZEMk3he2zVnZ4LVx0QJSvSrlnYz2MwFXj85ps/CPbJbaa7RD60LqNem4F/UAbfPV
g0XC9H4OV3ZlaqrVd1roSS+WpcOg/Nc7CFMJkSDWCzI2aP17M3SBdfA2jB/BWwiufhVaHJFE14cV
REFhA0SgZwg77HlkRBIITCpppzFWWqC/rs3cjQ1jhDwjzA6+8uGQasE0avmhuKYAfK1wgk3D98TN
QR27voopCtBThMwQHOUF78UyL2SBiz8wWgp9bZ5AvUvXJJ5uwa3vhghuyLg61ia7AzMqF3AjTAXX
jM8Np+k9RfrsYJFgCecZwEh0/CNxOJVmKWuYVLpAqM5HO+tCYXafbJiwGXDXGqLhBt1fiTEBxwqP
bMmq6Q7WE0cyB/4/URwEE2hm7T0GyATpQSVRgaUWpLRxn1b8MaEVla+dgeWJzBB6P4ooQe9A+dis
9LutcrtenbeWDxJG2qGh49jKYRvfgewutFHZiDF9AjVXm0sMSfB35fEIl8Up3e/nzDFJRfybR7mF
7RksCAjcc3XbZC7HM3DSFF9XF+7S74fOvengmZqvrwKDP95dLxy2W2GCF+MinomfGFYhHhm5U0Ef
g7GtNGe5JcrOuJRZUZIT+XMGV6itA+wDchS9u/WsVQD6hjItqZx6jkMrw/7mPDqokh/Z1k+7eIJ1
z4tftdPQrUambXWhOSB6ccC0395V7scPdawfkBdJKjZmvR60aXuAWEDiF2i8j8HilCzYnvsQCnpG
79PGUNxayCwmrSgXVAEHLo38vQbr/ulK6VsIWFNQTMgNWiLloNqfMmio88wwoQwVLHCC4tZknNEw
Nk4sKMsnsSmxpIQqb4uaDMMeqp8FwWbYXdgfroYinS8XtpSwA4juqRJBNzCSb29AXgS+GGBs2mfB
dKaWm4tHXKJ0ZGqANPgAmKnteT0AzYm9IpXuZ2odgkS7/IOvxA/AF0dnxemp44smoWCq+Q3agGud
R2LO8rlVyt/o74HSAmVBfWEc0DZEU/cznmVU2cImXDOpmQrUWBxQh+hLUQAu9usK3bH/PmAPXsXJ
l0T+Bn7oyOZOyC/F3DjaHJghXCxb4yuvA8HDLiSjye4FcDmOH/NYOjg7+89fvxvfIMaafXuGfF0K
0UeeT0+Xf0uRvHyb+7bYumMsdadLvi2RDYFqASWowZxXuqKTXilORg5Dn/WdadMKVquhaLPhaaEu
bHA/S9RJwRn5tP33xdPAnDn2iCRxhN+hrliDrtBZQaOBMOFxrUghG53HdOiKwDWnOkEZYbOHHAG3
5viu4MYVrlCdgsZVk4GllrJWwdN/Wt8OqHWTvOP96VXiVxxFRBZ04hqvUdbkx1MnUhhSJYIjnHc6
AvMEPq5jDrTlblD6BcYkuDGxj6PXxCB1J7PFdlqoFB4vkHqi91gx3T8qYoP1UPm/CVizIua/vmEH
AWVz7JQyQv3AjXmfX9W/6TCRRrU3VO+rhB3yGfaElv6g04g9dgnhK63FCE0PcIM4cMdcG14b/InS
FknrqTzTiGJqvID+ECrMh6pHQr2kxlK93O7LucbCIX+ogOefC4QQQxaXHP/EOETNzxqgIZ8J8zh2
PCbZzrhl2CCng0xdlkMyKXLKa4ea7qEZorIBcf4vPPmAIhNqZDz1pm0IScdR+2GGm//7mzTYwlH6
zIiQRRN8VRgC3rJ1LURr8gUvLqzKeHxOFFSI3jbveslm5zOtH052SamGMZxQdkAoVjAuHF2Tl0zH
hUdujNl7AqeCXjPkx2JUfhCOunpjqnESh2iT8oaceYXpGpDCZdSXf/IsEnSONPN76y16Hj91IRoZ
vub+ZGjEpp0aOg177R1MJEfOmU554kpP+HdSRahHVZ3kfQlTNBX/V8oiHZAiJEqWKNB9NfF/C6cC
bGCeGYJl1WrRsItrKHomW0LogHVISmhm07lSGE8WL4AMKHcu3qY+Hf00A5W9ENoZFoUpOBI+tfzv
o+dxcv21CuowRv6qY1lNyHmrKwGinKsb6EWDhjwvqWrkT52k0YwO7eZoTe/G8XKlFPLvr8r++Xga
wtpJ40JPr2Ka+f4J8rSufROHENgCILeK3jjXDwIyx+9wxO5zdFsvR62X8yt55BbXHSfvJQCiuYzP
tqyaeVklmZkSPsooYX3B8OvpZuwMNyux358FrDVWP9qsnq1ZpBr7LrSZMeAFjqT4PgY9rqp2pxCw
cfSQvCnvcRhDN9Q6GVezGgoYSidAXDQ0+HdQ+KAIXfBW94aCgS9aToenej3rzdzxhmnOfts9Ek3Y
9fkvSTgqmRIDzFkEZHU0vTJDER77Bz99rejAwEtWxxFvgvEAmKYnury+a+Vm4iPkhKiyVXs/VT4L
jRY4SA9+4YamwyYz+wIgFgO4Pbys4O4yaBq9OzlA4N+X+GDUziDYp4e/suee8IBeVe+UpLX08gr7
qB4ZSGmbdyJELNbjbDqKpTXajQI2FuNxM7xgj9PGDBmcusx5B3zCQNvJRwh2wxLbW/DLPqE9/sti
ZDMrCyAixCMl7S/o23WuiX0R/zuBCgi4lF6/XgB/JE3AJBA6kyvfd+oRPEKWT5L91x9CVxuvHPTN
hnQRKSimsfd7503dOkT3SpY3q6zgSKLYtcw9Klh9kL2oSe2fDlJarNQ953cjpZ6Cku6+l/wFdDSM
JNGAKvIKZIsi3eGRc9qQPd9itWvaYByoYhRam/s7W66TX4pLbUr9OI5R3zlEzf2fwJy4pEC3ulzV
bbxTUkX1lmIxGuBDt7YzJ/vFc1ItDZMPVL5sLbFU0cQIIuT9laWbFdL9vckPp6v+dipy5z4rQBQM
XfSRKCl594a7vcms5Yurq3T2WIbj1+j7lsY1e+mPiTA3kFTA7JwmwlyIDB9W0+bz9LvSRGeZZ4s8
jLSaOhtxOouoB4Dt9awE7bws6Ugf8AlAZ6x/erDcNJ8xNbVso0BTdV2PCR6AaNHdhva4i9nU/ayE
fF3GcHb/YLB7pW4TGJ7MTxNDtJALdVO5s+9MBtYa7wr1n5LJi2h10moXjod8bELh0iBvTWXnZZkm
hFS1tqlOs2GiPN8BeGQWbm2qmMy7EZ88V/Ch7DfrKMZaXwPYTDCGSqmjYNRNI2Y5Ytw4jpb9dzcI
97mFQcoqNtLTlkYTeef9WCNAAtuu2mbQRCedFJoPmwDR93lmrneZzo7JBIJr7E0DYpdXgWPKTiWN
2Cz8+d9ccgzZSN5/SYOUjuAwJr4sX2tmtmBFsdHZzIG3+eCPfQzKpTWruK5JbyIFOoK6lkBm9tgX
966K15CB2nfgyq9d30gNl5H2oEG9uctlzVYnjQNsXlMFtGNgtDqVda06vhj8zNnVElyuqrJHSrL6
uylQmV3sCeqpsv1ZIQUmCDHCR34Qhz5V+9CX8atD5p9qrcV4L7gMmBU+Vrth02N94UG5sBC1kKgz
IbnBSeSkuFNfLqVctS5ncnM0C1Bxc+iUMlbSRsSjWSa6/gB7fhExku2XlS/dp3qvTvd4bTbi4205
Pw4P+orOC9IOter4pMedOkNhLt8+pa25KXWszDp2lqgcarUvgfQ+xdAnerOAeC7bHkyrZGlt283u
15u/4YLGe8iOywq28oXRhK/I44E3aodRyoXQUmrpUMssey45t4GJW5WmlRkp7OOHYkgiuHB2G7Ut
wp3N0nklgCupBBG4Z+/QgG+cCh9ZpWbPTxhpSEAG/L9psoT0akT/DPG9+0U4yj3qbcpIe+jf2Eja
KCFBHLgm3mz9LpUpNvEE/jvNNSC0oj5rXJCYXBcIjkZ0VtmelZu66THYh0PJj2Ck/WFmV2tsuVwJ
8HxEOZLVoZx6YsnYO+7BHWpaFwHzEcALxghJu9b+a5q2ILyYqWozw9pJfjyf6j8ZeawrL2ZPpHTs
FlDtzTwfLnt/BnQweIYwaNluiU7z/nT2kdEAOCZuyMx5AAZInEICUsFBnfOlY97DJ2K+OCI3BbnH
sX8S0grSgaDHP5Ai8age+YZntAqElTllfFpHoIoY5mtsbofpGeqvd6g1SaTx0YAaPLR1cnUStdNw
J9vbhRzvZ6npseNEJO+mDvUqYs8ntCKy7b/olhUv0hXdfJ2yg5RCVhEtWBuBLh9Tq+5sQ8fyct11
/u1GSFJzJg9wV/hc3/0u/1zkhkJwN72R87wNpztu/5GK2t2U3hKWICSFEobX6h+EuSRU/XFRn0XT
2WBlzbwHbUQPJ7SPnG43DMD0lGgFUaFlTxW14GGzx2tyWtiZNBia/XvLvkvSfJCb89v1Rw6QevZA
n9rb8uEZswLC3WvEUlk9tD4NHVK5tRhFY0pRJ0yCYg17/fZpv/cJ1A0BsbrMWxEM5yh1DFNs6HpP
S/509sLLfh2n+blJ0q/KHkaPiNV8Nwg7dC/xkLBTsbFsoMufJ3K70qs/UGP3a4X+wo8QEB+CmUOv
xCFHDhOHhvC6mjG7LsVAvOnWLkl051gXUJ8zTCGvoTGtmIZugKP01o86aTPbp6o/N6foRXDPe+q/
YyXiS6q/f7GgW5rvXo9f8xX469nQmGCsIAHqG1oORsiXwHGwspNhSyHdfWgudz792CQHRmscLoU7
UrJBNHso10Ngk49NvUjVm4r736YvEiEEFqlfHeujoHFgQt1dJ5wtUbfO+deCLU2IgZPmjojSM+N+
i2PZdJXuDYCaxXEYTV4C672grFaq2KaxTk35T/QMruWFP21L2nM98bETGcCv6J+/SXuZv+EbO2XS
rnXNGNjA3hhfWhEiOyU2/HBlZKDKp57BipgFyNH+eHQo1AafvpdcrAFhaAmWD5DuqYJstH0SiLHv
KeXxlPg+nvYAHtnfTd2tfEgyqJTTvEqyZFjQGAyqNXKxK+KLFBnKLevWlVYcZCEPm1gE2mknrXK8
sZ+e2bwBrqcGCAGej/mJze22ksvhInc4jOuA064vEC+S4eIY17i0qoErdQX9/CyQHu3oRJT0KfV6
HjcOba114NRIQ5lXXJdmc8mV4m9TlTARTprqE9bP03dSOFwLtTlKhoVn9lDSJGhOlxE/lUqFpxKp
+MvwX8wNJkt6VPaO8HlZwd6Yh++An+TeLfBN4IQjeAQ1PLRX3bSGdtqO879h4ABzitS6yDmhjcWF
nPMesQRqz0LtrOdSIDcYwt/IuO7Xg0SW2wDoaAS9XRzDNrTpP2LbNJLcWP26P66uTXF7Ywr92Zna
tLSB8SFGlT7FVgngq9JHrsEkvadgE/jhqlEJUtLgSAaiYqeAIdojX3VcXcvNI9IFON7Yzs0Lzq20
l24SalFkeHBsfS9pYpGFv1I6fGH7hIS3tjQfF7o7resQ3WMqyufc8uXrXC4OLrMbfWxTIR/vWvMK
dIA7zpsuhEpcwN5r0qEYk5SEg4ByhuBlyycwGA764rdCI6Wv+Kna/lBWCeWfC/4vCoa8FPty7pHz
88jIfahBvt2gy/lUJKLIhqvCY0Y8ilobwDXDfLg9ryPyzB7JNZmYZpBdudGQAOfciu30kT/Fv6l1
3TQb04ZV+01RM6eQ6RTo8dIJwdmWSbX6AyjyKVSx1QPlsYzpZc3N3pOrSYZpMxSo/UYAMejxZGXn
bLT20vEaHL2BWjPh0cukPYG0FzALumm3FpjvjGcpPjGO2MUTnlrAYS7r3V2HDVc4eqTvQ+MdjmPB
hyxD9UlyZ5D8Lm79yvxBLJWdPkN65szl22iC7re78Y5xq6eukExP7xFETZgB6t619+g9HSc6hS9t
PmfjB/hU+GZ3dXc4kITMKM27rCkWgSJTMzw+8pE9baWrQ0J04wI3cUz1m2290HqPRlchRGmM02ud
stew/xIaODsJoMINLXR4PtOAr2XwtLufwB1rCEY47uWuIT1whFQ1h8erGwGxtYDQs7PqFhlVllOZ
RaAXP5qgEG98xeIsdZCQEvcee+5F4GX72shP+eNBPWx1Hb03pFD4VhHOLlxa4aSoXztqIQjlxrSu
Cu+swdurLchYzHhr6rZ+6S5AKKjEavG+PbgUTrKRdiMJjhAM8COYkP1sGuF5sAgo7e9II+yPeyB2
td/iD9/VHqHk1YRInQriZDdcN6CYd8IdX1zsXd/yAdiOzLpXSQfXzTrR6XZTWeDkuaZ3c5D+JwHX
LTdcE9EB+Ym8WtRJ/+H4HXotudWA7p8nQyh5cVjgPZMUDtEzxMVlKgR+EF8u6TNYXp1oGbsJq/FB
VqE40Sm6DqKWU9asA+Wg1bmMm1KKeXNkUi8cuZvdcM2nAjHlAIOHI//odZxWA8Ih9KWiqxzM1Wnf
7hC0QwR6/smp3Bmpk0EI/AvZ5KtFwTfyk7lMgpRwTVP5JVzkxCIntyUiOr6+0DEf4a2VUPH2bUXk
MJdktC9lQHT1eOQ/KYXTHLagRMByHV3Be4+xIR041MowQfd/ZojvsRdOvNPl1KtAN/f0yVjc+DgO
FGxm10rdVlgvhG4ncyfrbBl5+MWGsmVNgmKdW7xgJa39hxMeqKPA9znCoUyLdAJy9mVznFqJb3Ok
8gHdOUuan1Sx+3S2z5zEqg7tg7Mz0oKMwuSLikWXutCvmKyrnyfTxNxoL5g6P0C3vUYLMgLDipyG
2HM0ymI1PFOr9KaktjZ4y42y/17/auuqCY2r7boU9V1zM8Z4t+sD1xXoqtSaJ1LBzKVrInpPS3mn
ITKCoS1R4Iu51veBXY/1d9oG8JlT0408aSgBVxINlEvY4m/VrBmzoT92zSxBA34WPC+QQ/ZL77H4
cd/xKIZHpOwsyXxC7zXntpmo4J4zg2yHjIKPPJM13UUB37Qcbb8ICzh8gHi6cluNZ6mdmen9JuOz
XM2qn02mI17ttnuBpDCJXCjGPojqWFofjIskAjhQB4sytbCgEsYgqDsNnnYI2Uvpj0c5Ya4fKpfe
WnqVZbH4VmFt8/UiAOAxSwGompqRN/POGpM91XWhl0S+uVtg7XxWIrx6So3JpY6fSyLZu+1Q8cfd
WX6HrIL5GXzkNykjrBCoylpOQwo48mE2vJiTbDfQjmXnpSOHcYXXEOpZsvnVQIalZRLiEWjAdVC3
D90TW8LB2RaTZXRrpk1yM7gtwxBnLtkpbLCi48tFUVJGLXNFRdIWwj/DdGylIPc1lql9n80zfBtL
n0vMxdSQ3MBVqj7D3jTSbX+vrndZjBO2G4pudUIcsdnKMwWr/SjR46dl0pMirTbElMfikiy3jqzc
axnaYDs/iQJEEiTyPRZU3vU8Z8zbzVvFi6XS8SXgSl/GqBAo2k9Wvji5BTPDi4FQPACC767VxddQ
5Pe557ZFbj4ynRyT2Pvo/1ji0TcTgpELyGg3sWxYmtEF6NtG2gztt73zzRsmRPtPg+P3TEOsD/tv
84YOHNmCuzFY21qEg3UzlpIjhfFTWDYpHl8YsdI3MeMj1aGF+uuQxiPPgiGyqx91VKGE5TFd44Y1
SPQAXPbzwD8GklxBM81Eyu3ocO3P1dahI/yiMT2FpSYqZQ9Pr7xoBYfTUhnHu+VEOnr7EWJmOc85
fdOFUGBr4rkxRyQzCB/Nc1NqjXhE9H0yxPIPfTFwSK2fhJjF08O/NIV2v3dHU7bdU1kQ7CDa8Da3
2+AX2VbtveHq9wWGtAykHYDytvbdikZJr5+FvSSCKELcoHIOG8FLwF0QB+ezhdMCQeEEEYvQlPXF
W3lP07+MZuqSQ7NSwzwPE2N4Zs66Hjyc5j8lsaw6NrbCnth3gSpuKMjU2VxJ+mAJDeWcgDv3VjTv
5IAyuLoo1gz+7jYb2VGGXVeGwFS+SqpnTmLrHrlptFWihcxc0hViPBPYUqbf75nSiPJEtrTL6Iaj
3fuLHcNsaI3CMHZ3/+AjtTf6mv/MZF50QxS/KRQFLmmAT8dSIeoVip3GDHwBYcbUHgipYp5iLt0c
ipxHkyPgiDRzirz2Julot6dLP+LRyTh573a5GdidatMnYh7jrkU/HgJdz6zJghnTEBMtbwNvyjZr
vsPtPQEp4tI8bfBFgzYspy5WL3HcZAk5kScVIByJV/I6o8CkkyTY+OybAZQBgkMGpc/OyTzdSv0p
Tg+7qi12Ht4vIO/1Y9OBn3GbWPV6OSBXdJ1adOi2gFW3/ls79BoY6SgPtpyS/mSznRzxsih489NA
pkGR6BHOdcAqbx5P1My2KmyJXrVf5kWU8qo1eZPTDIvnjK8NmYBb/wtYH9ldiVGRMZCT8pG8KsDF
ajev9GyCyfRMk3cjo7TL3Bd3NzlZWdy4kW23rer3Af5UzRrN6Lvp6g78UyvmNUfUackOxUnDZZiV
J8Ns0AU46pnczgCIowdeopDuXtFkyZXvtCHD9JfInTYWGrG+QNdB9X2wys+xyZNlhxbObdWAiDwF
YMT4bIx2KJvEdnz0/znqq3k3rp7bQxpTh2KrubQMl8Zr3klUZZq4V2bF/ALSfGe2KskbVQ09jkyf
GMABQKIlaHXgw27YNSPHFlFwI+AucQWogmVZVUNjos4CIW+A3mWlAnVWkk37Wm5zbdnmQnGhBLVH
9pTksudkQAu86MTHlPXJfcB2DaHlruqqiWyFDl416Lbj6O3qClFxRohq8XUGaP0FBFJLUVW4glXe
z0Fgj8+vADWXX37bOpIsXQndG/wnEh1kt3cYUw/CTiEjKmymXP7TzdeZwp7c9/JxFwuvCvlxYnPd
/Yld2IQAnuA5yPktSvMURwmmkjBbZgaw0EOzXU+vjbjW843XQOpky9kiWemUowNx0ud6nE2wQyV+
mQ4RSRslYHoiavyTRTwfzrXXf0prJMbohABwUWMZEjyogVEcYg4O1NSQrT4csvXtUsYDTdFmjq4t
N5txpMH8/RiDV1AGC57D1f96pJYGpXSRPg0lzUThTDxphM2Wpon0WfttqCuRLLtXrCpjAneabJL9
SwgXtNFcD8E5Bg0i0lzpsltz92L5WjB4+b+7iMbqC26xuJmnlK6mfem4CXgWfbVmlWqmr/jKMuTa
ztTK87ZKzyI6Vo1ZP2c2sFxhU6rE4koTjK1Q107gNDdud4ZPim34Rg4/N4+sMW8X8y9jwv5qZJ+l
Nj8+95AWc1bxVy1qZJSn8Z85te+hy1ZgJKQqYXP0BMwBHsbrmwFBX4HsdZx/iI6iz5tkNaVF6D47
QKLn/V+oQS3QWqEXo8BqPyHbE/dznYQ4tGVb2//KmuRG00x5AwWLaw2kpS9/Jng/2PxhOe5iF2VV
kQkmDEw7QmWFajC8mf12NgU0jp8cixzxOegnLdX4X6HGk+/IvJsFh/0f3Gvbi+OUJjsTeLOvnR0K
qlDsngutxlUvMAdrZwMTfQkTUdNaTRhFcuXJNTyd+3Ppmr9jETvJmklpx60PjDrRABK7OwpgPcTv
qZN9tDX/qNkeNSMyROKNwCARtT97hDZpRchJmyxfNx0uJz9xfSeNwDLMgMzInuvw+YuR7QZI8VFA
lw57mJQWnjT12dbeWlxoaQsX2c0lK/heKIVEl3kQ2+uTtD64I07FS+nFUmXTC+m3P0mB776v8HN0
wAAvZQneuLi2OqFLgK88cV2WRRV7f6ftS5ZvMJC+13uuG1Z7XBFpe6SgnlDMz3m5XZtPjyL7n/VE
vVn/y4fnOLW8TeQ7MvDLxgBZzUkmV8KMdEn0klErWFVlx/kdkqfxxHT77Y3pXGEn3fXCd7XyvUoN
1LoA9LQPBYMcFZmIhmKEm4HWXTaINGv5sqNc4Zog8rCSSXtoMXPSRh+ogY/nlpfXJb9UEfReAVkG
m5uWNbWvAQZdJnWJ4DQBeTiOmvInRVV8jUh9wSe9cUxM1srsxu2lfNmFrDpBQGjfwbs8FGhbcJkP
MuOsNWvRsJywU3sE5Ce4EC6Carw29MJV16cSM7x71/N/WAGy97pBRDCnIgOuZJgJDfuF6OXAFNWh
4VC/9HXVlh7xxe4XonsYOXVLBCIIloNuv1LCgGCDAfxy3zB/3knob7XyKPLZ6qL39OOa723oWKsf
WKf8MPlTh7bKlRrj/FlwL5bkDO1AQzQpqnsFZz4kxrKZhMOZxzUo3ZXQJ3IdbdKN7vbzi8/fwZ2V
ZWtwWsJg66K3dcheQ3j7mSm6+vd/eW9CVbxiNCsdnfmnuBPVdNBXljQeIXgAoKvEu6Ng5/2xhScn
IVun/JYlCZzF0NgP74opmMV3AIEGqOS2YI4iL72MWpzBN4wV0D6OQI7Nz/4oYaVrJG1N6FWaHZW/
Kldoi0/ASOqVg6N5hS2o8022BNVs+BYbQKRJxiYWET1ya1imkONri25Q32tjiqVZP+RAP7wyVnVg
2sHOUBVmwud9Tf3m2ce0Lf+1Rcqy1iH2Jb6NR4swD9HTPdSR7UXjG4tbGsY7aNCD7U84w+hwarIp
oa9Mu7303OyJ2iiYYTpcg8zw40EesyuIkJv3OuCbyfuqQn+/2DlWchWe/UEUtKWI/dtK8Orxl6vV
qk4pxgHPoZk77hG0ZtSzbuEeD1BQx6lR2hqr4bQDIgQ/Bsn5JB9F6k7CwVhJHlhb2C+h6MePyCF9
2HjjfUyGVTU/WrjwJg87H0WfWj3SMprUb3miedTB/gxiwqEXG+uTCTRJ8syZaxcaO3l+lKgoCjHg
Pc7t9ExvttMX+Rw0Lf9EDY0TledePutL+kidCOh1E60tIWSAcV2xRbf0HyQgq4YHfpXkECEzTwAu
yJuKDEgwfu+RNRqB+cqpkfFNLQiTbURhkVBBDwahSefnJxDENXzYGtYCD2tLybutwD+qZimO3o+t
NV4C+/Qw9RKww30MGPOpaRIu18oStkU5OWf3rFPm+3PcEWeAngCjsgfVsLh0frOG3PxkTpp1T3AU
ItS5VSqxeqr4bQEBzQTdJl1DDwFmByuQv7eRc7M4khKm1Gajs957YeLhYaTSkUvD5RWRvO5szLBX
H7resCN7lo6ksYToxPIK+qwowwe5XR3DrN9DlxyaNgcS8dl0CV7LYWJvKJCcemb2jvC6mrqRPMS6
1F1wd19vZ+xZiHEc5Zfzmrj6a0OKVfI0RCT061eIrXSloWyS+J+PQ8tS9t40ggyeDKFglt9diOb7
8b4qcZo8BbSiAvuB1Y9wM2Z3O/5juj/taE1eAT7L4YRkYVsQsSMv2rXGam0wfhVk5gmTRzRMe2bK
Vh7/Xc6jum+V2QblINpVNeqwx/hNn0Ro3n5PVHN4YjShctqX8Tnk5T9u+gyaskwqaYkLxJ5wO4UJ
VTwpH9vziGB0fBp4PXz0C5P61rMRlIHz3sppAh7sJToky4WoujdAZydZd2Es5RANNZ3FPZ0cs7KJ
o5uMCbX2tMwbEHIEAaT4YwrEcq9uHw1Z17kA07HkOVvyMf5QCStHn+MX+fPKkhGl4FtyUS9HDGiW
xgQCKVcDpYmMfxKf/zHHkHL1PY+0lzO0Ah75026ewFgjBfw3lXfMmXc+44HsDSt3XWwnTUkZeMTA
JVoR0YOSo3/dkspBMDLLnk3113tzco6ZGIeTX9auwoXgQVimq2vk2u9MUsjkKMuarm2C33YebqIU
zyutcfWIPUwx2gigTPN/6Jfkkw3rfwVot3Pi160YszpnDD6DmJZGRxNkCTRi9zw+WcONTbZ5kjM0
FnFBrWrvrZOAWTzTwF4X2lnKGqkujVT4K8+XXy33jOr8AG2jId6h7sGIs1mWSWrvhWnVKyDD58FD
c3S9ZikMnLekftSNFqmEu9veCaqrgxg8ty9pISinSlpnRcrX3BSpU0TGuG/P1DAWxZT5NvTjuGT5
tDs/NxzNwncsCyS9jpM/yAN9qgEPpody2tRIt2ddbz5VCobkC3qHohLQd7jsa8kMdMbHKfVA3biS
YE3pntWuOES+Q3ukOZsuF7v48JERdiwqSukiJmg5GHF6nMmK2tt8UAj1pgviRtoegYK5XdrAH603
lLuz7KH3ZrXiPS6tfTymmjUwaBCUqVC9NPNwxJmucdQ8CYUo8qZpBs/S+2vAvriVmanLsR9hRvrr
UQRHYbTmZuda6CHGxaek7yMoXPlHj5Wfx3IXvBP2D4YIi8lmECyvxaOfh74seiHz9KnEWH+jx/1p
JuyyfU4zrLLwt2YwQb0puebHP24niywhMd8vNt0LtdLTpX6A10oS4hqxoJVkphEf/3+3C5D+qBVQ
GvpcDPgd9warji/rmLn7PmdMU3QJOajb+t9DXqw68EmoXCTC/kKZaNnYVcZ2W5/6Y6tmlZZzKnHJ
8YK9eyRFh04go+UHimStXkt6Bikcr1bp2nct1y14F0O4xuz26zxWUFse2Xn1T/wJ1a8l7CrwZcAR
Qsc5+cE7BbjzzoZ1Tdtkdkem4akGg74YFpf/JhPCt+x0shL6oZwjjZCEgBvF13kTlBRgfRZBHWu0
WoJUJpN9DKY5simSGmJCmzCAcDdktCTL2T4fYPwvHkdHvnQEZvLuW3ODYIYJ2xKd0kmxcPqAirLe
DtY7/prAT8nHI4m8USc+yBl/ateMOLILmmscdR3c35ttpzuMHdvoj8y2YNsHuBTW/XxsF29vtibi
3pUd6tZkMccI5gFLEJKnXyYHhASeGMAZHm/jl31ThllZS9RoHi0WfoeOikC2/a5mvsQ+J+fIux/R
caWvUQbJ1Jy8Ryn9kIY6OYLmOUXVmYZ0mTkLElYX1g18+uada+Bpqe0anmGG5SM5FZ3J8WeBLN94
kCqW1clwHxQAsK+2kmrdDfG+d9KR3IsUJPAY6+2Eq6/YGqIyGkwk36BQh7TPm479rfgJwLUDIgXV
bmgtJeHmM4QJqe1doMUkFPO5cLGvJTNMC1FEGnvSAjuk8xDpzrVPHaV9zWxxwyUiTYv2v2g5nSbo
IxwDVsvhqNDc7JdBkkX4oYuskUNwtyLI3Q8Ua/O+B4Zss/NDqkTJQd7twaOz0e/adLmipoaxAdot
x6ZAQfxYF5/X2Oco4BeoiBkeOy6aidBtRqXGfxi0ZmAkibJNK18ded0Qw79d5GP+9PJ/6fJ6J/16
uXY+PmV1lsAETur6TAAEOSWnY05gpOsLnvtU7YVCQY0SPjPRO4wRfV7xTF829Ej/C290cnXrhRng
mMSqKhBqSfS3nvUQisD/ve5PVb01tYVjjT2fejFnc0nd0q1XplSkZbErnKeFrK77cjbT5oV59CuM
HB765gIvB+88qHbNDdAhv2/SE2xSAV+V85EDga37gpN7NLt7y2ZeGkOK5cgnh/PqDTmYrOeD0ox3
4fffs8F6oGLlpz+0lQSOzqdinJ5fjxCbdLSWaVt68vp8MYNvy9rEFJ0lrfheqDgoMog6M/0cemL8
6Jhj7HtazOGFmW8h0HjvHXKcUPgsrtv6v8udqQRjegKEqqL7xU+NAmvSzAwfDJChYh9wazzfCjYM
3ZzxsY9sZSn1jPdqZpXHlZz2xw5emuA4wC4obVJIuKruYykuBmaNEE7H8ppLqYwjP8lFbduDrYiF
hDTt3ANWIqrkiHZyj5z1t9pKXhulZYy5g4ZFXiVtUL5gjxTJzf4KPptuU8nErxt2L+nBegtdeZf/
HlSVUy0kLbKjK4qtFbfeopBWXkQTXKwHYCT2xJm/ydW9SdOQvnXwl7IEn21Ncs3aEDt/V+uzwtDP
aazUMkVRHfRSlUYc1oezKUIoiL6561eKSjSqwjl898TMxLAMrS1LIuS4AFokvtqnr9yDsedCFTjG
ZlzOXm0OtSZtTZyi+nAqlKWCQNGyVsYbBGg2j7D+xyS6tVXVKG29HuXwXj9BY2XmPf0qL8latLun
uLoqZa3zyfhcZt1U9h0Bxbrgb5Oyg48VES2eXd55nysXid4A/8N6OgCioYsYGFTP57MJqLBF80bG
7Pn4gB22je0380Nglqd0ykVjXZgoAajQUHfQJz97rryk3iCvgcnguxnPP4MawYfyAqVHHHyWRiig
H3lLscPt+a2ibsmTpaNaqWFFYvzIVBl3I+t13oZvXZcigY3Ei315/Hj+Y3zLlTFhzWUFz4VJIsZC
TQinxLU8MhQNceL5zHFhbtTWvw1S4JX4/Q8Eg2oYkLhHCNkrg6MLJOa0IVtaFPBwfQ6R2VkkmiGF
Wxfuy1Gnj0EB+TU76XmE4N1c5fcKBwXR5ytKVAz5xQ7lIIujsDOBNofd5oans4FtHVLbW/7+qbAs
4Mxoqm4OzbhiZvlRtrSCk1zybcC9uBvsjpwM/CdHk1DwrexnAEXHE9NNlBBXr8ECx8do2irTI+pB
glV4FRndV9YekI0QTO42/BQaB9+YsVi2bcos6QZzOr6sCp5U3jfyjIU45FJD+2Z0G2lIQI8OUqUq
E5kvS8hdSjOa1+qAZ4KJKs16U4Ar3g4/ZHxy7nbUOCMRqi7J9nFg3HvLyIJzM7+eXKEpjxhR0aPp
54RgInJgVXW6PuBwMp/UsWfGqH1QYRrPeRFeiRcEDg3b8BgCscyTbrTnwiLpJPcIdWzxgU+OTW4j
oiCTAyqdbWmB4o/SuqfIj7QD/XZ40E+HgHgdhnCaAs6+RfVXSKT+HkPt3hYKiRFU/uGbhpkjGG8g
qLyG/atUPQUe1PpYzXMzFbVDsD8Wbj+zgzoTD0/JojaqnJd6tZnyBP+h14ecXABA6lFwrQA4L0yP
2s3I2r+wM49WcJX0BqXW74kXNYxJ8TWsSdumrhiPCzIMmdjjbYzr5Ug2XH1iTcKHjYsoplYNQ0Ma
efV8Z5ZsGI8qkkR0FvVr9j8eltm7P8KfVQ/ku0I6+nQIBYBmfFSJQvuJ7OyNr3vkz8MY+m/g/GlE
F0KeSJ4xDR/uBfwK9523aN1358S7TTnUcGUkcV59evbKjMbaii5BywKiVf7gnK7CE6TFEAD0s4hY
1SnBfuQLY7eUdcWOoZfcVzBefVj29jH00lETObRHLgN6adpflyUmxTvSekQu49JJptsTx2bDmI2C
pUXnR55s2Wi1jIOj+9F1ekHbQcVGzxHZAec+0jGSN7r5Bc+nYMCuvVk5UvNtZ+u9WIFGwSoWGWiD
U0dmDXDNaOhGWdX+/zA3rbTzoGgIRblvGRxk6R2/aNAyo+MyfLrjX/dOwmfmeB5AW1g6xKvt2Nbn
ggxa2rATq5cLnKbjAdCVb349MRbEQWI7+6za2LckklQLmDeUz5yGJTz7uHkL6uqIasrCqaY+Ga8X
dImUfn7YUne/LA7ZeE80Bi7D7EuR/DnzHbtOpNSKvgmjLa67gnKOqKMfEWmKU4apOdllk2TaYUVz
y1XT0dvp0tbjRaf5xqlKREm0+CtQRsqIZkgkZQtq5txMvZdiDCk1djxnbaBsstnsa238fKtF1IFo
+kFJQJZ3mUtSSLjtbCf9ZRX42Xlgd40iNk9Gh10aq7uFSDRRN0dX0pzlDiRm0XVOuU9xyDnbO70D
WZMMQidPDX1vx/8ZI7IqSlDvi7XUwJuBauDjpTMz9UIRE+qliTb0jmyIW2/KNxRAM6WlUHslg0Bs
mf70B+Ceb0qbc0J/44wS3mFGbNj5pM2N5BFIDYAkn9dR9z0ZZb1ernuXNrnjODXpFbm4HXRnP5un
nNWI/3P8OGHsNkKsYJXj6mCXfAhv5EBNd8at7Uh+Jr/8kcszci9RWAOTa01bMw0j3qBzUruYsZbo
xNKU5V5sVrtYHDQr10wk7s0+Yg7ZNnLmGYTOewk415B2rPG1Gn3A0YHJmF83W8cQVEUSJ+guhVrt
qaBbKIdGsYA+YWUvphjC41PIxTOQL926xaWCEO+B3ssi+5absuj+j1Q5JK3/4mqavcBX1NuPI/vO
KvwEpMZjfbEBkRdyE4YqkgdNQ60fp/tbVGIXet6vOI3ObhA1pf/MDPN4Ps7Ty15eM3PSIFEOQNnw
Sv0sw4JPiU2/kaq/DdE7LPW7bcyTOVntuuyt0rmHK0f8RgM08mXNWsWkF054Ga5kdmcPkiNHgTn1
VEuv6fJBtfay5xth4WAGkjH9Q5psbwnFrEdwTJzjwC51w5Fabbk0jMpJr1mXdm5TnwHQkIPTCQR9
EHpI+L906zpcFGIYXV8Ba5mlsMf29+YNlHpuakIeDFjYwGowIJwzu5tPI23Il1ZhK6+dSM73EE/B
xKIbYFp47iqC9khbSFyIwxmFqC3bV6py8WJA4f/ZHwrpZHgXlmtreaJWN8rwXQ5d3m/cgxx6lf+Y
uTB3P2odZI835cV6T/z3CnSKXNpWmEU5FY54r02Ak7+FH7oUMv1KxseUBgWdycd5VgzkNlOhYeK4
jq69I8LFZT+3T0PcuDp3nglNBcxrDCBiDDjO5Iug0OLObSmHJPUvVUVWu5eS/3YIkERMmH4n4g2/
PvPxkewYlzigC3Lm//+NvnacKHs0o7N9GxrDk/vKD093m++nmY0bUAh4tEs4ir4WYElZKo+2jm/j
DBW9PTzjDRZpWQBMmXda6sQHntoBZYCBgCcQyDvd1NIiE5sUZVNdfDwJvk8e0X34tqMxmNQPa3Qn
QIJIAm9EGJEQg6rY23+ry7WmJcrlpTpkVIMLfp6wvTP2u8SV1yFKGaSfaS3qQPYB1lPJuKlJ0LJP
IYHmCHZw60iG7ykoxvnmZohgP+DMN7/W/2AhHqgDnCfRA9pTK3e/TieWdBi98O+SMxhwca0EEBoG
Xsni8D0P5w7somhokEZvV+qmULzNpcw/iQ079mfdnYQlTWPwUCycpLiqKqXPkUXlEnnpflqvpeBK
dthpqTqu8NGr/Xtlpnl9RnvLLCjpJSLJDP2U1DgAigXhYnd5TARnaT44wztvrZ7iwXxrZZP47tPz
7+z3feSg4jwYd4r7yjGJ73QlFb3LsXqiw8cOmpkW5c91j16Q2jpjrFXMmEAC+82u4soAU7MsBLBk
CI6VbBgRCU/Bvu4faqWIpRbfBXaUhAEnj7Wc7ldd0Gg1UaTNagZtoqpPo+78e29BQCRS07pOYSrv
R8EiTbok2yKTyBwdNcY3/M7r3GaIKc6Ggk0M1jWNEth68T7aWaJQMkY0RAe+BYBBCW878T1io2Ix
1bWpBTbDuQRhH8p/K3uuDHgyFilO4xu41+EidLsEAAhjdNDSFx1w+wtOFBq7frnT4XCn39Ge+UbQ
DNW/lZx4nmCAa6c2rJUQFUJ/GLsyPdkOK5Jobsy48HF2h9bO/1YsSrS/8ZtoXyNGDaigTieLxVj3
vPTFhJfoCq/pZ+frGdlKzBSdYe6QDsxLLAW+BdRd97WGI89fQCeYtBJoN8MoI6NDlrppDv5jAf/D
+mcd/r/BDj+CkcAjD0KNbf1d5RCvVfkXXTDudY1sHsPhsYfM6j7MbD1i4Zs3Yf3aK+/iYdIH7zbY
HFiYsuIlmNSo8Tz71tVVNSr0xrNlMmqL/I8SY2qllFG1yjXyLItsZ5B5CsQC6Syn1ATF0atCLk/i
6AUa+VRCJck2Iqrci/RsLtrGRvtr5xwGilVssdQm+pAziU4OmTk/2C8yw7fBYkzt9/H3rDEsJYWq
OYCHmndNyqTaZo8SFBKlPKdqRQSK7T6bXTOJpOXBFmfRGY5rMSuAlpmOAT0BMW8cGuHb5cSo7aBs
2mav4MNPKhpf+reKW7EwmtBgCgoctVuNdGNKnzjruLsEyuX7EkFPZx78ydqpBxcKiKhA/FiVbrtI
dq2N4f+pQ/DfYpG1jrmudbcV7Hi9WjlKZvEzIqAdh3OmmjQ0bjzn2Un74qLdhuKPHzbnccdV5grP
NnMQv7E3DbDhanY01KnX79rGaeCLvfiIWk3MJv1Ko7X5YGDY3oK3knLdzRkNcvKGOjjES/FovT4t
tNxpGbqLOS9ZYR+fMIqYg340VAmZ0AbhjQD/YKooN1GkXeG/0qlJODS8lotFmOnKsxWPdlDsHZTF
gebH9XMwZafxbay3grcgElLGuS5q1w/XTdX/66m6/GNK8bb5K59T5BliT2UVD9K9/mQ4JdxauexW
m+GyshRH7yqEeoueRCRsff11OOjh5C7DLcMVv72urxKxZoCwFTgSUyZyu7BsxyqyQxs9B/SS4VYf
D/XqkpdhepV9mgbE6zAZ5+3FfKlM/YZPWuryqNP96zD71M0B9QX1jzQZjV5kdqz23XKEqvTL/twK
xsg7Db3iCa8pfVhJ0kEJ0jKi1oOOxpKb6cxl0or9XozMJfjSKXOyLIzIfLGQKaA1j5N7C4g6zEZ8
GZsuUS+qLxr+9aagwJue869klCAn8GEfUR1TU2RYReW590O743svarMrSa1/E+604lDMlDyRmOzC
nALzwrc5eTJtzbsl9Qe2+JgRrSR8m96tb3HK5NOb3A1SXijnFAFOK8lT5Lk1vaDWJwN4vfBi9PZy
VC+Odk9Gbjvs9q1i4zTym2lv/ZjIvhvxNbtCBHhHhcRMN//iPLNfxOaJC11jwQCPnFXoNmdDUm47
t4dP4COsUShiyx1btijWlFQleKCCRvDDjlv02IKEZ7WJTVV1e+F3Ude0VIJcyAmoISmw7r2aAEVa
tsZvj8EVToh4aAGAvSsK+DsE5z0O5Y2MvvC6Bd8kXxstANn/F4hJsMchRS7LRpVn9LQheMmoj82E
+9Lvy/U5qJJS2wJLS+5BlHjy91/uSZy4aqRWnTtbt1hCgrTgYnALD3f+q+ytrtn0SqrOjiOgqP/g
CgLvTkeuOLu9S/CAYwcqaivqkIVvxKw+BCRlkyLqQTaXLydbu1t3X/mF06LXc8F1bt/+XJxYTrgk
9MC+ik/+5jV1QLw0MOPHhSPjhMmHqrzHX4U7kYCQAk+JL/RwegxlSr9FhTY10aJWdQ8oc2bnJMJS
ES2lfRlRxc2eFZN5sVrgZJI7lWq5xgFgFel3upQf42eQoZiakufQ95NCZOuK6msdaJykC0dVADdc
4yvoX31I21XxrvARPW2ZjcWM9umO+S37AwYGktT/Supo85VxqBWsRGy/WAxOI7aMwbZgiG+Q8I1P
MIlhY7LLHOzJ0Pekzud05cIISCcr5Zk1soYwF7kCtlxmZJumv2o4zq3iHKSxrswmIDc3SjoUc/ez
UTnRFL1PeXGBpWCVCpQopJimLwNNZSXTWM1TcCb3KwK5xPG/050ynAdqd2kXEkt+TAr+4M+7EolF
nb3+z4NfsxFbfRt+1ZkPygHLLQ4Dx0T29ll4XMlYn0xK4NrnAdAQuCHj31oklGZtwj90U+tBmCTJ
2puaH1f1XnacVW197/ezbNtpjZ/O/caza3Vnk9JTV1UOypBrnIiaLndqCF2eit4rDJaLTpLp2e6B
R36xbmWkXwsXRRUxXQ/nzCan4z8eNk3jAk9kAVrGY1isCRJlkf02M+hyJMR0gPx4ssKRfoDlp3qZ
P52R2SNtqdwlMwvSPpgve2p6X8zayNn5Yk6OoRehgm09RbidlbrLrvO0AizRuNvagOrGuIYvYyGj
Pc0ToImlfMTQ76t4ZhcJUzUPEHnfbmhbxk1phai7MYG5UOjzQTu/keH4IpEkj0ulA2tI6lNcDSbT
f5RhoqRUnMaBAtX2EtG7n4rLcYvBrt8WxUwLCYK8arKG5UWXVNQm1z57Qb19cCqxspdzp9k94J2f
WjpZ8QygtjY/HuJkO3+hL/bwT1CrMQVsxH39A3g//RtgA5a5bhZhNDt/uQDsMlbHG87kiPcZtE4C
2elvqZlB7ApOgot/DPDnEg+rdO9+7e2cFPrZA+Cc9IbxyExd3iCuaaCpVny5vKOHqKIXYHwSOdgt
rukWIb/+kTN5FhVMkIv8noMFf7MyJXKwt3eWXFvWdY6ZX8FQZoLJ8U1dYffq+S7JQGiRHlgEq3oD
ozuris9EkpwLrvuOCbMwns7Eq3OgU8hvMGN9n1HkrpmHAwuUuxSTqdwJUid5Tclgo+0m+BawYx6m
w+dPMbhM8urQpZwFJELKNzsvwWPOLUPhy/ZIKbg8KBRjZkV61MxBqPQiUO6i2o67wIu/rI2pW1GY
Qy0f/eO+Etvko5TS08eVejCzmqHvFoWxpuWBBcEJKpfdUDHBg2EEgV6s3G/Lf6IJLVCHlGGMMGyt
5cwGJtdVYIfyYKFI7K2YjTzxPyrNUq1ageAYqrCy6jvkytjy6LKygnhD0f/3Tzgxsy7njKIR4OSH
6W15rH2M8X9t6N6X4RASvThEzcDq93lvb3+vUAgw8A1HtvFsXZ9e5ljuVnFzlyglQIQfiRado51q
rfL6530qjyABye3oynr0vSv7i+ZMf86C9FTOAtBXfDzjanzBlD0KAFPtba2K0oxD7Lbitg3TcZMg
8SabPK0AZZrlAoNMg3Bp6/2VM3n69qOsD6u0a9ML6iBQXbzc6beacQlCZO+pCSMQ6QOyf1cm0M7f
Vq0IpisBzONpaHN84bPlWY+1/uwRtL56Yf8mNy74Acu0EHIW3YDscKZ96Nf0/DNKWBaIGFj/X7lt
XKL68e7wlFtDlXY+1C3FT1eXm79xNv9SghASgSA/RlJJhry6GKmOa5LLXM3JUIVRjzQng0AJ3a7l
BP3NtSdbixWocdQKldfzSmWjJDAnVFq1qLFHL0KSw5o2M0kH4DC9IhnneDecE0vxG8zE8jFFgR7p
EMlWhcvDVhlEc1RHM/bzy0v3HSz0GtelY3wlE8J265v+GyyOjfARy2WdouZXpJRdOX/VErgZSl/L
EIrf4yyfGadX6/UCNGsJ2/gAAP9KBU7BaEAZlpMRTUl8H8wsg9mLOeScyvEZ4TcrN+hE2aTHp/uh
SW2xUKDKY3li8/8zTaT10jEAz+jd6IBbSrhJVj1nD3p9EHLjmHgjNxtGQ/jCIDoeiqW3zC7k5E+7
yJjsbR0mYL8q9g/ZTV9JmAbjxvtGG9dKqD5JJhilCtIHciOqE3dGz3vrFwFev89rJhTBr0fdq2wT
G28WeWhwshv+FUmTAvbYrwNbHJ+H8LMKpA7ER9YJawTt78opjPLTZSjfK038yup9qIIjzQ4qK07q
3KcQqYmVqoc6O2kO1JDaRwx02zYu8WKkmbi5GXY/43/IF4IfEEmu3/a8cahSY3ix6WWTMgyeL9L4
691beM3zi6NLVCfrH+BtT0y3ToSn7MenjevyezS0q1Q+cAoBOqTGLpDS2eQghGymPkrEsxIYHahb
TFPHTHSHN9Z6uUWXv+HgdMbZm0GKJMXUE/tRO4XJUpXtqdGgE5xOfslj4KC7Jq/5ayVW4Rx2rPuc
j7jbJRnJhERGYOKYZRWZjlgdwhAeo5diwRj23dKCA4W90kAj+C9NsIIlFlwCgpCKwHiMNIkJFdkS
+BmEa1BVW/4faJSQ2iqG5VLuJx2LIOCJ5WrQo/3LNliieqJqCwHnxTQAifwHBIWe1/5Ta8f1jz9H
X94gM+gsZjhj4SkNVtz1ULgfqMZtx+yvrkOjnW52Xfmsy7ejZuNtscjtEKUIVpFQwtdBF1kMmdTi
F0YMdvrfgOPqj4Y8dIo5EUDXHcDkLb9rXoXG+IPtZiTmw+huXnH8bkktSPmSTehhPDf+FRSYnMZC
7TzQNvFLrtrmDht6o3Xpl7tOcDZZdE5zqRA57GSHG3Aq+wuD0NK2N8dyN+mM4NNTqpRIkYG0YigR
DF6r08iIa0/NsveRmLMu/VLFeEM9Ly3/WJFpR6iBa6CkB+NSI4es+7YVSIoRgev1IjTBoitqgtEr
A9SLcA+GLQnZXIl9OPCwVTOTni1u4QQ4bzC2LPJ1ZW8w9M7NWA0TjScKfuhjtjY+tppCMy7BjWe3
pc9bbPPuf6FWxyZ2eCJl6KVdZQgxZw8Ir1vNfC2vkq+D5kjBX06WQ3px5gSCqzF+2UacrjBEwmCG
XGt9yw58RD8fRD6Ofmo611Fjk5ZLFi6pvEBhs6Eqqa1WeHguDK2XCxlqjjHggxXyr5B1vmtdG382
wJYcpvZwM3nPMYeF3gnEfRdRaLYJ/oZsqBpdSrhpfvjmZetLm3ZjB7i3dZghTtcx0/k+tJPWnWyK
bqn2XwaPjF8CYhNs0GWyF5BSZuKKu0cGuHF1RorS8JXLd/5X64L7wLmgnEyN8ve/+5NKDxI9/8sO
D3FFYzYsB3f5++NyPonx+j7uffnjpkaWWumUHj/+Su5roVC16wKK2MpYJVbqQF6mUK55JccCYUvW
ChUaVBaqmTEtyc0/GUGAxwmpNFJB2DEm4VoE8coX/tuS6MGPCzkqNUk/u6w8V418hxiyKB7UwBLr
jil/UTfJCjXgA1uDtSxwoVna3fBZ/Bnue4UYjdB1C6JfyxXNvrN8VrvOYZERaz65QIpsMzTh/yX8
pUR5jwo7ueKYd/TB/Vf18l+vIM9BbtaFrgHa24dApavpNy2VgoPLxhKmd9vDuWLpipzxY5/rI3NX
kSvbqj6AIzXhtwt1pAx/96nW2xOaI96wO3qk9yzPqtXfhSLq57kfYfBjZTgvJIgjjYSsY26fy2+m
hb+c3XKCS+9TWoRKWdDiYSHh60ddKYV4b+JxkFrpwbiquTst5BW1XaEkECeQZW6sCaBwWX9es26w
HoimUtPBOt7v4HJH17PZrE09PLKQJQIZbnku2KHPGzwammmQPdJGCaOE8hhFJaWPqD0xtcW4pHQy
XTWPSACt4m/u0sFX90iiP+6JJSKtMC9nXVHYySY/IRT39snZDohTA52X6+7ImBG0cVWjKdy5F32F
RdylFYPAj+lLObu8d/uCikxycYCtaTgDhE0lYFJ9qVTsemco34jDttnLtiGFFiHeHDpQdIUg4OE1
zX2A1yP2JvfFVqKJwpOWOutdXS0BEJPXdfkAq9NaA1bGz728FuO2RWyWTmYqlQIDB510EE/8Bm61
sjN418ncByQluZi4Qe/1PUw2WA/EGhGWbBJiZdfywHkRCqM4wO1Zovr6iTwhuVp1CrogE8PyjqBw
6zhNuIXemKv7inZFoezeO9Vp3xVC3Y86NGTEALmyiIYHLsofb9ETcRLHQ4/kOYd1/WnO/Tl9hBY9
9ZKDdOviQC3g8xDkQBmHVVZMaSdjhIdfgajWVY1/Vb5E2QTSLPDeTM+bkqpNnW5+DzcJQJWnAOVU
+5Lk2jm/ISsWUr03Jsae7aq8QLe6MkHAFExf2SZMWtfbvroS5AMWUc5yXG7i4g0I3IfK4U3N9QLQ
bQDpRlfjKfHJoKmAw0n+W5jzfUaN7BZgAhOlZMkm21JDX2qv82JvcCbHnvpZjmGmMsX+5fNXAUOD
qFwSBkpgw4xwdBhfOw5duZhDYvx1qqbbzUaxdfIC7kkpu9jwFS2QQUUeGr7Digam9v1q4c1U3glQ
mJ1/CDndqToUmyc+KaSPkKAfvLMQPCmYACo+MYz9B1ENh4vwS2GGwyyiZtXKGLxwB0nB/LP6CZd/
vQxVT8QsPikAhI9Gg1E6K3l4mxBcjvWbfvkgydyQlC/3Jf0wVRIx5sYlJKvjj3IiocbXMosrRIym
8w6ognwMprx71rZcF6wzSMZViJpscEJmobt/e5Z0WOhVWq1d51WbYV5DnmhG6fpWYf9yJXnjlkTZ
in+Abnt9wRp2aRnutDRQ/d4ubXmGUTOtOmDj572VJfz8skAJ8oxnyUseU1d/EH+v0N0Fck8dIaA5
ZRCPTjoT8VOOVLWK4joIvoNM0L1tp06kqs3a2h2vmNhcpcoCxCc6dluJLRJg/GkJ67cjA8gJIYce
OFcxGEQmEcGdUyMdGRl7W8skjccgiRKcUPh0WezK1mAi62mknhUGEQkBp8YqFv9XBLE30pGhWuF0
O4Ag/J7RCwO13PRS7Y4jO0+XM003dAQ3771a8BGJZRzOGumQiLOEtcv0897UAHF+J76j+esnj6as
wbKPOXU/An+ieb6aiX0szX5cDo+HXk7/jCVePpiF48zzH7l/DonJigk4SNqjYboMbMC25eTARNZ5
sj0Lrp1jvYLBAmW5zInxzrEMJN6yVd9cxW83ihtY+G8g6Jn/S4liBfKFvQ2w1gMxqFkEVp1z1LDx
yi3jG86iPhrGwFQXCF4yHV26WXkTa48oF4k+LjzHud9Fynur6auoA3JaiVnIbK1GjuOSg5tuzq3x
SqptSQSauz9T7UNsJoWo/bZbAGSphib+sRZzZYZ4A8ens+XU9P5QW/SEWnRc2UhPfUlkSu6JGX1T
rPTCLIisw4twZiW30uskuXIzX6aWOjSeaFTPN1YyZzm/cB+i5zFjKBFPky/YPIWRc79mRjbYCbIr
nf/7QeAqxaXfzshkNeFopCp3+HdKJrvxwDF/MbVGY2vR0gSPwAvNCfwWqn4T1TsVLdQlHmjC+uGJ
9gOnghN7uQQAjIv/X2XGG3bvIIVZ8/QHA/r+e+cta3IKGQgPQznsjTKT5hgJ3MrrzrGa5w00EZ0x
iXLZRNM6TydwMxEiY+5slZUhcqwJqGFGPl4CvdTSVX5uyOZRLBh0mMBhBQLV2/vVu16z0ysYYbkO
BkZfNNxRKyhwbdVLPJUz60xzfD8Fhlbtc5hbbv87Ykvt6DjPca5lJ6mXDH9b3UrHkh1pP3py1XzS
1C37jL/Dmccr8TlzEpKwWuit8W3OshqQUCYQZXmAW0gxXUox2hgIkJnamnzpjmZzaIB99z6h39pD
Zgt7fYFFvzUwJP7AO0gh1tsdxZs9vWb9TeAihUvLHejZt1+pILF+Dsc9qo9BUtJl4EDa0wrdaJxe
XM/AH08HUkH81ghEqbL0wer6CGtHJ7eW9FmbxMeVEBxU3okD+ScdjF3Mort9WkKqqNRvcwRwf283
Sg+8skwRiXgVJxcOHZlsi8LTfx8VPTh96mi3/TM8r/M0uwrgNLNEvBkQrgqjBQsLVuNawMyzIW16
RoP4r0gD2/qhxza5ovrqOj+UL5dOY+5lwokkzSUe7PlNKbepI/G+wtNe7VLySsE0wCsmqsD5DS7u
SzRPPODbvq5uChoruyDwoYHUP6J4NTujU+8715lXS520+G+9MCP9NOSajjXTsd3IP43u4RagR1qT
+nRNuq3/eHByuTTJJaKRz8KoeIQY6c8j9k3TVizLOPjHo2k41svM2HJIGNWZgNPzVKmEITNvzrZR
S3hIkX5jgt1NcRsXFl0gbIYZrc2XTevpPeK0sd3D4RHTq2lCll8bnSvNHsda4gR3WDOeUwK1Wdvn
kskfCCnv1BoiINTvXqilvm2AzbSUfYr62Q0DGnVRLiM5ocliXuxabUtEV/fmKy1oLNMfwxGKvyGK
hPgkOzjijfTrepdpfdbxghBUYKOK6zd2CdHDfOnD6Evv0AcFzGH4ceqyqWV4aJVmDCukn0hhwNkt
pOw9XC4tAxbYBHzr7XYDQY2ZMIFN64fj2NmDzQyEl/4xkRMcH4tplEbNRIFpu8cQRko68TgmqJHC
ZkL3e2MqJxQQWa6iwe/KvHPN8mzZECzVa11OhgKnMujbEoPymwJ//7IP4bC3jiinJR3khjgilM7p
4tcehGSttxiP9wTjkH9PMunG7/1VH8OXf2CQouGvNwQt/QQCTSBtH3a+rts6FpSeHR3vs3thbvJF
DaE5T0ZIWFTh+XIMlHV7886JnvOm9S6PjNWu5CHTjzyW4Xn9W0WqzUNI0povhVD/V5ydvQvUGXav
NNkOgWsL3eT7YfYY0G+E1nyOM36po4ipPUhfS0FypMxzqDbPM+hlQiky760VWEitJ1Rjl4j+7yih
l5qsC+d9EQXD+K6/JyqmQ9YvSaMwYHSCwFqteVpW0tGx9qn3tgKHLhY1IMCnBZrN7vgdu1FZomKX
48nL+cktbA98uMLAFUiuOmXyLmoE5rYjAQIcgZbi09DYs7Tg1xIG4rH9YeGuTyx3KgmHPpIPCvFe
F+n2tMCs8r3UEr1Tw+Pn1lflDOFop+O26nrimMds+IxF07NaVt72u1dzlrPfarbMA0cMx0Tb+V+0
L6uNvoaRhhuGY5eeb425SALqTQfxYZTuyZRg/9IstTHmPOWZR8MBK0x/DQyOK5wZ0SBMOx+MORF4
TyxbjrlsHUdff6ZLwI+zMa0yv7YDU8hLWGtp2gUMUVdUJC51dLFyHmRIjhl6TsVAIY8NktmWKGVG
KOzJ7s72lHx+3m9Mt95j4Ons3XvaQFSOINxAqcEB+7JJAP4uzbkED4lMb0bpaYNI+UcP5rw4X2Yj
sggg1E2g17lNaACWzG89849/H0Y0Cc8CalOzLkdLanJexGP87rVZ/+M1BDIBREWrDvPOcuM71Pnf
hrkPtzQM+lO0fSNLowfsLNsZ0YTWwxXoZAZiOra2ndbYRZn3UL5KF2uCWaJYKVq8oERz2T65dt6E
s3sIlrxJTMbrPzuScnSao41sTeaAC7VzBJ45qdDa+NnYUkUaz3zZPQkdfFSkySFcap+NlntBtO8A
TAjkj6tLP6yM0xiuUylaEUDP0CS5ceBjP9HjCvKugoRk6QTasXymOqt5m1WkcuG+5eXDtnkOqhQB
9t8Uh6k3TZKNwuSK/ZF0AKxJqcmKZRnz9ff04HBoenuPvZsv5p/6rQRFjADUDOT9OkA+k7xJFAxA
DZguCnPGaeCsBK7GK9uKwuPYJy8SGZf278HyIR3Aq16TdTNH9wgLwXDkF2MlHxq2d63HOIBzQggT
LGa++XQ5iam4KgmORP43PBoFd8pLOa775g2hl34SlX2Dotv08XvmYHWGbYD3ALARtK2psGzxw4Ba
WWXLaJFvvqI+VrgQZkWH5083IUsG7NgRoZGg4Wbcq0K7g1MUI46INhHxEZCHJaYdWx3YRzou3+9a
vXTEP56Vfo4Aqh+U5eXQbfmuN555xcWnkdy8R+TbffuZF45Kn2CftgBKqOle/SeSHSnCWeyGPQSH
ePWHmZare0tUUOYLuJuxHQ1uj2Yss7MIvgHwlLxu18g7ESdTODBMriB8bAChg0KbQtUem0KkfRXs
IMVFIXqKn7I/+9Vnj98Op9T3wRQEv1D6wXpEhaazlmHtX62rM6J87Q2aWSkg3ytCfs34mnqeqvc0
Os64mw2M3clDbTJbmgUqmacvm2s7i0HNJJc8Ic5KS8s2G3A7D1zxBBZ00Im2a+EYYPMq3rrPMAaH
DDIBEfHZ+E51lUXaYjVP87HbHIq4ga38phXvqKw0isI3fa5Ky7JM0uAvl+5ZhK214OkGb1WY9PGj
7XlpSEqdMzEA2EjCtmUiZC9376U9J4S9E0gwjRU5VRSHZsdpab9FjP8OvhZyZ+swky9TbkLjrIXX
Pdzw4B7FMsopmmxc8zE6TbLatogtcC6yZZECmZpguifSq5Litxs+LJSGGj9iw4zoHWsVa0j0ycGV
QO202C5QQAa5TgzRN6YHVs+U7Zj15gEBH0Vr1HwdFAx4ZgNKD3UDFpTojSPUHUbMgAub9brmaIsE
4naYkpCelPLhOfQmUfvwvNkHvH6Nt/9iYXJ3TEdbYozcinpK6/eZl5eLSfYRFOfafwDaHiDi9VYZ
K9/UY/uzVVrg8Y9TlwINmG3rQ2fCgd2ReWdzTTh9wA5ofBsLptAiHE7XcMPRHQug64Wm/KYavqYq
C1DqtERVss5IeEdf5/MLnpRxNOfVHH2rPU8gMd8+rgwhnNQEHcSoke39YN+2aq0BC8GF3jv470iS
oJlrp01fL4FCgYzx2nvsx83MqFA1GFqdJ76Q5p7GYn/XyonPqItB7GjCR4lGsrBPYH5hJM/LDJzB
p1FUyOddbBswFRdnwzb6Oo6WZ8jNcryRIC3jrktlhD7Z+UnTBOuj2F3LlOfte5Tpdl/7ic9zGcH+
qBBZDJDTAbiweK73AmhSGtytnJJGEaYmXzjee6QST4HJxSf/d47/Ilsx55a7PmAxtmo3smcD8Iab
6jZut8atKJpln7v/0xdha+lObyXQk0jIodwi3sTwzNX1iVLnogGgtIHPlnJGBj8qp7Dz8GIcRZeY
H9pf8TyHzE792u+hy9wZBn4OsVTZnjN1l6Du31xm7HIO+lJSPYGQH+A10qvcnF+iQ2SYF6437AQI
54Ls7gTSiJAkCCJE5N3L9JUCuHQbMdK4F4P63O8r4rDGFDdCNfEeHlrKl534l8dPuCAGX2mXB1DA
5ZJtoJ2GZ1G8dW4XbtuIU7u827zgGcSXrPCjm2QJFW8pZ4OCf9h+1dFSrkislaqBRdNj/BaFnefx
oHRT77vKDZ7qgQPQgvKNfnBK/T1YuWYZbuEA7Xlc6GkO8sQnN/mBfCN0qhSce6ZOug6IHvXMAeP6
sQJXMEN4NNiT35RggRP1VoRPWPwwpnMQVCu/Rreg75CzWMIz2Ryx1/ef4R0vXAD3Id6baoan+GOd
xHoV2AGxv4nZe/5WvQxsx5JhKlS5zjpHoXdKzEu+HSiXsanNC1s4SAeMKh110oEAgAni3rzCT8pn
XjrJlZXlRcCbdcPnHq5RlZpqf0L4kBNZFF3MyUpL1mUU3Sguv8Ob4YR/QGJLs61AbGhOwmzCcNuC
bTX2Yg0waVfuSrxgPnX0SSDoyCn46+ZefoQC/frHzLm7iU32C3DFanDvv72TOjIA6fw9BYfcqu8I
Hjy0rzqpSL80BS7jULeZX17Ok3pjvGIPHt4MfDq6OAFPqxH1gnbVezaw8q9niwKN7R3jJo5+oZCo
FflxY+Mfee5PTAaNbCJF5UW8BPKGoHsB2Y+tpt94yJsnuP2rNiLRl98QOBcdfH5gUUiuvXogYzQy
mbeifi9pumAKMLw9yYuqWFgrW7NOlIVyaSyW6ITnmitd0MBOH08hNUQ4VPpXpGWicZ5oPTEtqQKi
VAlsD4pIEH5bqzUvd6tSNRmrR+5IMGWP5r7CdpM3oHaZ+FolGOZi4335n6iTeHwNsQKH/yYmmO2j
pXY4ztF6dQYVgnSNvJF01wxxNEcV8FR08cKKt+SK1LQttozPQV2zBurUuSfLHKNelcrf4pLPZdFb
w3K5A4hjO6Vs5/dbeTyN39Wtw7ZmpEYkFDhKQsy5fb9ff4AkgkUku0PT/NPKMi5sKBidtW93dP6d
RqlcNRv9fGXStTLvj0uuXJLGu5gqorC8b0l11OKW+8FZXJ50oA1mFewvjp7jC7/eh1IIJgchOAqN
DKNcqldICYMhH/VXxsw83vCUqVfVtX4nIT0rvJvCj2QvuUBjVkmCZrWBX3aJdJBnSKiZZe4pg+bE
nJPY47cwgPaYpL9NTV+/HGDSpf+qo/0jxE3VJT2xjWQl6ZecjIMtL/pZdn+ZzjVcMpk3jpL6B71z
ljzjFf0xhdYtoO/8QpON/krdkT8RW3OU+EUYcltmG455oviNT/1pDiJP+/JysWwh1wbfu1Qn6Hzc
kow9dvAhrVJowe7jblHff0kNUZYp4VBGYXD+jgcjFb0s7gwVNXxb9JmICHQuBxYdFv4GiUSLRRmc
rBCCiFZzqN2ylymSaFCPykyFqJ7r0NQGGBqiSHo7iepV6zNINMUXGSSy0oLXFx/u1rBhOuhRWaFV
yDzAmisPrgh5eDnNmKAq8hD/yXXZRpj6dMSNBcGy+pYt1gnKK2Wg+CvE8eE3qiEQd8g2KiHqbjes
tNhTQXY1AA07H+XoeTi+F705af4P8weLkQaFzVNxT94ncx/4+KdvJKuWebxKEXi6aOpksW7aO2aC
MlkVAnvrF89TkX8IjAqS+oTVRRzGGK0n/lBQ4Ve+t050AzZ63KbID/Do9n+jUnhQNrrj4PgU5nVX
jr5sbM6pkfiDHLPoD7G1u/n7/WapNGxxlUQsGvB/FdmGpYsrAC4Hy+DoekQbxMtPviSK8VNPDl48
Ri1BF5d+kIflonbVWhTOHUV4jukInR3TkkSYRW/a8xQVfpo4IP8hfTO7gAjC7hlwFA6kG+VlSxDk
zw0hQbY6hgIIMv7dMyApnhKlnTzBt2FJpv2Z5Sb91Rnqk455qfreL8+q+1QrvBdE4ZSSnCQs2MNA
dptBxzX3/B2gcEnlOzJ79hTSXuZny2CHLs98UiavmzRxEQsSzIWqaKk7CmKLCE5xHat6lD7hGy2q
dnpIvRmfHv3mY1HfIyQEf+DeGd9v9+hBZ5r5Z/7hFYTyH8Zl767ySP6Rrfh4vqUwSLpb3SVmN+/j
rwmiTJbzDexAscKtscJOr5qaCeVhFY/hZBMZv9Fsg9gUL+CKWVrBiJWYjrxS0uK+tF3UlXMKC/KY
Z3dyzcC4lXmIQh/Vd1EUD30Ca1xb/ppJHYMUQeAD3VkSGXjFO0wSL5UIIka8lh5sLsRoaubpvNsa
64yfXmr+c5Lh4t1nSHnvrcofgAybCeMel5vQaHnFtFtEWKE8bV5HVWi2MLQNJxYM1Vmsk5Dvi53+
vDDtkN2NzlJPEEhPRpIEt9rJdQVVY7yV2GqQrhjKd7eUbDNXG1FaMTtqfJ67pu9NNq35yAgCFRj+
pPng7V/ffN9B7r49VWpZcN/WUV1BobVSQD8k6/Ut4xZMBKNu5J7bzHD1idVcHJAV3t5h49B8f6dt
eR4AzmT+MKbsQLdpx3yvlasXKffYM3Zv3rqFC+eb1tWP0h+aZohse11KhpCayIMH4+3pcGORdzpF
KwCTPfzHODzWZ05WGFAyn20EZxt/v7rHmGVJYk30bAfH1tBXY60uVqNmUwkqp7rW8zmfjuzHEBqF
kQNM2hKej8NcSVHBn1h3pymKFOT9n63gXOwZXfcBbE3YzM1Mo20Uz9R2m6gcY4WWgPsE7EX/bU2W
2XnrJIXvPae/1kjtg2Ffyi2GCQPjqKIAkhFFySXelROfuzqJDRGNo+/yTeUTi5dKToYFc7o8WEfF
GAjkvg0qqG7ioVIISx8tHc1eIGSkwL3otJ7aFf0fbcxCwzgj9X/mjEAzKU+h77pPAAt0p4CwgFwT
0QV5bPlmfpa6TNJ6lG8UgwE+I7an/0KTt99fKuo1BRo3sWR7Y+rGmg+fzYajzBvM/IqvKLHydEOi
p5sk/hHvvrB8QME89MuEy+qJTC9pQw5cU1x+Phz3xkNBZoeRvGrxPWV+oNsaBJlOOHdsjiHV2VlI
7mLdGoMl802vgSby/Wp53wc+Inb+Amn/ffxI54xae12sbfNMlSSuCvemwqs2etz4ZvNLcXNsj9HK
2eXLXQwhQsJBPbgsEgtwFVMG9NL8h2eGcb8Td9k6nmiG0m7wEkhJDvdNAHHfKn1KioGTFJwpHEuX
rQEcAY98P2KeEUxRF1jsXuhXb4kNqK/oIu1Bt8Tv8bkzdmJmIRIu9BTfmsjDGhS/j/jr7UAIc5OD
tTRmN6Hx0ku5IGE3Iw8N421zYereFl2SSKjUq/8oxYDQXefj6q0IfSgoIFLRDOuPgnimyUqiEm8S
BjAPUF5j7fKk0VZtGVXevjnfZNXJlvzJ/f/umwbhRm00T0QG1mYbWkcA+u2KMolmEUqVFdHh9AFj
J6y9vd4OIpciiqpcWuSe6S/AGdlelWBI6B0KsUBM5rOFpqkkSkN0OB6z5udfkQ5UwX+X1T7/RSDU
AZ3WtycocB+p40GPwBILG7DrUjm5IU9JblXn6JjIoqT0fgfjwvNfLS618s+dwFroRzodClPv7ilS
T5MfBckkGDnb9EON/HWxh/FR/kA3PtCEiecom2ZOTxOIMk02FrCeiDhtksOKMiWH23QF9SofguXL
Wn+B3+cHgEjxWB7atFgttvvPt9uUYJy9TWvlAL7e2/0ApsoGJkWo5ORWfADDBYWNiFtxoquSv4H0
fI+tDwAmSv5WkUJdeOjlUbFjRy4Qrpw1NO8TJQfyxYqWRScYcNyka06yJKA0/Lp9S0yQhrlGJZJB
c/cpuWyFY+sFY58jC3h5VWDZyDLIF72oMvWdxtgT1P56QbQ1zFB1bZ4IBgRqZ7h40dOVdC5L4dE9
lFaF8UiJkximkIQpN9zqFQPEls/tsKtKkkIR5wR3tIETzPHQ4G4bMu/rg1hTTmYQ3OqOFbHeaD1g
RMPEfnSbtQvLFG/bRsZ/zzTVzyud+NXYurjzkZJxb/GWhZZ6KvgMbErbo6ZnvXsyaAZnrKK8KoFz
1RwiXy22rtPRSCtYpy+69sC2JEhgPcE6jKvnInyl2Ohu6nH8RXMGLSMDxt0LfNgjZTfIWsZ9IZbf
JICUZgPjh/PACjQZmijncDQIFyJroUyehM7gOFtcyvVmZobADIquo9j0umjFbUOWVoIzyCdXWGdz
6c+TzPwu/r4/TiF9OREdR36x8TwBoaX2iT7xGqEdpKeCDY66baaYcZ/X0prTeImOduhyx4L110um
A5DUcyjh3U0GpQb5+7K6TetFWK02jxWHi7XCB50jMEc4tMgBT/L+6vEa0mDDMmZYEdR2pI/EJncA
XoG8W2pT9jNMa3VYou+4LwWCIWWJa3+gDLBvVtM4xeSousJ7r5hADBbwmlh4Oi+KhTW2zNOtoV7L
8J/+/mj0WHzgsABw1/nzaeYmRLPrnWExa+8h96QkovvBFLrnAQF75Ut4uXhP3z1fc4ZSSgCY6gPr
wpSO6usJniX9d9tAoZzQ2gVnvqiOJJFD/T+ElyC2Qh6LrtOonyK8YF+Fs680WHrIpwA5jSxZdoJ+
1LCaAoRzgOBTk93I7ZG9ne5+8Zt0F9eoRlcWbvVdU8hJ/Ap5gGK+q9h5MvzkAl9+MjDPPLlJDLV7
14mxyQB5Aec4c8RGCDvNH+kXY0Wn+fjqFTLfTYfHoWB1xi0Yx4pXBZ8HGi/P1LAnbuQXPRYMiHPO
ypFoLgJX+nGSv9Rse25+yw4Rg0EzlggUPVsYNJhCzm//OiL8x2cNAnHGWsrOlSVn6pylEp85hKaG
IpSsvsyuW+M8w5UJXcPodGbxXGd3P49sHXiCOXYrAihoM2KSWtVF/oRqglHDPJNsWI/n57Lns0Vf
jqM2cB4Y9qh3fCcsodkitG1h3yC953j38uWD0HX6HpfAnWfScXjeu6iDm58zWLRaO7Iq18ei+0uh
g8FbeaDo/bxZn2sTjuLuVuSuOIa5aRfOJ7X4tKr2DbtNTDOjZnlvRm2MPbJ2FMEcJWy7auPtTT7V
q9k923Zrq48c5Mq+CrQH1OCWr64grTJ1nt1Tj73Su5Omtu01tsYKrfY5bmE3w2ncRo/akb3Db8s7
oO0YO6Ysf4rQT+c+1Y0oeTjr5B+DoxyA48iGkYbUIqn17txkOyVAHzpC/Y43LSqEGOALC15dMnva
n6TvIbSf1erDfBWjQpHb0bL/VyIF9rcIcwcZ/3nNQbqkGX9ofwu+J+oiR/LFDzQ0qpF7CViegLsy
PG4zN0JH0qCFjTQrhe0gv154I+YmXfjhJqrEP3u6pwekjfY3hUqG1+RpJ80NveZvwNRML/sq7DX7
ECvUstjUWquYHCk6Lq19KmqTGy0vxW+Hh41cHUhqsbAsm3mqW9dxaV48lJUqW2GhTQbKNi3ss73Q
G0P1i9MGqd0Bd/zu6NBQY5HBMtupjMULmZhkrUv+gdEDelTiRhjmT65ZPXjjuIHL7baUsxESZLjf
9pERxvPexB3NvVUu5Zj7MFryvg9+nWdEJcpDapqy6TC16uCCLzsX629p+ZPSd6iVkMM3Duf6fBcm
hzB9eSkkBh36Ev2kZPCNA3fVa2EUlN8h1mFyvHcpYy7dMNztYhiZuiKPswrnJM7XRDJtr3l6Ocx8
eCh1puMp9fQsMU4tiY5w8MxZBdCrnDmuYhJ7KzKIxhZv9zRHtZFDXiLqDYJW10QGLNAoLKLghrAd
M6NVqhPOO+trCflTzxA/VEqGLCmImECbFtXSH6Qw2APQwg2CB3qydL1RUs52PbnzdVvsqZKpvKI3
l/hG42QQaS747gfKYwZiVuBHMGrW64H0pQh/IcYxuVZaYwuDOrwY3kUoMcEGdvHQue6bWoU08NED
TRhULSu7iHB8hcikDzcz4+GJQplytO/aWPJwy8WjjDTBeSzJHqzGa0AjXTz0yd1ld2Q9m2j1GrKx
PlUbwzEXAmm8Ogmp06Y4kvmQOZDRGH5kcXPPigcc5xECaRjaqzmXQegebobMkU2nn12RdyMELF4Q
AmCkGMFQZ4OajOZbg8QIbdopU2m5fJlVJ8XT6cQd89xPtPVXGDZfXekcBYDTitK+X6SPmqeQ/aaM
ehGV5szvyxDKr0Ku2thzDmxz4h4DykeT+gJdxuAoT3BQLI/uijoGueP+mRRfOSYUJU73RBN7kSIz
G37+aJECdMtiTqj/9WC5uAEHIT3VKncrCFjIG3hBvpMOAeNuS6VYd/Ui4geTxdtvz00x5W+8RVqz
oKvdUYWjDzw2YgSn0ox3XeiLiWX2R/p1AIN85D8rE4bER7wg+43YfeZx4+guGMVBZIGfXjYD2N+f
X5SgVbsrk1WWCZGg5Pi3N4zsmiQmNLktrj7nUenwy/MeqCcFpGS4FqfxSdVXB2urJa/ZpJPpTExW
ysQdf+aP0uEFyYJmZ5jE77F02Ef4vjGlHRjed7KISe5bYosbusCAutSd+pqqPm04kOCYiF2CGtqP
33p4tmQLFpssISM8xWMOz6S6gYXlhW6rcJO8Bn9OlH5TPo69UQDx/xAO4wOOvmdFX/cey0Ym2vN/
9Bk5UWBtm+o79Rq5K65sC5RNC3iK1ML6ijBrTiTwW18+z3x11VFmhMMFio7cPPQntqs2h+AggDtq
aC247HoWXtFHCkrWKb3GtbH2/bI5WR+wdIabvXPcHT9gE24oAQR1Op0IRGsc87f+xWWsAwuZ8S2p
GCpseALNdRM3YUr+l0xowCxMZR4Fjvs9oZWCessY1mVW81/HHPVgBQwmm1kvnSR4P79vrgQgsPcZ
xi2iEU1iMpWJ1xIIT1SJdSBPka3AxkJFuE7v850qe1sGMDINbBgcKij5Nn6kW/Gx3ARxfMKtEoow
vuWEFFvm9BbUF14U3g6sl1Tu0V19XudBOaCV+lKkmaScOPaR58yG8B4niDNUIa0nOnkDy25HQHr8
q8hKjo0t1Lj3DN4OZRTOhQSyz60gnLR8Bi6b/+6H0DkaZvtgrHo11H+QeWdcLC1xW3cZTvZ81wKB
QDsRgazVmBEsVXv5AbhjuvF96oXgxxtmDKCP2XALR6KrtUhIeLnZSU4q4kmnQ+ri3XIYflL+rhOx
vbJthtsm1lOjFZg2mKnw7ZhTIHBEv8Vlxh+giL0ffAvGDKsFBTUpWVQTlV+HSOT+v9SUiM2QEs58
E20LI158vSwYiQgy4JcHCjJR0QuCf6VpkDWUo9vf9/4lFGaZoxVZSBR0USVhOGoL/CWWsEZYVV+A
XwdPe5tY+DZNEXXJDvK6spXPh8/bC/zePHkCIwDLHBA4MFtY5OVOJgaAjfpS4ifvWW2qjNMxOl4N
U7tp4Dh2uK21pIBASGj0ggWRV4jXXwVQElnq/u+J/94r+D+vKwYTZf0X8iMDigVoTPbebYHZHILq
v+6QZXf6fRfzLF2CMl16r1pXyOBXsrVBTHh8/mPdJPaRNiIEXRt5ezGTBB4YVjTlXREQ4a54stMi
VSTAoqEfzpBvUQ9I8jm3L5PBpeQ0Oln8TQsbUIEAEcUA6zRDp6NTOv96+5ZgFQplMhLe37z4mbmc
E7x27pVUCGAvWnHcSloWJs7Ah5f+wFgk/P9/tN4sJvWDhm3vnPsqE7IUYBtBk/dZlHS2s6Wj+JMB
EIQ8yvKjqMe3vULcAP/xLMR1gR3cJMPcwS7qXlik+GMkvbId6X0Q/0TAScvhh1PpQizyHkL+qvAT
yBe2WXu/tSaBHteNCURCCMp/z+i2VfadJpX+beUsLRuoup9t6uu9p2lNJ/LwqPSDki2cj5w7q3aJ
lLAuRB6NyjEU4PMbhsEyGZdHJMGx81x7x94OzqwpPPtsd4KscYB4ucMFeQ+4KgNojgiMYFcDlXkj
lkWPI4HciLV80N64gdxIhDGPxNQIyU2ZOevzUUsty2d84msNsTDswV6wiY85NObYJcFrU/UkKaLQ
0ty8dGJjIiD1ixYHYRe9oXOY6ZYOSht9wON8s36leP9uxgcCq337uoR/R3+t4tAP5fV/iiW77+Uo
2GH3iTYX90vaIOGgr1soNinrpjhAvsYbbLQlYJJM2+0MEsjA5KTUn8ItQvcMUgXXju7MXVISyk0h
4UfFtiUpGeSK0utR7tJtWnt9iOurYTz0LmlUbmLdZPo7JBbjO/WMMKPHdtnAAfi3Mmel4DNY65JG
jFIofFz+I2V7rsTWUNZoxEkM9mBs2Su2c1zhEpt+ZKXOydxcVJUuqeQFSnQnBDvftpjuNlyuNepB
ynZ64Y6+bWsh1NRnhpCWXRpJ93B2mOa0yLp+LLFJUwlseUQ+69WFvovaB8nQ7qZX9aU9ZCTyvY4r
DHPzgaNIUHe5i22NsN5A+sgeP1OoiqPxNEkuNvkBhpKMbCAGu8RvZIiCQOGdLAS4kbbBY4qXYBQA
rT4oxdK2Ol0qK1xLuhrcqfKgTkUGnU3MCkDKCWCS2hd5GmwTWq93P5Vg4cLwPgwzf2/S6XB0h42y
+mJnCuyfF1QFiaMVfivwlzj2ctlKDmjgTuTWkqqoan8j1pwJwep7pMEuYnvTBdsRPA1mK6Ng0oLe
f5KiHX/FRO+bWQ6/E1mC2pHFmfeZL3VkduiPCXPCBPvMoamx/FBKCXmFu+evlm/r0USMtNdF8zsv
aN97CkDrZhopYi9cqLTG0E8SwuxWBeti+ecSB0fy0qSjyXhzpYVAF8Mh3fP3AUT1oxbRK1Tv4EDH
enOFZGTbYWu3g4NyXik36P0wW67igDaINGsLY6kepK0mZm1J+Rp8gO0xnuI2v/ppJiQO8rksoJci
0MUSCqy9pcXmH3m6eudLdx4vAOYvFCMnhnH8ShuPI6hK3R547QQs9d3LnCXoToD7z23alVEZsYpV
CoCYCwS2Cl1hxobv1HLuo5cKgxG0aSaOz6O9PJIJPHML/rHDlvRqzilkZIt/yoaIalTDSTljl5I7
ku+dKjcPEHnLgUC/aTInoZuCyQq+jnLP4bekv80Fp1nD89AspI5KPnBRyDrza7ta0T/JirJP4lEo
Mm3avKIGGaM6RmSDDTTcSysWGpY032S/uCw42RMjektAfcyvg2kwHzzyqvNLOWiLe6NuBfJaA7dc
95244s+s6w7mvnOxGwzw6NQyvX/g7ZKBf/YUGg7TnDIPMGtmgZjBJC62ZXGD3Z87wqhQvYaF9/Me
Tz8VGJSxflcz+iE9b4x9FivDM2MxlZGy/4gtXTdqV5RAaTrBeSF3d78V54hoELOT0E6u3QnB5Wvi
rd6hfrdNpeRHXQsZB3uszChGRWVc3HiUDz9M4bIVhKWAU/wdTgUBT7bcmAY3e24TRU14QlNG8jd5
sri9UsV6ET/v4uUYRgn1VGSLYn++BOx4B51+6Qk9I14yHYV5YqxvNWFn5k0JW57aIQDFACy0xMS4
7W6wqrMcedqRGf+LoE8kYjWi9uYy4PX0gVhdZVYgBVMlsgU6zwAaPBn5COWsYogm2sEP6et9x8Hb
yqbUHgHPvHY+TXrDa7CHPKYRh3mlv3Y4Gbs3AeNeL1JM5X2Ty75qplBNP/4c7bRUGxOdvQ4md7xg
hapmrlfzLNMLEipKeXOz3k92SHyVuQB9kul+SiSV7Fe2UpMcob++FXo1rNYVV9rHTkqI5Rm5TrnS
J1UqX2BBzifnKsemul9x3pi/9pH8+r5ONYigfg3iVf9NpAt/iqIu+cLv2ZxiappneBqCZCCXm87q
TGAqy/+ecedfkhncCCdna9rWHwlGtQjH5RrCi2pgW0vDzFkA7+2A8ZhnBa/WvKuntlp6Xe62qtXQ
+rJ6IEF4BxtHdsNPSXwcHWuYGYsTRB79VY46y7EYylTfitRgIDZM2DRjU6mqMxOoCS566dg3xCi/
EHDyYlhlpcdVUd8O/hUAjY+oqM+BMdnU+LCscveI5I5EbMEFqf3WEGfXnXdpFQrdADuQ/oDUr5e7
aSq9wA21enx28VourH4idsBrC4FRl1uo2xp9YUZZrFvD4iwtF5+SeJ6BA1crg1xox6gIa9IX7ByC
EzdaIO188DwCHNHyvQyiPUP5Gp3zP/UqtPSieatlJ/ptBMVZiU1Q/lCRR7EESeXvLy46v9NFPsS6
VQP1HP+vDt+VjwAWDhmMhuHgvo4opXEcfLAVgl8NLHwBdmVADFG1mQVhREt7OFlcbd1766w3tQaE
jSGneNFj+4TABnj6djDue/yJMZvvpFsU75lAY81G4j2r53ZEEp0rfZ9T+uymEaEnjU7HBKmM0nTr
JPMKJBdoz7aAhIEYjt1Y8ezNesZmneNax2MaeZW30tZhc+OHDpFIAr2ygQD0Uu2A2K85KRECzg7+
l01jzsZPR9IrDtYUOQvINcNtC9gv+wP/tyg3iQVaT7kkf7DphDEBOcWxSw0Skhyh4kEz2CqAk4ri
wCwld4ENOgEGMgonh3Lszqa40Ow8Oa4Gc20lJoNqV3DxBmifXRj3FHNKvMLYQmqEm8bAB4xXkMNI
OLq2ZNNjC/4UlkfM18djS01VnxJp7an3Ahf1Rqi2id3HmXVVgMjeI0buh7YCciGbo47ZvWj2UUO+
c9RYH5bx4eK1JdeiJB+p4bfBeJMFl4g6q7k3UotzuuaD7Osl3KRSrpgFO66n/hBmn/pUI0E4Xrts
4a+D8M28grqUsXth/zzezPfULE5ztKLUU/XpFHsPrheaKD4amZKZlTkgb+2F56EsikyuTjnQ3waa
wT57r0CvdYbHg13s93gWCYjNCYjR4CDhrNnZkZapfJO/c0X7gRhVaYB4DdGFAU9kScJt4U0HJR0E
3094zq1fbsraXtNMd5ROUwOZlOt7GtcCGWOx/+ZOPgQ+GinKo5bwvo45weDNNpX0v9qFgXulyAr9
mTHINHkXh44bno3klJxKJ+Y0V6j+VthtjOvFtLhPjtL6mBygWDcjgrJaGsANr/y5qGexRUaXXaeB
yv+A4NOZTyXRbkCEmk87GXSywwxWMd9unJ0qgC3NpcfU0bbeLNlrCumVpU5FCwGPSTe1x4CIO5cq
Pu24KW6JbRUaHXpiTK8VRYnIQpADsOCfSEuHFMO7NxXIPMO8Dp3KU6X1NRrkYQf6uinSZpWaoWol
uyZ8t1HuoMs+UEKw7y7QqQ6hsHuZwJxjSK/l4qq5hKWiPVGi+Y7xL9Z/IK/GkvbSrl6NiS6fk88Q
0UGD78clkxdka/mVsMR0suxM0ttT9yzIvTB2qKb6YY6x3MESXembYYypARujqGb7C7bAR27ZBDL8
v3nxzwOnDypHepKDmJ664RCKRHz/VduLkAp7aiaGRG7/C1fKcGsJgn7yougb05GlY4SxCXgFVQd9
jnXIrPoFTn103MO/lu90cGL4VxTRE4+5veI14U1DkCC7C++fZYo2leAqfAfzaLmoi+w/37cz6TKr
hFty6F6YcuS8OF9/XRutIAuckNKxCh3ymMV7pql3WvkkT40QFTAvpA3tQL5o34wBRd8BBX2IXB/f
8TTnSSQ+L5sLGkpsRWlxPJzQk6iSSUqZy4k0bK5IIgxnPyWYyWHSyLCZb8i2RMNDjaMfiTcA4xGf
U+FzCnkE3Qcv/vmr14888L6r8lwNrQ0jIYJP5Fu1t4SHtY948FR2lMx12CJeiXmcNkPhJ/nti5M8
mYVnniVipoQ6eTQMPPMJdDDHTNiJ8ybQEXo3axqX2B8Mt7etrWmJUK9+un8/qR21oSnKp267bob0
KVZ0NUk9iFJKnk8psYp5Y7IYX/F2RwmkC/x8jor22vycb4WTn53nsRTBEWJbIy7Yd3zR0qixrK2Z
niXR+Qj0tfhLDEX23P2asw65Q7YcQw6cUa+rWL2WAv1XjrS3jXc+XZ2Vn54/1Kdj2KyBOnVhW+s1
2Wq5cRtBN+mK0S2X3saAgFa+I6FvRSfb12xEjITeklgjgnblzGNzcMGyLkCy+8E7KSjnCS5904Of
oL6UL8PCLtz3NG1x+Haj2Mi+ou3s0F9G37mBWaarLU1z23n/YuYyMhCM616KZb+WVc/EN+LxO9lW
n9xru5TmiojIc9j4GO/L8NdBo6zmFsQ+YQcpOumj3K3PEBQtbjYqNa2PkvShTxUGWjfN1+L57CLm
hZCFCP2YQZxsHsVJXyhnY+V0/GNLxTwOANRnEdnI7mmFg2jMRhL8BEwIVKNiPOMft26S9Uc6jHV9
MSJExwOg+pAbeNRG5KT9nxtJrdW1oKwSHYlvUVIBzUvELOBiLc9gzYVkjwAEI79vy105llBh034h
2ORIZBoZcm/27ZRgGmIlqubPpenGNF124cCAXb0XQUtGItsOQuVSep9MPCSpWf2dGz4Jtlvct8Ip
g61A0lsD0Fj9Uqr51PtYXN9fg0DJyckoc27EdBNZx6yqWI3hlu5c4srpUsSrR/x3cU5T9G1C4d/x
UdC7w+9KS7xlIQuKmTUfbOfWh2UYywwT7HMTtwHMSSbWoKBDUa3qp60yFphe/PEtjMzu72kAluXJ
ODC395dwyKa17Gg0AEYllRvA9FANmb65EEu044KLrTD9RoxNioIaGwBtx0M/UdFJj0ZrMeC7IOrH
uZwaOsQIOhDPh0+67/5XaUMOZ/OIPFlng37eba0Gl6he69bCIhH0Pub99/2gfb6MQjqP70wtEz4P
ECxKuHWbqJIjUomsBsRQXjOdxm+t/pGz0kgmJ19VvbDvNatB1Vc+xgypago3Um1yXiQRVJnLoEi4
ycZCqGUmFO05LjB5Kyj4YDYlvXwHpeDRfJM40tcsQUuRcW4Acr489AXvNdnlDuCVR1EvbMMjUp4S
JGXKOXkih9Ndcke4zWoIFzw4WUXkxz8zvWZ1EZHETCVGV/4qD71TmiaRQJOTUdC+KNIIUzrQ4XRo
MOjpq5s65GYL39w76DjR8M3MNEO8XCGjAfzT/bP+ebjbGb/woPzX21cVTFsXG3WbMM67L2onRBks
7c9uhwsLDX6NnySyoFdfhKmabbekmT/8zotSSHKNDHDdMS+aWLuSqmtrU1EKAzoQe2FpNlpVOmmp
L7mgRVbuuj0sw56AxrqHnQR4oV7fMnPjUmzYpR6/nG38V9nNCHnzpn7EAg0XQYC/oJGvGFyYjaUy
W48wgsJyQlf7OecduXxYVs2kSzBKi23/QqHAhjAj8TInOakXLJYsjYMelDGUN3kA9dOqhHSnKg+Z
/O7dqt8xZJL+aQr7KZ1beEYGFOkj2O2hblaldOqXtYWKnG2T2T/kSjN130F16CzTFFZBYfeuM2kp
AiKd1WR0eWJHADGvnFZDBznuBS2RJBnW4/DqROlvOh8N5ZqvamqYqqAeQrBN3rCiBYliOdnBczKb
bncMBb+NSgXY6zGH/bHh1WnBZpQ0M0/DaMK3Gw84vtYf10mABRrrWuVQHen09qYbAB7tSVIFj47+
zej9o59BMNuFH9g6oAYYB1l1V/a93TscxcM8IO+HIKOcnnQ2uUfbgh9aHr+p8GK7Y2zGNNL7p8J2
6ULln9yRZ9CzGsZHAOxuEDQEYYZf6w0NQeVjvDgU5MajpjA16ksNIS9YpACF0i0v0zQScEsEsyDj
1srlDbd1oob+1MsOjJV1OhK469BBfxPNr2dqegV+ltsA8zoD1AKr/J8SU56tJ7ciGzY9eP7kO75N
iYQ/QCqqKKXh7amc/6jDa5cwizCeWFRvw8qkBEVNMxioSF4fhLHDotz7dOxf1Jt6VuWsNM0cXjd/
ac5PFtbR7ppd0w8ugR5ZxhjtJAO4PbteoyjE6E6lYv3VpCPufhsy+rjJPyv4Fy5BJUwcH3DAoXxR
nKSf661G4p9GVDaES/zu2t8tp1nEXwQkg+h8YFZwm32FZ9jhHEnh5zsozZqy0mriDTCf/sG4M2zg
0pi1M9BNXPoAiuzFQjCBCq0UunB9QGBzaKPHOyOmuFUhuu++l7yWbep9aWimcx5vstYsEjTuIY1k
75C7TIyca8igqXWTH+Z0YpY+skfdCiQPudKcGt275LPNWLIye5go56pnMNol/jmmoCH2meOWm2RQ
KdpJjVaRhepqnTpVgWCBsqRmO9GgDsrQFH9WRad5c5eLfJTi40JigN/kPLzKCIVEnzYiQDkoSTrG
ntYJBJc+Zq97jypKeyJHSWgRDKSFzXItITI+Z1GHevHMkhJVACXgtmqZ/MC5oOvQuqAMEcAOGOjW
4c8NkSMuJz5VQttsPWoyGlsXOWIcD1NOPb+5XcgtVGQbGp3VTSHCapu/txtS9Kj0KZh57aRxevQG
7ZpvoLs9MYSEfRWtXC/OnuWhYq0TFaph95MRHKMUTDJWHrf+t+7kUWRazmkUG/llrILgiWfXS2kD
wXA54mtbD2jMxXVTsCe89Hnhe8mxmqbBJHGt7KZ/iMFVsfYktBse+yiZApEqsqhjgVQRMVwy4v9A
D/XD0Xp+92g2OaDio3VtJeMZamdQ7PC4dfII2A3HGteBXJa2S3LSSAlAj3hqhr1XdKhwN06vfVBw
sAfK+5tSkZq0KbZV9KPzuZhYPG52rk4SmjVdR837uvYm45iHFMgBOwikc2zAVn9fDdznbDlzyFpG
vp4Hheblr6reVeN64MW6E8xRFvGFpcZiXyUbuks8+woOzWrmYvEIeFxAR6dA7l59MdRGXMR5xFe7
RDqyypHG1nkVZnW48RD8DS6a3qPGptrNkAF5/1cnaJjfMqjxQQh2v446KUuRoSt6sLRFAZmefVUd
YFymVhTGHV31IhQo7ZZWNrPtmjsB0z21gczHcWVIOXkLnplh9ZpXlls2trjcQXIbJc8TahxR3PQi
7KJMhaxBilnQkTMXfeTz5WT2BDnPfFWKd1sjib5/KYN6AnQwB7JJUYlkh+Cm3VBxhzyKAzYVMUyH
5taSedH2gnFAAu8cNFOD7Z+1pJyQ1PrpzXJfCozVJ12qj3H6VPLOqT/1Ta2DGmmRLRet/pX8mK+a
rjgqSYVTiGdfuRGOqDKY/iNy7Cs8ktwi4HgcF7X92TqjjuiXCv6xsSCwWjWa+Q9zdM4dK6YTcYFL
2do/Ywe/XY6+PfoiYn73m+VssA3Ej7yfcg+Y9tmxsgPVB/+DlrbtnxhcFqAHxACUT4Rid4LJGEdP
vN0wLbwVZIuMIydnCaRMcbRylbfw/k1GqpSkWHwqCCbIG0jNzdyhRcVZMDS3MozI8Xuf7xawMMuQ
BVLvd1btR1b7gvQav4DcLeYFaqaA0o7ahL634WOiNeOQAYs9qZXPgZGsTIvW2fRy4lat34ojWrs8
xunnsV45FE9adDKcTCufTYiGk9ufUNkHahW6FXEXp2KK2IkLukK5JRg5OmYs6yEez8Ix/cIwhBaN
A2s1x4k/EhWwVid//Sn1hu7dUEMFt6X82+o7o3Yi8KVcAscEWduiIKuUk4YDOYv5aRneP8m3ImLf
ry6rob1gSSePKnVJVyhUWGfvGZXTlueFI01BlBKtimkD0bt/kIB9ZXdWV6XxyU415VUscV4Hhtd3
Xz/SvyEcA4K3m0DYyjAPT7D5eLTIWdV2d5MX/L1VpciVE/VIPx7MlrBNIVEOh/ibOXvChOKDDP3Z
1wAexID9rwxSnkg3RoKPS7VmrYiShBoUuPiYJVoAKqzfv+i6928WTomDaQ3enmQExL6FnkTqMMn3
SRUVZge10rQdAYdbhGp2ALp3Gt5vupoUe3t67Ke0OpNBz0VYrxAky+Usquyd+pnetSKWlZaAZmKo
cxq8MB+6LEegiJ90+FSEWuuKoc4lo+u3cf8TZchaM4TCZbtOnpkfg8axE/dN+eFfan6XFBe8d96B
CxNIuBLQMTBWG/re4NL2c2ExVTFDlhcLK4E6NyoPkoRcB0WzVjBY/BitVrm6i4+yKSRZqKbQAVaX
SQKH3ifI4e83467g4iwlJvTb+QsJJoGSvEwyDKSVVio/3EV63dNJHCPU8AVXq9vgL+lDw/bAPKI/
LtwCcYdGQjcZX0AXF+91GSSUwmZUtHZfnv7BrXko9S76aJVuLeSIDCzhjlNGNqT2vPcXY0NUtPIN
vMKYfDijO45eRbQ5NaSq49s0VokKph3ctSMNDNzID2rftZUk2PeDruHtn+m/DR9ZMs4TLGPrsg4h
j9mQDUXoE6IGplIMS2XM7bFqxMcJZIBuzJhAqXUo0PAIqQ3910UaByZicw5kohyR4nFCtgHYmEi/
8oL3mZV5ldeiaioqNgJ96qBgrlgxnRG68gQytfUeNqxeiShdchrqLgjg9hAdBTcpRIAOODShAXIN
6mDqL0RSjPH3IVAlvThg/SqaD1zxKquW3J0CzfVbDi64g00XbkYN9FSahuh+upBg8HSnd4GZjzSp
A5ev0tFgqwVTkgeHkSqXlS4W7785coRTU2bAsWyG0SFOqpJaLQJS0ZVOFtv2ZJBuqs021Ao4eTtA
iAg3uWfbETGg2s5VP/VYJZnJ1tVty+jJfd9G8rDm460vINIZQ6MFv6TqfEMY/hUXBigCYyFDUAGL
HJlMvwJCnMfVksy0gbNUXUoaNbZSGVsVZS3/B0wJXjhpkdnWuaJeKyms+796+t9Bsv2hwf6EwtNE
zyZ1OXl0YSh/T5elSIXOG+K7xnudJ0is9ND9ca/YqqeqKmTJhdqi6zdkZC+lkv7IlL3UqrMSTexQ
9wNGmKhCIrEbyzA/gnxd4t4+SGva/5A8JM6qaZ/VTNMDDFn3zFsC+tOtEqxgn5l+I7K//WW7miiA
/FqqEM73v3kNNuRXjTeEytI5G4Pp3fICHX7JfMAgUW1ML2hQX0hK6xu5L4QIlDjl0l9QZjzum/9Y
sM73FVWTm+3Ip5K3MEdYNhVt2DcVaxSuHXdYUCaavx4rzd5HX7kiguBmKxfjoUGPhC477A8J4d8x
cCLE3a+MtWXGeaHB1YHyzkKtpZI/7UCm800UAjiQeVE76t6VOl7RRf6QRDvbIv/zodMOpbKPHGEs
xDoWL4rxWN4814j2SeUzxWkqoW0qUhLWgityJ9dZc68z/w7Vg2RHv0PVEJmPqvH5p9xWXBbQBQLD
ueQ9UevMeaDS8Y2oUZ6KV+wDG54s+yHSFtvZnJ915XyZR7PnXcSVZKpHo+PERCsCq5l/2P9hZMPk
qQKpO7LqzP6GnSRqnlnaVn5YoWMiW+MrXeG8UJBgW+Ru9LnSxId0NMlSCFyDGZHrDR1mshJtcDqx
2Gcz2gGO2iiy1jV0O76zKkJt82/1FpTKOQmgMUOu+tRH/2RFWYQL5EYaL7XPQqx8/Yg1rpyWO+g3
GX9m6gv6oFhf7Bb0j4fVEm6hGtDtiaUnnuUiEayKyG7JrKcqgkNmzEqSkPIwsUI6EZY341kLJmbO
JWJ4bn8+Oap319jdiXhZ4b1wP5YdqMQz0/bsrdHaUt554Kx+t8PQlw7OTZRiu9GLFNJVUaYmOpT4
gBYW9fwn0y6YAUe7BnhTStFZHYff3C0megwn8RvaUbGn8M+CEDgty2I2fzTgf9SVKOx9TnfKTepA
/zLtEmWjsHEcI/NzLHzGpPoognJr2IIgv9asV3Gvlpp0igRi/Xv21SYXkLnZFQJ8BYOYVq+GlBRz
biC0WxsoclFPtR0cPTQAQeFiJ3YD9a4h1XSFhNtgbW+tZ4UCqN9a2cvXm3g6CTd++p66V2FUvIVd
MfRi9oaeng6Kv3CBmU/NqiUEWv3HqbJqhMDqe8k6Ph7aK1fXp5bTd4CwKg5Q8vJqUBkxPVqIh0A0
0jpA4VoPRhOovgd2tQbJK5brt2sCRmFsYecrEJM4h72ps4Hc/XhilTo3fOqeBZVA+SU3ykOd/myZ
VYwt/ckes8XD0Utj23KVENDoUhac5irAMFNyz4MP/5JByWJ4tnUpUGV+Z1lT2maBYANPYQ5QL+it
Mv+xC4wEg0j9v3Fc+A+gG9q2Cnmwbfud7XAxD616Qe3uBTnTO2FAcFwIffTyP3PjmtFxlHNT6Pph
VdsYtVX3qZd7Qkn1o2szN+L2hxTa/9Itn60dGfWZu5JsEpo6WcHHoESWwKWXYB5Mfy6Fl3NGovla
VEQoaH+9TRjZtpaps8kWE7mDxu2NCBM1rYOuxQibQJgc904xygVolDkzOcRrEIk5a9+Tw29QE4mW
RMf9whi9fsnzc7yMaMnI2HAKqxcoJCLLeyzw/GOhKlhN0iJLHeqGAojE24Nmw4kOWycQ0z/SDxBn
YNaZhnKfkhDS0UBDEkoisMdsdGvnF/305APcWSa+1j9pC68yqlDCqHARlbud96NXHYE/6ils1BaF
3l8aDRh2awSORBWk8Ogk91DPxyVL6KxuMvFSchX1HtbrzCexUGKRJwC2vZtezVGqSHK6b0+Nj5c0
7GWqx4eyDx4TdxgeJcw6w77xvdKlCQa+Db3mryf4sG27dZJRmNhe66PI0V8yZ/r+/wRShUBImCez
RNKCv+hmN1pNuz3MluVzLwpKrsKAtOc3F0JCQjNQgJvEixsIJKah8WbNFdae4u3+44p2cPAAKUwM
uqg+owY717Zr7+J/SW4QA9Ay3FwR3RRIvdEJ1V4aSr9C6VoaokHu01Ktq2nqACszE2w5/NZ1i8Kf
ZNW/8LvczaHnO6zv0HDHBNb84Vn3aGXZPTV/brMHKert7gvk1m9qTqB4qR97AhyKi+7a37AEQj1J
EVY0+5LEf63LVzGihSYGRx1FmhJI7r9wKyD7Adp741/8GMFc94nbasU6C/yJMX2heIy0cg0J4l6S
lodGamQZ5RTnRizhF3GfV/2LzGgVvlxPp7oKC0a+eQ009llRTFYo/qPck1KU8MgyDboZJ1GE7SI5
oJkkqvGGV1rBrTWgbJp+Aq4T8spbgpKYJQ4OjlKkicEVeOLRr/BUskPHN1J6osvQ8mv/pQtjE2kE
Cmmq8nS7ihVQsxx5JnON+cqrisa1YzWAP3wlaNS8hOs8l9h43TF44O192xNEN9YCzlT5rug0i1Av
6R2K6Pd1TKtJ84m3a6KFXo+tMD+BnHTueoMDqmfB2zskv0P7enpHP96zL+5Rm77a/LqcFwmb0jJI
wQLx0/8GxQVFOWWAAScMcGxNuym3456tKQxTzNI6nAQbK6eeImbw8h4ZWWPxjXHJszaP79pP755W
gIazk0cjwjH9kQVhN7N9+vl5ZoOsT768jYa7zC642UTjxmZXzaJDH7yuIeb8cNGv9B9sBv2VYwwT
jCeicIz8RZHGqKTRYI/H+9Q6rABABDT6JxmPMp1N0K+7oDcSgyXdZytpoze3Eaxw8MTR4EluMgJY
KqbGz6yQK+w62gyo/1TfUe8CGGXJSzg1rPC9NLA3+HIcTQwUUvQGRVS/jDmvz4XklUlOGp3o0r2G
heSq78L9SuLhLlA/4PDYBKUgrfR1HBcJTy2IsbaIrIh2J0KuPj6jXHTxAg+ZmaXBQKdFgceEuQn8
tN2tdAzp/VdMHQa0O77MlckwdhPP4OdnpxSRhP+m2GKt4DJmReMjwX7Kmj/fR31+KADbLJ2ywKlz
vT1rFATK3V18tRELArVG0YJ/Qz9m+uVUB/9CyNdrDXbeaYK+DdHCoD5MI7k2QMTBNYNM6WRV2yup
N39lPriTsECmRcnEqTH9GZqkJvq6/Q6AZyQr3I0/l1fR2AE5N2nC1+IzOVO+mmg6NG1vLkqZn3ug
Wc4URIzPJ2dwQf3NdGSUdNwcDVvLZMTt7fA1rJ2GyQU6jB7yqgyBNSHxCku9SsM84td6bNAeB3Dg
JSYXO91mO2AQTYUmvFX8LYFtSPNHYL9CjEBeiYvLgxRogHz8P3NOL+C1kTDaMwiZPkJ0OCBcuFU1
WUCoWmdJ+W5hBDOOKb3jStrnLfKXJjRnWiO95qLsRrcPivXO2bAgA+cAOtwYFrPsEVuUaMScad0G
KBSAb03pNKqs6FDAXrW5GbdnapPVcupcJN42a52wTHW8bmm78T8CPPCx79wo/+Gx5oPQ6O3rGm5Y
sxPtk4K7lT9Xd5Ju+1j+kdG8cp8nkTqaGB0v+HZcux1XfxHlWmlIvlqIPLJfP5i2+H6fD9cuOpnI
OtlegitNu8s6vo0lVMfyoi0jP+hZCoKYMOJvFN3wrdLDRl/UKNYmkobu334eqiz7MjX4QIWCGpH5
rQL3zw+i4eOLTBoeP6y8ejf3oknpdr1gtI4FNZPIWiBnRn+N6Rn+/csZ9fvb9MYUFZ4JTa8j5Z+2
yiIo7bCje3DJIhPWVaydtw0BQ7GPsszOUOXovrl09qznYQWlIgjaV0DihmbG1JCt2mp8pvGlRrMr
hjOshCe6iMDfCU7TzAp1pxFbu5avKj0KOKW3dyWggLQSRpc8WDCRDyHH/ZRw1tfzqRQ5YpXvXIwd
zpZQytYVQvWevUoT0DgHebPwVUwt8u0v4+8ysyLeJUVvoL56d0fL7emvSQqE8RWr+sT/jm++vVxk
sOe5R6pSXtj5oTDqPBKjyoeDXqSPTsZQd/SyILCp3BhjHZcAYCBTjtOuSxChBhbO1fMwuy8reu1q
7C7S15xc1bhtvRJ30AtlfXSe2jZWijRwcYm40sv0nAEbbldW4rH5/NHjpyCfUXbr6z7jThdqLAjZ
03MWmKTsHT4w+7OPg5dkbPr+my59dwNAC+H9VElafou3OVp783ZUTkcjXHs8KgbeG1PjCS2bxHi7
Bj1TurqMEOyELdeY4M/K+p8nLTr+/0ekw0xLH2oo/iED+qxqTpdF5TEKhAWII+YPJripzPyyYcEe
F3GkScABjvGLb++LySRQhRpxnHgz96YgLd4h2XR9dhfOb5rdOjlcuh5n1APMnqS4nG99VrgJL3sk
MvmWGDlZQ6DQ+eljrs2fx0AOQghGL6lBOwZNrU7DDl92I6B35pAQyPSOzMWa1Bu/yc+sW6gOz9ke
leq3TWun1dzGiIFwvM2BEGrA8T+Ly+7yi94S1SNLvzZkBXnqkLg3o/A4PF75rTlSX7UknNEtmq1f
5Ws4VrKmbQUBoA+lWlSTCZ0kMx8UK9p3VFqSrHv1cECufL/my9vsXYyDdSpnGkK7/u+4A3bhvHYz
CkpyuJ9NeXagm/atyR818ik1lQbPnYqK2QJmxmyEemzwbBSodz+dwOZw9L+XGiFX151G1rT0qPEO
cVbU5BkGkgfA0jMhOE0PSZHiA3byRcSMZ+KSw0veG7f4NUHLd0fn4NZQXXvkPUFKL7AKV8Q5b/sW
PadDm24NIKbrB38xayVDDFCyvs26UWhmQPo0e+8+LvYcM3gO7kMPJX8RiJVdirmFJ929ElmlLmC9
mmHC9ssDVwDxoss3tbD9rYHV2+WcD0JcxmIICntcS/Ihdj105kyrqZ8whLuMGdRmdNKW+s6K7eky
YIE9/BIijqov0vcBqA7J+v3au+/Ak6Y7EmkXoIks+02ASkzqNlQ7URWCuoj0ra0TFOrtQF0+IuHw
lT+VKka5P6tfaw9hwzlJ6xeapztSBoJ3qSk3aJBTArpda4IEBfvonliKEuAQOcijC2WN3BpkMASn
jMG2Gzka1T/ztGgcgXzRjt2gSEypl4MBKFGY5J5EZY0WSkm4z56CtTJ1TMaN4Wcwbl1HXPqI1JTU
+UuGChHkmn5CxSmmyQxeszk+XlCZIukNViI9pDUx76JsY4YVl3tTIwSmUPit5duARk8BRJUCu9Ll
LsWiEJ8CiHkzAVFypt1eLofQeijFmjyLo21o88sFoOayAQVzBBKNbbBF7jYdPN4984puqoNk03Ys
oMC0HbEl7chgsbsZ2yfzhZPWMCYxsXcpiloYXCqQXORcaJHnp474H6v+7IVE9sEx19LjPAxJos4U
r2ov3lopw7UM2v/yAF2yGJFQ2ZXATwbDQ+yJHETXe9hJ6UuPXFjp3TSAci5EePBjt+klesnEspig
CU4LCZHSUraf1S+FxnH/v4fHgwAe//fUKwn6LPLcV8+b+2hviZCETrzLlIuSvYBI0wrXXnfm9IhK
rtd05gUxcMnIJtm6PMnv2OM6jlOiPb1Vhz3lWawtOR40K/aDzkI1VmXVxDhL8rbbia0ldIBw0eHy
60PiKsgvGj5pVjyb/cXk4R8VU6wgQ1Qqr+E/it6HXAazJyOs9Z5keYodIGxFSZEl9+DNF8gKNRq1
mx6q3hHa96tbE4FvxDU+MrbzDeYwxLY4mupzjsNM54e4ncBXwn+0/sHSno5twQOi5dOwHa/vLwLJ
qPIaVl2fzDrYq/Cxv0IdzXC0Vo/cfzeKHXtVJYP50R/IWwiqBGhpv/OZ6EsMefT+bJGGAYiu5M+e
P0GVUKNXDV+4Ku+V7V3hRXlEpJNVEVpKyrD1JbLeCg3zJEcIF5a/6bAy0wLTSHHJWAbDxWosE+T1
8HN2+Ay/cV+yZDNsNUkOj2rWq2xs0cxqt/NAC9bTFDedR8jYRkWzLvBt6CBIHIm7C+G+8Ke2j7LY
E5gR4oN+WrNLmPB0fiU0+Fy0sd3BNgtEtjfbjD/0+rBSH7nKbFgwF5K2vNk9xQ9X6kc5Gk2yStzx
bnxexA4SIrUgiW4Yw0EkbF/wKgCWhkS3Hh3m76ZcNxHQLjJ7GxzV/3wnYZF2tB55P1zksIDmkSoR
Q4Rl/UjzBG/Ofe1hb04Ok6qXWNcP5zJHU83uEW+3UmYTklm20ZxUOQ7ONYCaTa32XASXrlBY52lu
hRaf1xdqK4TL7Tb0Rm73ltaPwIvr/DTQNF8of9eKNA0AyjFflWoMWpfd50ZEUKtVQ3i70YsiaIp3
xiYVqJY9bcLdea9Ycfg95vpZOLrf8zgbxOa2mDBGwDdJxIbRpjkiXIPU+JP2S3R4Wnaal4uf8krN
RwAPza3SCH6UK4VjuqdM+L91gGtSrDp9TJ0j0x89XEuLBS7/n6XC28xdeGI3g7VyaD5yuzr9OgKy
cVW7Tm8G4EgEA84iaAusyMDZB5zcoi+7ZsZET8iWVFb0FoQSYtXb43KBoxiVGHAq7J2jC7Snnsq1
7veKeySa3woOr77ggfpc4ZXZTJFYnUB2Lo+FWQ1pLz88pSeGOL2jsCINFsB3D2PIYfSR4YwMn0Fs
ikR0RNegwETjJMNRi2GWlPwstitnajqkQS2/xC2oQB36gFnLXC/zptRQeLiVLrs4DqPcgKBT32uZ
lsPX+68Rg6CVRiuW2vhtlYp0A/aj2gWa/uClVhGX755CbMhoaOJfeWZZu8pAVOC5gDuAGWX5o/B9
Z26cvRjmd9o8CDM770z0KHM5y7oaeMm+cWF8YpwaF/aP9C8CuKDRhwqhkj3NRfqshZ5ZFgTSA4k9
lcy1f42kco+Bb00PWRmK3vuF7DkZGHGCbRLTQPZiaMH10WV2pfEhCPaRzdgtEgJVuGPSnMvJpxnt
iFOHvCgsVaA2mmvB2Bmd/Kl8OxcjWaCJCAsWbyFS/lzztqSx4kwU/EAFkJTOPYRrKiYLh3m/KYqC
U3SERQJVjmphtoAUi0wPwaZ8GmJkE6ERWQgmU1/SpZLl5xAz5p8YnppSoct+np1XIFdTmm50zZx0
0m7Cxw4HtBgE0gfDhXccitLgFjBCbGxMYu1ipUCitLrI+fEe3EWMUyrttYcoiFTFCP/ivxzR9NnK
X7Dccu2CLJg4iqDL0EJwTRS1B6fT8U16Ena3819H468t8jtMOi9hHukpTB1Yyea8Y/EtoK0m2uhU
dbu0Gm84IMt1WN/Ook72u9bf2XpZ15hbfPod2cOz3yb3m79WWiET4f05Y8Y9KAixAQudK7BsBJa3
cODtrOqE06pk0AkzHe8ARU+dcLG6A3REglin7vymhak+0q3MPKOcTutgYGiemtvXEa6i3SQPh8ov
+NNVaZLG1rIrT2ATwr512E0mAmQ1IdCBBX2RhgUoB4ObKfmoheMRZ3IFhY8uP5EPtfoU5q48K/a2
yTRcgD1v+quM+YBGCCsIR4ibg/pSAa09VQMi5wLj14letx1njMjxIUD+Ml4KDYubwB2JatGlWhKs
+2cpB/4ZYOfbSeRoew3ENB/3ef0KZ9jRy4jbCrradViUU7j7a7cMCcJPX5GCgx0tPiSyjzrqrZza
NH1YbxYfJoGA8ieleKKrvgEW6I0KqECq/WdjP80uVsziSUO8dBdnSJcI/yXF5Aj5euB3UclHV+gs
uiQbZz4/4ewCRpBd1eAD5TVvs+snKu978Kci1zC1i/kh3Z7tQUXTEaB0A0k13PV9iK1pSy70BWm8
xHplvTrKb/r4TywDg0uN4/L9XXNrZiLzVHR/SsfYHinGOLIsI0zJAxGwyeTmZVoa9S568S2pSwrv
DMH4xucJqtNyGEXbmowfvVWQ3fp4IncXlYOEGeU7DTdDjHxUvOpID5T8AGIbuMBZdIZrhaTa9LC5
hMzd4Xhl6AeDoVQswYtOBFWbQ6vSzixDimRdQAdqWJ3z/UQ2zVZfW36IOOYDBXTQlA8VSzdr6AKl
xZR/9BzxQEn93Icg/1AIdMLszY/o/6U0JMsPOtAgFK1InEkkfop0BLuZThqag26prsv+wOTDVmSJ
iHxsnbkkmUlyTH8dLbQwAyLd4YmnM2I35batCVDmACyVq5Xtgakanu7mR/xsnObtdcFbzfFDAHBC
BEGxgcI0JniVpfO81NqoZlaYHjBkC5Rg/v2ayaKCSmiKASWwyRqkevguJyBS8pkw2B9XSHgNJIqS
1UFShqz/5zXTuZONWLaY+QO49oIpCsW01+ZNbBaPlVb1bH3K+xHwCYJAorRvO9GYdbVhWFbFr/1i
Js/gqhieAd1OchWysL93oxMYl/ip/CellJJ69OwY1shH08Lcf1koEDI7EHz1NsaUNMFo4AVzPq3B
beKCWu3l917zPLhlWZYPuQutafkH0zcHqIo5v3NC03kS90mnMEeEF5YnAuK2RNGV+BjAPVbdTjzo
RHeFLZKCj/O1spHNHWw22EYF0nNUgIM9E1eez2JiKsfCxPxAV18MPjCJE/s4ygcvt8Dpo00c6U2e
f+olVepTLSnGKnC7Cc+hdg/R0G/Q65ttKOZldiB8AP4JzBGzX1mxJxXJVWtFWvUvnl3UM+ciKeK9
U9V9Uiauz//F+gBRXOtuUKbpJB70VwKYtuYLXA78UBxzB0tadWOUOs1HZWnegVYygrQAbUD3tGbW
MpEi4yLiKsExqjkcBs3B4cmq4oZZUdojFWeCcKOs1zDJvAJoPEwzMTPjZgAt4PzAvoIIVPqiYIlr
k2fBxsBlE2mYXZyKtcPVpt2x1AvccIJTusDC8/4a9/mVIeB+K+7xuuUdvJq72M2Bjn576/MzJdW8
ikwIPUIZEIvm5T7bS7qajFV11rKbBLTCKhvhCCYQM9RlXOyanQtlXMW8wxIvTDIpPtV/fXJMS03D
DJLljiqaoxMEiBBg7rBZHI3Ie7d+I48Q06vemQAbei180dcPkT7rQejb7OnDJ3Hh3y14R9lzsjqz
XTQYrbjO3eiKeFNqpBqhq5Che1dvMQCvipDPzsU3nF61hY75cPRWrjpGwHkrRr00gYJJo1afKRJy
3DFTfNaUSWegfijcNZO5LJEtupojXMj94QgzW95PDC2HgtFRa3f8k+ySay6pvz2GI5QMJsbK58Sa
UkDf0aOCGbySGKLqYxK+bnddth8Zcb5pzroyH55U+NidDSW1idiQh5qp1laBB2cLikGG+OVZ1Ewg
ELWv3DzlwmqbW7j+8+xVFXSi1sdR3Tiq0zF7HMXsuJgxM+ZsJicgF/rxz/P/g6aADRMzXfibDAlU
/yDqjMMHtS5MM62aHhA5IuvCiQwrKm6tmkotXP0ecUiG73qSWOwOEyYDIKC48zbJVY3IA6bpRTus
EgdIJr1G2P5dMdo66sdJxLzdaVVBy0OaqNqb9oQzm9rj/635YVcUL+cXDk1Rp7UIrvImAr2tg6jV
gXyydALYHYdUFe3wM1h8C2w+UoIe4AsWy/rNmYmtBj4EsGDdt01sqHy4V5CJ0OjnqZyBgmA2e1ig
MlISHWvGuVIezV0veRynaZGjyDxOhKXVpGwpo26sWKoPlEwJ3Tet2F9fVjzB1ZFFAUgEbWotMcVD
5gTgmKetsVcU/q4C5AA1XyMTQMFzSuZq4bCKyV1JnbhbSDkpTpaBRLaJXiid/h7+QzYCFFP27UPz
GRHR5BfeAMlsl6MYfUIzCYMz/PXl8mumxBVg0twtLEvwH5mBHoAWiklzZcdqCEnW/pleTziv3pd0
gKQ28rygFCHgnt3HRl5UKM3JDlxtuS89W5ZX15KjL3DD807D4LDFm5nZWMmyg0EQe2Xt3OrObucC
ljg5C0+nanNvJoKbFewOl8tnj3sBY/qpg08gYUR3AInt78hLb8kunBe0AInYGbCi8gE5tmo13cYX
KhwiS7ed8iVGbYX0pNLoqaNnVASiTejaptjWVil9ed4PsOvPuJSKs43J8W1xXytL4mGq3yugVdr7
xpyAiD0I5rzrp7clZa0li1qvLggPxR8pSLHK98YVOjd+mA8jtf4oaVyfv5b6wLHDFpx1fPFSs1u+
VIZ7jXRfESs3FKPaeyUXywMINA3lMZvsyn1K+jyQrSIZPZ+1ArGBN4Z7zGqvkOxALETM2hIoUs6f
ie4EcTrPKMj1VMrHL7GP2lotJRFDI7v/Uy9HG16xfC1+VcugyFEH0K3PwP0aNXtFesTHyvIlVByV
dB5wyEEZA3K+C7lt7HUOAMvdCCdc0nkB5+n+GAVsxFMuURyzPkn8GLs6F1q+N8HmRMICe937cy8S
RMuN0JTqvmtQgvD3N+9Y4kVOdmIps2/hd33kZYCxYtI4Kwr+oKo78eSE3s9MCJkLFi7Wwg1N48BI
iruPfeDrTAq09N0yaV8xWQvpkai9RiM3IyPbGM2GhA+R/HSL15+pu45aDrCBIRnCF3iltCRHQolc
pzXIApM78iEGYrYK1VY9fv+Q/B5bx6gFT9z0etz2ZZAIsmyCpmdvVjVeyGPZVIn38GWqZjLqZ+CW
VuZo7NMD9vFC4It8xCIAG9U472isdQbxlrFY2u9MZDlOzzHJchF3wXpfsZ4RwnQF7Z0GFoV9iYC3
ubVe56ImNj6mBXu2S+Uwtmwtc+dgcwoyuJnHziy7S5nAER6xMrjt+YH9x0CbEhI2Us/6/cp0Zf1L
f/IWCHfGfkJsnAyBz5AjSMa6TteaaoxNq6BRlfS8YOuG492Fefy24gew2JDFf7jXMH+7fJUvjJru
VeLh6XY0GEkMvYg9AxOYCJ1GDF2RkJrutL9NIr/sD85UihlAh/dpEBmw8LzbW6pPjyalwz7jh29N
ZfwJV0Jc1kagLPg5+Wn7bxkPU+3QBIxc/x2GfBi4OeijH2AyjoJGCQEobrBy1PCep1tSjPc+gEEI
qf0dHhK8GptgAOgKJKvYObe6ISS4WX7AlWOHx5HMSAJre+gXUv+iEsKPKU2PkCGgC7uaqaPVRRyC
RZ/sod1USyfqAN8PEV+o9hwlXREV1UZSZue2/TzxnJ1LOI25mX1JRRNDgJ6z2HCWThobF8OxOQaC
rMWZDz6xKQq6DR7uR/EjD1PjIC3Rl0I8gTxFYxU6RRnZghmUWDwRdGxy682Sek4U+5CfdNSLK0zu
EWiu5nPk7bYMlYUBuBhE034rX+DBjbiNsGZSOhvWN8R2bTr/53OGRWQVo0/3FbmzCbtRNgF6aF8m
nSA0cWr7F2WsPTvZ40RegTlmEHPlVp5Zn6w/yEIXKRTFA78jg+nUVLZa+4Kra0TOtEugvx6rMzAc
KfZxIaQM9jVMb7vu3+oaWM4JSOJcqJDlGRIBG7C5qgsaMFzuCyf8LCYfGaTl4rUvBAWKgUtzL9+p
+jWLTNmtUP2no1F4uKjJzDFas1mYXrDKJsuiXHmii8JGKnMUt/rGZ/oObH74PaUbBfsHpt0+smfk
pJRlaqjfMknIajMOShUO9ChpWvbmIQczHFLU1qeSjkEW7zka4nzJhBd3/eTNPdccMOdJfur4Qj+5
PLnm079Ug2GNbep8h2u6mOcLYoDwfF79s9faWhK9sba+vd1AJhacij2y6KelWhHAjOtH7Tm96HFh
2xkfrpJoG049lo8yXyjjFJdcSGnq7x45VM/6eetAJ3lgLNmmoJ77RvflTV1bOKerl/ZwO3qfochV
eB6HRIMw1TUvuwMCokzbQK0GE6ij95Hy0oCbamDmpWZc6BRqWmEwBFKD2VSON3TexYiMh1CTyBkp
fS1Jh1BDTcUEOKN4OpPGas5mk3wO1QW3yU0gGhqYG3NP0DdwUgMxg+yZTOXG3PjB7O/7EZeJemh7
K2ZSMHLh+kQRw+BrK5uGZ4x9bb9S5PD6b1TedNgQbdZRwnHj5efxybUZqsDr8wQ/Yc+XhHhxtygG
JZTIv+OoURt3owF/WvghJVG2VyRx8ICzsbvJhNt9XYrqtaDAoLPw23eqKZd+L6wUIKy2XDdLY09A
w5Tiuij+feFNCZFi21ZSmphuOQqTfjR6sUei/kO7Zuxl3xBIB2u6QwmLNbe3iLjc/tQRQgixbjVC
T4SjAaaEwI46YS+Rxjob+Wa269AOBHkQCTOXHc2ssgmrH0FHDvsU06ucWL+iS8cKhAaqqc+vJm/d
nX3z1irSCQkl786NJ3dQbt79C3vOqoqHZIV30nxPlbuCtTR231N7fN3S1HF9K3SoKwBsrtdWj/08
2WVSgG1usBYWt4ZkAq72ayKlgEOPebKbU7tT83i+qE9Y5QxhT3RN9Wd2VpVHNfHI1FvPjlmFRFew
9DHm4FHj8iOvVzcZf71+k3VLwGmEJLbFT6pTpnBeVWQtkC1gKDfPazEu70sCdx7yFtNdtJTkpwVI
2EBImVzYr4bN3hh6Qg9+vgpy3FoYOU6/jnv53T8sKfezSzeGdvuRKqTXiCzW2xqgibMm7dAHQIzS
W51ygY/XRs6c2TI9TPpqyRcIBQbTYIxLfFZ4CWhv3SNxihJO/Dtv3ipGfLCpLO+kCfjr2IV/01OR
5j6dGX6m2nOZ2y2Skc1reOjFAnF4hDr1SwazuTwLY4a8jFMHuZQ3k33GqzKAOqLWWzHmB79Kbwx/
CQU1ShDJTzQFUXX6kFLXL2rqFRRLITEevVPRp2LzwLji7sLyvX89x61S09jfp2/ws3fdGzjNroza
oJxOw7Ng5SSziRtt23QxkzLb4I/pWyRWQ6R//h7FBeVHXexB8XTIkMxwyFhFbbJJO/ZYcY3BrGUw
lFjnMM+hEidaU5tD+Jf+iGNjDyfF4VRRMcladeuTWlIsAnafcJdox85g///AgmXXd6/hwhuePgR9
mCaGhpLx98I/KifOvKWkQnC4Hl7GNTq0p/pMhRR7eUvGdp5Y7sKKVi4uRoduwL50D+DRfA8tbOUz
87fRu+vaKhhma7bG7sKlLHt7ToZBXhBIbT8EI/O5nWS5UxZ3g+nyoJx0ejRV52ZW2sFgT809x7wX
10QGbnHlJGxzdQpsxSWCEMNIaDgy6RpCPJul9U+PfJCSiupcAHkOgukSwVWWiparklIlBI1X4iFN
G0LH1HNLNTrOY4n1a5P+1l96/Bd0U2Vl8qQksepSI8ACWYYjQ36LqntbMmki4lyrXBymQF6val/c
Loc/r6xWzFBFsSPbkq8SBo7n2WjJwp+JKaSDFvjIIoZxwizvfJbH069iiML/7cRrSVsa4pQTOqPU
N4AG3cQOHicIftgRp4YDo/mXsfbEVMekVvdFC2JAMDIcu4ny2YFoXpEtt0TLm6v086VnJQ0a2HC1
QF+TXvxXcvh6ciHdsFdqSHActlwRAKqqyvR80gNH+0Sg6ltBtEVHgWk5t9VhcipI3AcE9S1Th+zL
pX2kyyw19GUPaU1euIp2zKt6a4EYcWEMhv77xogbor7hTQnU8acQeT0OMEL7CaHXzooLLQ132f+3
MKDu+oIAndN05yDJvEJBh3HGH/Zm4y77kMaqcJcr2aFnl4EJ4y0S06R7TXPVNm3UDMHtYvBFtjZ0
7IG2riS9pzyTG8eLHjPAykhpLm5407vg7C4ZPDCqZOw/Cp7z0zizqSNPXugoIvMvb+SuWG1zWTOQ
SmQ1Jzj5sFOw98gZQCzEKztiPPxh9OpXo3Q6QTRPDBp9i2igBMxNkidZrB7b1S8geV2AiDGnrrfo
+wiEThy3H+WGI4/MnISqjvXwsrvh4mFZMno3ypEIqkd8QWCtuCiFLx8JWnaMTKX4fD+Hi8gSQ4Gh
MPXPV6Uk2lQ33IIlQ+8EIneF0yCR6qSDIwrcxChfO0j5ObFC4ZWJ0B/IUUsWGarsXnnO3yhTT0BC
rMvS0t1+1RNz2OL3zgzyOhze6+0/1EDFaWSNtoHO314W7eFGuuPyKT+YTnH/yM1WM/GWhKwchNrt
dOoQpJ/GcVpT07b4i11uxsrxAxOP+yBAYV/A+IoPyJeZfJ0XaodzRRytCY0W2h1bLoVntrG2i87z
zTqdTUahxxUdPzuB5aw6X6lRxp2h82UTKM62WMhDqaQqLLZxBMPYI79AK3RQu8rq+YKYrXx4Ma7k
/LVclHr67zXZ9jOJmq/cpaia5VWVK0dwLzc/duWzxowOFmgcJ6wq97AHz8uW4qjGfzPUrVKZFu4H
ApcBUHQA1IIed/dgiCF3AXTnzpbPnd2gPbH/ixmXdk4HTbx1t/UfjlSchsfaYmR/TbwiPTi9o3+V
rUfViJUvgDFgeSQeuJAdxI6/vJD/SrQWv0gcC+/9AITs5ucImfI3TLJxCCy/gFy6vWSx421rOBcq
Cdk8U4Z1znWkbCqCZadqi6t3kC62oR0u2kdd/1wmDv9bXPOH+IKVDmFjEQdMHAe1nSKUy0/+s0Ps
2qVOwfnDKq/wAwkdJRWZnIm66NxZ2W5xLTTc0nbewOrHTKaGt1hSyzavXYulf3IRiCRAL7a2ruF/
JblWuBmzTnoCPWUe7WQBhTQB+CJPntM+i4AWSBQm+uTi5mpBHRxBrVeFbzpKEmh+iEbtZ9PDCTy3
wOSxlB1fLlNQQEse6Y8Xn1KGG62gs2ODn2ltBWZQqqR25rY/kQXNAV9js3O/VxoRpTX3uEEqyFBb
1RaKvP1DtqoeFII7ascrvNS+BMwGVhIUoPCsYdyB/Ehj2Ov+pva4I4s7q3piNAlbt76+7dZTgf2D
HtPIbsCnwteTmiK9C/7cZ12gPHZyaj9htUDYH7gtkpdnVIrLiRMJHyLv72h0DyDFmf46JY9rn8N1
XeegNqcsrwaQmdyR740hneSsjBFaxM5f8ajqT9Dk24DXqKt3vRthjLhEAg7AJn9fSl5cxeQUrzwW
KoWEntr8O3QDf4NVDOtsGVUnb0SwvEXDBasAHMZs2F7pWno6EeFbq8V51jyUiQXGfWMaBWEOJTyu
1TlXbtlRsa74NX1h/KGQLKUq1zvGeUmoURB12Pfr04tMEtHpbDaYGVmMqVWU63xHlaasRNarKx0y
CT8E5i7KXoIIFGgb3zymi9IkRGDf8lG9yYCgpDcBmuAevVPY+xE7L5YkXXuIbIOHusohyw/FSOqz
SDKCuzM27KtCZOkO6J/50SFg2U3flk7eXSndTbpTrIw3Khaqd9kBLJ57UpyXkadvEE0ZUwUl9+3x
8SCoBFFSkjlXYW5a1zV06Sbu+tQlybSOn2ijN7bnvOpUPaXnkdrHmpaY46ofS4Bap0H0eDr/micG
MREjbRjCErpZRovLxHrmUVr+0Ku4w0leoMdKJ/OcuWQgsau7/97mEhZ7NB/FzjwcY10h/UnfLXCE
uN0p9wCr3sv6XltG+4j9DFfbcm7gciD7ThPrSXw1TnaZOMv81NF4fiTAyoWzTs3TAVYC+ZfVK1Mg
nBVyOFzvA2kXj7J3YeldJxBa7S7Hxqxj81JkA95Oa8CrH4u1E2LdYZKvX0LmoU9RD2eBsz5dTGPZ
Epj5vuAPjlGQSIzbmJxCEDMNbS9EU0rsk0xTXeJozdeCK+rT3XmSOjYSJIYdEzfBZpuhQFcYgVai
0BwGrFL3Hc5+eR0OLCLLcnqLE/cUp+TccAMg7G92a8OKd+vnvKwxbMxgSNqgXGlJOM8xOgxgyz1C
MI9iZT7gxCdn6DA/1mhzxJui7HQrRIKIYL6Bic7vbvqWROTfzTt8ZIoavyogKiZ/St1U7gzeiRMj
qsvIGfqpPcDmuawCHCUlk00t6lOx6HuRRatV3RrkaAI9ZJ5RUoxddy83XVtyJidKS0w3WiPNnLNp
gGYFX/XNUUgewTGmHQ++6gdPTE5AUA+LsltpxRvi/pEIF5NVI2e9YmAzXM6ISFZRKo4c29PDqDQa
9G2flYn2y2YF6zt736UePtgvrVGDHgcc3wDgNJDxj4Hy4rrlMl/eZk8DK9GNOXbMHVyWQBQNZ16z
UU7AS2+8lICcLTCvXuDU/WsevkknDbKq7ICmORLy/VfWRfLgxZizj4HrKsj8IVcw1n8E3iolbXk3
ilDyQlR3ac3XYiFAYpUAEywuziI/DDF/dqU73Gq69dZcOvcVk8bj8Tg1N6HR5slZAqwA4/eMbx8b
Ql13BxKUMeLA5RoBt1zf0asIbJf4t/MdL6L1/YPkcm3gMHY7DSDe1zfyblf3hX7zMGycGhSaGZvR
BJ+ufIkHx+X/Pmb494dCR60+//TQJNXatC7GKLlzejfT5Z1hd5Z+czkg4Twoix2Ye5wDr9/UiR73
GYsFGtnSPkwHX5NHNr8oemmdUtlAU78qtatfDAqtNslzr8diAsdUK+fWmC/i1aI8/VrrSooM8u0R
5EDd5h2A0iJ3wmy4K3dlumsWg+40/S6mJ5RE39rOFxJVxnPE3hlL+y86vin+ZeJOC1HAolCTKQFP
Moevr0oWnHuATSm+HHY3J4BiRy6YgfOgcM7S3bQC7ZGSky2xJImtgYphhxsmY8RG/gLUNTPq0TTD
P6pzLrGJnJ5P6vYW0NeNMVffPSjkiJm5SOwVrIoU+pSYjOpIwcrcdvRB2rbjNHVCC58v4RAZA59m
dOsZept01UUstI0bHv5nxVNtFRb6vczrpwO5D5fryq9AefgYjcb6Yg95AA5DYZPgDh7rC3uyIbj4
HBUzBzY7SngcpViEk+bs+yMR3oj6HvxjgR2obC147scfvQBKG9t4qtq5S2J4YftyyUUWqIrN2iGS
odw+D6l75WkwgF1oPPWZq3+2LUi927zfGb3+wiPM1Le6o3wZHeMmmJktyngWl4D9ej8nIU5I0AZf
oBKHdXHHN405KJjUiK0fZOjQSUtdmsR6QqTwCLmVsyYpKjyv0AO+zbGS3/a6ULc1H5Wa0DCyn/KB
MrTtDyX9bztQsy5oOK+7/jnsI++xpRyi2ShGgrzoRrVYN76XLD8jTvWB6QIUkc3VE9+FWGKecYA8
feg0t89Uz54hgL7MMjLArLQXdSDJPstGXuA2kAbGjzG7e2k4xfBlWuy37Knw52EaKjQbABlzk/9T
GsUZzJn/3ls0w1q8PM2sx/lRpHnhvEUM70MnR45BWjU9nuDyz+/Vqa5rHb4cgcJz1rK3JIL8FHH7
26PuhecQyUm1e+MP/2Co8gydps8POQ/Xe0B5chJ3FRbKHh0CQ2TxuOVAninMCh5vaUxxRGlilsf/
nEUT1hQmkGOL4hXYOjP5JQn0lt2Yb06uNPaJJS1K8UfrzSrql2iE+bSfEaNCiDzY/9V8FSDcpdbb
IQ48YE7UJ+OYpj7o8Wcmy8IiXk2H0+K91uNkKLtiKOyP69EL073UWI5jkWV506Dc+CQShqshls1a
zpV9itS0JtzBkNdQy1sPokhPqfe4kugYvkPkaKqXgNDs2Sz+XWwKajMxlCgdmmsZHX85P3Mm/tuJ
gREEjNHtCmIu2QFrfiIDUZ01sikH4FNisWiooB1wH2jMcggQkspCvPrXKGWhU30UHPL1ZtXWvzxm
bZCGOJK0MJZG3+lqy6zxKtzaoaq99B1+dCjDjmwrkh5bgAuS76rxH9p8aOQFW2C020XgaMQp2Uq1
hV/MlAeC/qaZ2yH4g1nUpRQxfxyve1VaSc+yBG78XPNJU0u13yvVx7ICbGNR08bhyl1Jem2MfDU+
wqvkXGw7vj4sLUDzKfWWwWPJlAFrjNHDVz3PkgtmuXxDhtQinuOzU2Ev++j8AdmdXewGTjsCYHd3
ch3Hxrm449kYwEwOji9ihhr+OiiO6KfO+wR/taNJHpSpgAlgbc9wvTp8XfgpieZdsO7iZ5Ofuqs8
5k4i+kLchGawRbivhonxZjfs4kliSUWLorEICrWeIVEjBs67bbsm6ZjhUzQxXxr5JXi9aArcEPkU
ydWFj9UN05PMGX/rUmClfaYMPEliFZH/RtzGDtqZ8mpS7oY51aa/fgq7fcWgGM385lyInyDCRw3y
Uht4b5SiqIFvZbi8BlGrZ/d5ygMh+N+cXfT8OisbbC00Rwt1aKIjHw8hVjrrW7f05q6LMLkuY9DC
zP/LvrJLu146SlMPAGb2PAzRFcbBWEN1VMpKTe4CIqne6F4/1jjYKS4c2UuLwErcbZDb8M5PsiRp
zIS9x9Gkgt+fgNIIxxyaRNsjTxAxj7BJLAl+k6btoTYhn2aUJm7QlLEPnzj+YwpeOH+Hxi7xelcd
Nv5ANxLE47r+vGSDbH7+liDXzqlJOBzC8KDIhB8UN9aNarQtQ6WWG7mWfbofSKRet846iI4ouOvE
EVZB2gLIvkMMPIU3PjNjydvjkEsnkCkGkb9lEjZYGpwloNbDPwmkNNW8LTlGaSHjRB3GJrVPOYWl
SVos6Kly2jBY4M2SWbpEf5lO2bXsVrN1no2bkOH9zq2uiNjaF5av7SVJ//NiAFZQHRx5YP+/lBRA
C78jolss6WouxOLt8BZRoVrOzGqR1eWMv4V7CTxzs19c7DGVvizo8hNz6Z2l8SLEgcyIQ7LlR3AU
RM+MAXmXcECioOl3hEy0JsMjnpD0f1wuoBCt6Xe0nnSGvYrCcURtp0fD/2j8oiOW6k17cXXOOryr
9QW0KtdUujquFXzzAMMcTglt68JwOJ5yBHyz6+WtwkibuXv3zihdKvy7vSPGXWU8wtZ3kapnvFJP
85Zh17iDfqjWvB9SIAx49txK4xR5nwmX84mUBPGhpk9oQiuCnqbWcv6LHI30fjFi3YVr8ANQw3Lb
dEzqDSDqjwK+wKMTns60JTu7xgWnwIejtth11T9SgPbD/nb9Zg8KifUzT6GWXvUJlMTriQO6Zf8p
mWBKqdBrcNtswHl8McZbwVST9irpo74/+V1aI6uQAY2T8zzBWbqK4bvC0AWMM9QUfVXO0ZPXBa2i
l4k/wywFtZ96fWDKIGsl4i6BuzxaD6/Np5SxFjI9r6eDnantusRvmzGGINWCSPEw5XcZP3Zhaxts
cCLrlcIn0pe2jjXiZ7q4mZmSXZJ3AvwnToWrpHZ3cgVAHHMXd6QaTIQziNSUda55DI1Cuf5UYkvC
eLl6ND5OpkF/9yeZsw9T1RyW+GtM6kkoVZiee1sX+ITraKXC7Q8N5jKM8MIzkBXXEefDnGcrBk4V
3z01zwxZ++Uhoo5VbEZJFy/rh+cQYlQhP3Sq+KiVguLfV+8RO4pU9S+DaNGA8yKxe+TqQpAA0Uxn
ZCtGgIm4htPbZj67L2AxSTExTH5ezLavcTCyj/qvU4eB9dJ0DnEXbz7de+mjVAylca8DhlYW2dt3
dQPTlYdOLp2DDPJUgT0lf2TW+uaPfMBfzd0Su5PrgOK8Wm3V5s3+cHMWuXDGI3DkB7PpI0lhEEzh
1QNNzpdiGr95wxrDd/WRs8DEL5g1aVoP/5O5EgUajG0mjPdq801y9ZVOBwHzq0I7EdxnVyM0jS4x
7FWOmmnWd32jmRxXbDFdUYG/G+axN0ZcYHkfEb8c9ZO1rACoOOL+K72kS7eU1QXayhDBJJdOCdYU
wbMeywzdXSu6CqX/ABm9hLiD/BSuQPtdBoD6TclTTxbIsEW/9/8JN6sYRo3QDNpKwkaW31weZUw3
rzf0ynB0ZsTwlBvvXuVd0nh9jFFasr9SO00SjzzpV7swPnymNdJeUnBAK/1CS+jj/q1xaxANb7Gj
04Bgn8Y1Qe0evbx7h8LGDApdx/fCMQzGmaI+wCVAGB98KYqWyUaGs7SAEBKmwUaHjq1zQI8MjYrW
KDu50eYRMT9+wBFbSmftlg8xXfeL3OUVGu2weBhF7N4EhVUZmVq2Gubhg/zIAPfPdNZblBx+CTEz
gdOuqGe4GkVGJ+4CYAiC5ENSr/qCk6LNREiA68h1sEPCVg8gNY0GIA4Pc1bmZUrJjvYzyf6F0cO7
6ZFrnO7CK2Umn6jnGtp9oauIYtr80oZqqoYDk/AhPz2bRlFksnpDqfEmD25dsn3u8EP1hk5LcXgu
wdmmK9ypgPsG9WtYXWLuiIUl/nQjHdcFHFwQmDZbFC4wKfDNq/ob08sRbgFsAuTWxvSCtPp6TUcx
TP8jRTuatJCWB4+xrJg/txTq+PWhAQlB86aKUACB5EjLOktxVNDKhXjPmr3DXT7WGFlCy2DOS7b0
C1addt2SWU1NNwxhuOkuxf8+8e0aUFYM1fWUuyj5MhqWM0tv4AuvIqm3NCMvlq/RFaZgv8810VzO
yyjgAjIGmYW2HhHL0wgJMGAqrjY366W1tD9nVsYu6Ly9DCRdPujru9u2LjFVpUbZTSBrqP/b6mvA
NtMzvN0klT43a/6S7SK93WL3MFfDnYiuyPrHBd4t1dAick9Sia/vKv2b7oLuJQ/JWN5gnuHq1oU+
Ttoc1/pj9fkyr2aiat9QYJNmb7nEk6Qc3rJUGsfl9Am/ZPrFsJvU9knq7OYL/aeo/qCJsxujQ1Vx
i+b+OfDy2+VCgSG6aZB9z86Qj9Tk1sWufUSQb7alf66miR8PjKPELH1CpfXTHeIVBuu5fu3xZZB7
3Li1IQ6Gx1ak8mbZABUvpu763S+QPx8msAxEPxfkenuHN1ekJsd7LseYukCx705CbPXR+trSp3LG
wKTayT8Sa9gPbAA3jmQ7wqM5bXA9ljNvUrAcVAcKx/woviRqBDCWWtP4QokixLPo06HQ1q6ZMYW+
4GW5urdKOd+WP9mS4GNVGWSkAtlZq3x0QOB6bak/EK06njJMypLXPG+NokdYE7DnBJTbd0Ef/P63
pepSV6bHNanz8kHnYYADwZPVckOKkkafDmPqxg7xu9ik+UBHyAEFGkJ0jeiq7j/lEx1h2O+MI8Jc
PdFDTxv8LcHFBrPjteesaxQBbm7uD9w1DzwfhFq9qw6IzmGAe40TXAoEqzER6CHYn6evcZN3NTMV
fC2TGCYTe+TpRuHIewyq1BSZB1TkfNcNe1yHXV4w743/ZJrv6crjie4sViHyxZ50zcRVbz42jmRN
f90aiG/nM/CPmVusmQJg2WGk68UeG6uz1IGNrWaVbeyjQrnnQJbpctUcHvs6++Z9T0WE6RKqEJOl
6SoEYG8KDT0ygytM24+HQM29hUmi+mKU8MWtq8QD3CgMXp7rN2MK4GscVbimwht3oPQKUueYj7S6
yuoN2liXrr+70AlJn4kQ40Z362s9zoBbEmajWTlgp85ECNeyoGWNl6IR5itRanQsSKo2xMFnWejs
fEbGYDkTeyf/h+uaihLwT9Kk7PebZCt2EQ7uG7yYpWAlJN75gZQGd1VOcjJtAzxb/oDlYfdmhubc
y9m4G0p+22qujScHJJ4R3s2SVqGE2gfgqYiIktTeNQYJZR0zdSzE25le7kHxMt8dmak7sqLBbCqK
/SB/asNl5C+cta4OJCWub/OhTmI6Bm2rPjA5hKzBgJ9wSgu2A6OkEeZmqCmzvJVe3yOwJckHB5L+
xAcrNXmnkBNlbL/2GjzIR7ZrnbiYEo3SofKHSQhdh3Ywiiw2lre8QvT+FmJXRsAuXgLEqDhhyVbH
kTCFjCRJtL3Qtd07tILNEnsirNfS0WW8mWMaf0RGpihKoSEKKt9snBCovU3XrAQ5sEf1F0HVyOVu
7JCS6Wshn1Hh3h2dD1UAWsncoZ5vlAlWoQTdoDTQ+9Enr96z5MAvvarA5EcvFLaYBMHUilPudDtT
/A3sK74lecE2k+a9P9kuJ7kqPQm10paKWzO6NmD4jjQ9rzEYRSglZqNSsDmBAW8Em2VSxh8imWix
rfO+Nd1AJqQPuboqQudLjLdm/MbJKkTRbNm+41S+VRiEhIsuOg7h1pNVXG/gIf9eaOorSBQPSFcj
UAvtGrTnQUNk+3d86pE/3NI/4VldGIlzELM49wf/mwfgUHDAOziehGS+zTVUYKctXhmCTNfffqYS
p0/91+YRAoIwEXJ7ishVdiqxeFXWGn+2uYY0cm8LpTF/ikQpq5KyjKKQ2aJbSJV2seXt6hU5oNHw
JIeLIDJ1Q2+uJZPeXpHhO5VkY2BDAHZsQXZ5Zci3BU/KfSG6P+kJmThxulRhv2vKmtOhnXBwMEwN
FHoxnWFEWdy1dyOru6sFSnGiLo+qbrD0b3KHm+rlGVLm//4neUIJz7tBsarzpNaSW5/rAEPMn9TY
c9Z7T+931u8cOaxQkoc6Sq5WAhs3PQxw7snu47t1vNKW7ZCNRYItX4KkvLTdFeSH6BnJ/ehFGtXg
s+AwcYeIaXDMBQM9vB6SglkuDcJAsv3D326+yLeYYN4levohWjjnKz6bWpP4FZRqIg6XECRMRdxF
dGVMwZk+gcah2R+jroUlMh6+holWeVCQq1DZtjoLLQIWaDB/tgtRum0/N6NJ0ianyRHpviPxLS2S
dV9AGZ/HUIdMBK5EuZVsVnh0x7qNNCcmLl0+hP+OmlBSg96jIFxjlHPyYBjGePzBnsF6QKl8JHxi
j/o9rvlw/m02QGjFjFz7PMuz0iO0p5VjVmt71rAzx3hC/tD7b1GCdk83PCleHD/p+oIr5X28iDtS
KMbuP0IE2L2o96T230x2voo16bo5nePL7jQdrWvYOjQgdv0Pjz4xsrmWvMysL02N50wgVNGLP2T6
vPiOu8NW8E9TpKdmUlO3q1cAIQucGVMshrH2n5G48NjqjkRJRAKoskqOxjKcZDPIR1NKtpnsxoqi
hVT7I2Xq4BxnN/t4wS+sGcCPgB5T4KnffrTb97xjNRpl4r5dtmPW8HKCB3XBuqMB7/dzz5x9IqyJ
VhsiYCmn+Fr+YFQX1jYFJg0+RwkwD3r3P+QVpfePqZJgHfK0p/ejliUWCpeUtCu7e4M0JoCb+mkb
HnE5oSGM7faoC7DwuQ/9nhh4+ALvc9ATAn4/IYKHtBUUWRYe7gCL26nRsFmmMW3U+Orkvw0q6nvD
zyGbPfH5tyLn50EpODpPzv8PvgxWp4e0Smf19POXaSP7uA9T6XszG75qhLYNlX8JJWBTUD1M1HtU
ZX2Q8tmMO3NEIdrgcQgscHtwYRC1Z0UaoqgmAMjObDCZnZoWuEH5WmSBbkuDN6vqJMxkAtGBQzZM
6CE+b/8Avp4mu+CrpWHSpP0gLGYzQGauRRBPpu2kPLiOyXBXDxlMAuAIe2aLkckA4Sl85TnHfpP3
8hwySawoF9Nt+CuUVekq49nKKtP8dJJ+1zrFIhO1/m099L9om4opYD9PlguQN7eD1e6X2thuLJmI
Tq3Hf3GmGHjUdrkiOtT65ChDI3hJFCJ3xi3EHzg4wu2ZEWyvebVYZyaZ+yhh+WJ1G7OcNeBmWSzZ
igQNB23coS6tIRDrkdM6Er/bQfOqHXm016DqbekoKYPvvhl9qrupLMAYBSsyA+JkxqkTbEiA1l8o
eeAF1VdYE/Q8dJ9T95Sps1f2bOIzgJKdpHZK2Rl3L9nZD9CRHE4YZPpts/E9Nqni4XLwplWQRpu+
n70XW93BXTs9bH30s9otZUp2/Urx98Ifnwuz3O1duYneOWmGrPtbrBsmI1B8Ew7IzenL9m1AW4Rb
ylZjIZxrZOEVrK6elb/qaj0cOvLKWZBK7PgnlG/poq3268WWXKOhRy+30ajncZwOSftKogf36GZS
mxs7rfzxl/cf4yk0hCDQ018u0yuJTMkrljRWPbHvalfXNsyA6AjR3Xtq414zcQPoFdY3fVz5336C
bbyFJb8zz03UfxgmTg66z/byxINIH760OfD8gJ4FVfHYTqlUaJebTq345jygNiDkGXxiRBqKMQz6
aNtkHfLbf8DYgAFaZyTv4Q7azgC8EvEKG25Y8v0Vx9tMhrij4zJlTRzOzKwKIv+Ullz9pyy496k/
37K0GJTCQO57BHnvbj0IxFoGQXG9Dmkjip4DpH8pruZ4aUuYLl/MBcY3O1UhROUdo5IzqilM4nw+
K3jo/mxq+7GEznU+q+edv1gFljforSD3QWjIl8s8D/n72J5vGZ5Ndn5Xc8wKmLF6r+SD8fShvdpS
SYsOObmwo2/w70azPAdIZwjllJu/wrflJelNZFA60FmfnrJMbzRhRzePzPmbVMK0vYwjqH1naqGl
ijZER80CiCJN68vERM33MQ/VoUC2DDR6siN3cyMMYfvsB8o7b7SQLHBT/wxpL8v/wtPYKCASfgOM
rj6O9P1Vqc7bfj8EA46aqK9zfV6rkwYyA/aCvTHMGHWHAgZBIq95QHanfY5oBRWV+ohD8RQ2d4xK
IaVlqoNY7j0Gga95lb/spUxrJ3CsBqRDIAn0wvby6lEZ8N7ltgKvt3ITXdstBEb2gernvBoGqLt9
K6jcSBff5fFu91qQzzlaDi8+ewylVIJRWGjum/BQyQzvBKqy29iyqLkfp92OhY0pH2oFaFAXElUt
JguwRSVHyyptkPQyWBSkxrCnyq2Ei40GjhIyQes5TQQHGmSyLfdzmWgJDlSYvvmQkh5Mnp9S9geo
n17v+WOzditGQfrpG3XKZ53ubmiqmfecg1cVsESz1JweP4TsctaoJCAevgcoz/agEep1bzLguY0y
0mItQe1Ot+oznicFwg+qCe7NpMYmYtMaxsO7i7IcJScCm/Liu6wmIT7qYCm/Q3h/blI3h1JSElkx
7umzsmeYqMQ/RraRgea9UnFJA3xe+fvt5l33OZxEFgzlIquS6WRPnh1DuK+XcX/F9cvo4VUWI2CM
3GWDuC1drCg0WrEmWaxtlSIp0WdnbCt6BB6o35EIiIVOVI8jUoltWP/DfY5v8o1Yd8LJuHtJie3W
FEq8FN8QbKDzIKwJBLM4dpPwZMV7YNahXw9o4jky7yTSJj1sQ574KdZhOMqkYApM7U2cwsGrfTlK
9gtKD9pshw0Aim427aUPQHPDBIGWzIWX7BJ2b31z1WPybgMiT2v5hTJIA+HI3z314jHD4cCoNk76
46paAsF00eSimsoc9UDub9Q4ms2HDykiWbZ5DUc7PZemAesi9JHvmxmCvLG4iaJje65rIIVJj+q/
bvehy/Xhd62CvjG70SLJmtw82Wd3dzams3Im1YCOc8Hiw86QWcIoPKGuu06GCF/LkBSYqRj/C5nb
LxG5ho2CndQU1RgugOa/IfjTY2iooLk/mv4V80ceNjcobsuIcOIibQ5/tPnIQM4gbmeYZNEqv1jz
BlTkARhhBK9YYRsBQtDda+ZU4LYXRdwqkhRN6SuZEnj+w19nlsZNEv1bOlk/jDGEdpzwzn+HheRZ
oGQrly1KK6qU34KHKoGGqnnrTidmhzftgyms1bWPc8SmMMP8jk3k2qEL4uN0QIy4OFvEZaF3uwip
R+6IGRYE9cth52dge63tPJSYifS4P7g2bfF5t54tyhuSi2Z4tnJYAx9ye/cAw2zKgTmCX3QJqlWI
HNysrTPO94niaDh7r7z9JX02h6K62o3GRquo6Rny0ibnUuzXBxLC9ovSICklJDGRd3QF4nIPBV21
EncHhCwOFFwLwtIgEZHudDzUA6ZOXWxgYMolMTQvM3sKMyAg9TWlMKV9ITaHQmzq54x4ooJUqj8Z
gTWu4+o0QCXRpFrTd/2kRWctw+3H2aT57vQDSj9YbRIoRyZRyHVxtNaCf8foNsgews2Y0LP/EsLZ
4c+MuFto4qQGG69uOn4MjZNHQzNcc6BxY9A1sySXwMY+wpR7j+mjPDU6IjpmgyNsLRUslNmSd6Cg
opUmi7t55ZkYMvKr038HGNxcCBWYQbPBW7sV0tNl0HzSQLzJ19E2ieUkD8Wf/KJtx5JilvrwHqxO
zC/XbZ1FA0qXqybxGVJzHen7BTliGS+Gbwp8wtMj198bHT4k9m8H9r2gUNDyElKiyIIZL4FL4RRv
cLzfa627R8t/xOlILIcfbOkLJAtobLyop+fx1TSRqZIyD2GatJck7mWkQ/PVntLUmrnSvIi1kSN/
Sv17zMAfh5reP77jk1hVCgZGpYbHmHA4ZLizBp5ZfZwJr/lEeQJVj8C9AaP8vZF1KkISq6WWBJga
yf03VdykRsUURoP0a6hEbPEXSB/dyECt6CsbA9LMXktMhaNejMBG+SYLLDaRP8y8nJsebu2X79ej
RG2KQH+WgXCkrbCJBQgJC5knRkk+6mvJyZEsfGChp423YpgBQBAZeov01FX++h4m61iQAm/e6dfG
09JlInBqpmFopr52L6dlGnkcHttYTKBMYTJ13yZv+AA2pRrNBGl9bZHC3TOigTArmpkg5R2kMImA
sesYbZoOIR2pKCwHUkOvreyRFBbBOriKMXBEMUEjJqjxOT/E9sWO8eR8AIzUsh2aJhSX8z5UB+Nt
vZ8oF7bUDDv3Fn1cKjxRJkAVPiJFxQdsCpSsAds/C2uHrGvGAWulcD+UE0Y8OB68Knw41K2dHQXR
MklQTFUYuWFkEtJVRWe1VF3qF628nF+rMh0b1wiqBDENeRNMKwHp+ofI+vxFFN960+ISXNk69rDq
lA1gD6UOjVVfD0GRQPmZ02Dt7hy94w9v8GATJAlcLyWIBrEVtojawYSQdD7p4dE/GfhXIddyFHJ2
0L5oOF7mrGkze+3hDr8ywg5xQBtHgeDZ1lMuGHjTZ/Junb8Glkt/5eqBBx/r4zeWfPh1bGGHCoNQ
Un4CxTSaDrlsfPVS8tP3JDtPXtP2WUzPb67LMUS2P7lHKpZNqv5v1we0eYk2ErWSz2TDMjCD3bmO
EXsd9n+tTGp1A4y6gHdbKZ2uc0Lo7bEmgUHkSFpC0fxfYxpV5Ca9ne4jMr054q0LiEDNo7QV49I2
kVfdKmsMM3GPte+B/uy7Qwk2N8rN62e/j0xMUhqMzDPv8Ct38+SIndWP9cX7tIOJi1j1N+riIImA
d7sbMqL0ZDZ9M6fYCqtksQL1/Ghie/XdXWULybieJKPo6v8GH3v/Bml05CXW8ON78OUHOnRI9/tj
GYBARfK91xkrNSxgmUUHMvfB7+qCJt4hzhuzOEXquHXb3eOWjYHL9aQCAWkyM9rJBpBiWKYwUjLb
MCGFiydiZeg1+EGOKVPEcshVps4DzS38EIu3KVqFUEn/BwjLH338i0J4+/VGgOB+Df9ZXDv/B81T
ny7dghW4N/elE/Ynr6jf3q+RA4sGd2TOSe+g3Fj9B5KT2QJ35/02eQr8QtZauFkB2R6GewuVslsF
OVN1dtf+iHCzzt7GlIpHgkpGIWnRT7VyjJ/yNtkj5ZG8BbcrP9A+FTlm4nmftYr5D9a9iodHAJHA
u1SiWRCXx9i9Sd8HdCX3saCjrJeAd0PwkoYn9y9lif/LSdXhD2TZY0RSV5WT5kVBsexbspNQYctC
TJ+QGeEQzs4f/21q6aCwmd6gIJuPXfVFUfNpm3YQravnobJR3QoB6C8vuvSE2N9abucGAENNTnkx
oIK6KHNGPB/a/8/sz1k+cHSTS6DwkfMLprIbfT4b8Fd+tYPP1D1eUS3v1dg6vPCU4/qHgikyTcuJ
94wg5xMzzPleNJXTIJ18IrjKH3NrpZ+Lyse3eYtyowVdhy73lN5IaEwHw5GZ65Cq4BlJNxwXTWkJ
njA+uM08qeMs7Q/3541dJmE7Hgc8CQusZxKJbx2j8Yd1osCuN518j4fem45DnvWMIKVNw7JTNfry
6p+xyMmL+7ee1wIwSW75Yic+VT3OfQqfYmCpVufWgg5G+L4ObXuZWRfl4B4Zqxdb/iACsRMIV9zg
cRUXejl8HknaoPRkB9hK5X8lLqBgwAnH/p8zUX7+AU/A7z8TqbK8kpmj4xLJCoaIGzpHya/tt/30
q1Y3C7o4ijSkx32fdySLZK0StoHcC0t9CatyxYBfh7piqONUYikRREhAVITs4fOlblMHg+c8fXYt
Y2vxbTJRp8yPTQqZcDhv6niVmDMWInd0iCIPFIqPYcDlebd7wJTJkQkBfOZO4ZsDo9eoSkx920tY
qSbuhGtJIdQhAb23ifjs1xTuktPgG57jwWH8gStdS9yph8iPpBwMdksn3MDaZOmVfuVnnQRjk11c
ClPJlcUq31z9UWt2HxpcZOK9wa91IB9pu6ZVTOAjdDix429hMCglXPRPM06jScp8pN8W842Z/0e4
N7xxPs5WJZvRyvzBU0VDVgxqs6UXyknlnEfyBxTirhrwf8ZsE7aXe+h7Sl+RrVWf7im8nmZH5iwu
b9649R3Iqy+4KbMv1+NyFWNlSg0cp8VD1z0x52ACdmrDv9+oYL5Mp2BXaz7Pri4m6A/YO4hVbUHd
olatJAQep2dyodhn7sOGPJ5Y6ZYYYn+xSyX+MYnrL4iu3fqYkwq3LD7w42+H44tK75TlLG8JznJK
/ywYdKkd+eAgMezB4zyg7RRSb3GujF4FM3AvV0sk3W3hIhjkSGaFJf/MAnYNeS+x5DfwEvnUEtES
2fIGDnWcO94FziQbw/Qyz9Qn4uGaEkt2NSBW9ns5mP/CB7a5Uzu4hUEbmMF6+cKwl/Zc9fnSpROb
Bgs+B/6MmwFqyuEkkKSmyphl7sbB7QbNpDgakZlVGy0KQmFo9XIRkJm2jVI8CPZEAmTNZLdEWTMV
EBL7KlV1CbkMdPNwPykf7XH4lVzzHpz5Ka4LQcwvXuPbv6sxQQw8Dnx2MQLTMW/8KNRfLrbwb2i6
L0aCYZed29cAc+YnVl2/+AdfibkYZYDHFz/ZaUZIHrXAy9CrR+iBeTY+Zi/r5EgzjiT2EKFUy/xj
OCD2bWOpm4rQpPQncHeW055jo6VfSUX/s+uotDgsUjTOhC3sarnULt9G19rwqgNXmy5rVizmzUej
EBxm2v0L+ymcz1nNcHklK6RByQ2cv2xXHLW7S2xlvfFKLWMTMAeH1l5swi8YaIgkCNIPaKO9yeXB
80Ok73vDmBSIVdumuczd8/SbnECRiBDY3yhoYe6Kp921LS7i7EShWuYJGBaukmTu/Pd7zsJ2Wq36
L+IaWXuBPID0FtaQ1VILMZ2KEiIeVro0M2sc+JQj1/2D5aTALuVHuxNygBgzlQIdACgTzMJCOtrx
G9wlHoqzRVhT60Cbj7fES/LePuKsBmZuoKmreb+J1+Hvirb2OPADiqwcWWsfbiDhZkcsHpApLDeS
t79QqT7Y2C4iOXh2DQkeXtL1zgYScMGB16aG1pB4s9/8rZUphKG376XJIUBwoV0G7zShAaAo0a6X
y8CT5cGTrJk5z+irvnpgA9vnuN/rZjPz5jZStGXQMXvW0G9NVi7I57YUaMVZ8XvtT0F1G6zQzwhQ
s1cYFS+vC4445jThXkQkIMTaRaptcrpVz2E2S3oYj0RfQ23uBYktLfc0x+PyaDcE+WHaoTvpG+8k
AZPNFJrw/S0aPNNIyxTcqOb6ofRYgVC3Ag3VjmJ6+CLnQks7gWA664v9c6k6sUYdgKsVo71WzDgj
KH7J936tdoVRcoHoTKHBKhWm3VPY3iyRw5tcsui8BBaZVJU8F37YDhslKSEZPt6RYotNyDLzrHr+
qfn95A/u4BxsB4nXW7mn20Oj9iUk534yrBoZRYT7gyQU1XwydqwqMalvqgRH34z86FR52vdlnvQP
QxKn20cLt25dWG1pR2T+UHX1o9YnMSZMYl03xXObvqhO+pmJKswuZzqiUAq9CmfiVxTGlaC1sSm5
J68wwXfSRuPJwpXz4KsiqppGblIFAGedD6ucEEuL/Y0zSSFn+d+occ6L1RH2xDE31LvFXpiNpF2D
lrwItFUU5nwSP1gRM9HkApEF+qPCrRnrJzuhQPwv0Dl9x/y+hSHsEW5Y0+3KbPHdQeIblV5Jbx79
wwVqxmY2oGaCs6kV1eqQifu5cWJOkpmzDuWZGC7WUkNgyYnXCwo/1IW7fBPNmLgszV52SOBeLQxJ
3+Y1dFW8Tp8WIRR9u4Df3QQi0ico4GC7Wx3po+0WiSE49hpWgFn54xFUt28RBKchM+XsSEwuNY9/
0jyF61EvYI5Jeja7kqWb0tC1pL8328nS1SgyuDlY6QGVRYZs7XwNQghxdVDd+WlL0OyVINft+Hhu
kawa/bryyfax7RO3bLz4NNYN2BwulZCy9DNJ7mtb7sQAHTnSJTD7oD6pCM6gz2qCmlZWEO1m2/8v
CrpEAIsECZDxS5IAk40atjglLjHQVANgRN7ra7U1s77OUnI/nYuAYcYG8GV/GsM4DN6lIyH+an8a
OVEq/6mDAdIpw5q5Tvod0+Az73GmIQBp2E/JK5/JbWeqUEZ0ylXOVNvPa/JrB60RT8ugfeJON4Oz
nAUjMEGGRxNDTbj8VN2n7qa/FSMfQCUAdiDwwKn7BTRJlJwxP7b1CG5ITz6NIW1zeRsgF10/HvRT
JCQ9VQf6Vjd9R/8GfitQXzbLgv751N3OkBxgIfvLNd3UFUwBqJmd9wH46mLEDA78uqBOTTSmckhd
Y/tiyYl+1xC0XV8XjiAa23Oz0PDXcsaEn3MFJsx7GpxqGrfMKTXRamveOannRUx21xHhoENS1mOv
tmfmlOhvUYadcgx/FVLYFLvoocRIGYE2OpGw8u6dmdvYTgXbPkdPjGquvjLY+XoGXYot+t1CYcZd
eOTSGXDqnn1lA/kpbUnmSPQkAZ0F0ZNu5SyjXQ/VZIGs00KIwojBPUVx481E9UfuSwmSFnFXzNmE
u+rCQ6PmUmhKPx8NgW/zoy6TuHtfSSLyp3r0f495V0U5ILpW+MVjparvEfu6uP2A6bFx72P+avYp
+I1WZ+RHFvidHh6a9z22F7yXOpwINHs4BG8QKSaXZapszXuVc3oxy0oLSxKMXAFX2Q6RpO4B0EFT
Dz42wumeT4hpWfdsLWQPdeCMS+2N17kqp3TjT9XAwHTvWznOMu39/bS7XdOrMYqxlNyJJLwrspjb
q+Nzka5VoqNricuTgqa4mk3uRz433uD/a+5Ml3e18flBIDk7oHse+981cCWAhGUlDRP0i/TvKqUm
riz5p3j7Se0tD90O7YioAabpgecnbyHI9AuIkMp8ED+OXc1sFzDeckZKmPDpbwmiau7yrfR1ThCh
av75G0v9nGVh3i/oAEml+a8bK5+qqNXd+h3ekhm+GelcnkxMjiZsgdNg+2JCnmsBJZMvESuzQUKy
R3/wknyETienR0e+xbOy2ifdbd639CJn78bQX21PSuh8fPxddmRAa0UMmLJ+C34+tbzb87phwV3e
aFewqJhbKhA1mbJmc6UbWw77aUve16p0Yk3LaeY6MLFdCYU8yiufAJKnJTqqWsf7cVndvsTPsB9P
l+/QCOQ6NgXZNcGlu5I5gk+gTtA+4W4lIkC7Yvt//bruYmNpEryJrLKtzwqylbvFycGZ+Mcw7y5A
TXSJ0MgSz5OKlH2nIP07g0fhSwPhk34vh5Oakz0Tf0oJpgt1QzzPbm+Mk9nkLW0gVvPlK6NRYrym
QwJPq+wuNYVLVjzUTlWvpqa0n2pVXHGDwZ6EYI8lCYHoVNv4wMyXGR6eHmShqeIbLykuzhnZaG0V
JSjFLQ1N3eW/KIuXQqKV80JRiu1moD3W7BKHNidTVXt5izUSWhHUFv+Uz5U8td8dVO5HT+yIp8au
g3Z0FMzEVFNk9s5ySr4xPvijeViJTEm+NntVsLgFKgqvAcdVmuAFpSLIlP/jF2/Cz4LU3dKw42r3
vI4IACWP5VwS3nuqapluGKE7DlkpfF0GF4d72onTW71kBOabUH2xMUc+W41QtzRdxO9OZxJR9oiv
OHPdLkqNGnjjZxppU6d3h5Lz2UKrr5X6IlW8q7D/RCloyXpwPVPd58+BEqHBOfRh4DC5+MgXe9RY
+AGPZZeYXafUfR7zDDJBu2wQ/S73w+C3IfDdHRTNbYW092+VewUNjcjatgHI9qXrsmTTRcRkQEfY
Ccdh3cauhSzeVM2CIjF1kqPmA4VGz7vJ4C2IMFQ+n0BUGKEmi/vqoZGrfd2zdSZ+xMfbt33xMNcU
Yt9oZsrpX4CJ4lYm1LDqVxgf45dV3WIoaM59479I2XcM/ZwXCFkhxVTYlCb2SOioT+NkFBSLFkbz
8ZPhOi/rGZauiIH2FXqIKxmzNQOWpZpirGZNRQHe9j3gidJa/49XDXetKbxE2NmvNDvYNbynITWQ
+IUiUhWwqKMWtBbbigFoaqmtWPyExCVcRghMlY0mGSgR7zL0a5s0BnBu91nQ59uhvGzKXEZR89F3
8EUOHg9fFcTbYA6ATp0g2Cur6HAkFBWdmf9lk2iLdBpcZR0stWFj5YzQzm1FFBxgtatBYAeOSnTG
hZJVkQEtHexWJbDx9nzreaXf3EGpr68DQfpW7Ooe+EUQnQdbXsmPIMZPT4JdJEYYln3vjSsNwuE4
0FAhfoj/sdvqp/4Tygj7frVDGKisP32fxjkqhG3oG9PrPBerG4TU1kmoCWRzIKe5YMR7MyeF8EV7
KJpwypJjlqd12pFWfxAZV0fe9d7krymCbTVIAHRYX/msD4uqTu5f1MqeRhvh9UyU5qxhP+2YJASB
ZXrAugQUkKLXnWTDE5tYBZ+Wo5+eq2T53gd1MF8Ywj0+2SOP41/xwDWgf1N87uZWiNhwoMz1QAKs
3Eks1wcuA8GqnYXjxmsZGTQLYwKKp/mtAaWFFUqQ5s97ElSpltNuAk6B01zmoJG5XQnGgQlob3yj
iDUwJXQaBi9EiGMjXnz6zqpPEAfBvPe5xIh/lzeRjTvAjLdo+EQnnfugt9qaMNUgWDYtN8UHAUYK
Lt1tawFTw+GA8UC9uUu6kL0EVKHWzaA0DaB5HeQbk2lVKZa5RT5HadvICDkJrZodgnuNJFn1ZQVa
H034Dn+jRM1nA5K1xpTeXVaLSnxfyrOYraN4I21DPCdn5w6meG2UD4uwufNRFKTto/Hp8MKXjxSs
IdVXGHG+pexqvC3SJdUTHG0jwEOGzTaT1jef2RS6UFKqyQ+ioDjDqX8BFumL3Yt1/828ZMkrmjiU
+6Mtzakg/TzKn8B7LjJb2iKm4KmGUoK5AVcp+8R1rnXP5MkS0QOPYDgSPRxhb6Lc+lG74FLPixKt
uxaayl3zIvDmuIIWvEbUg9JC0hdGn6mGFBjAF17e1hreBIuid039HgSWAJMVUbLZkn/FyFEU5yBV
3C/YCYqdQNHHxSFRrUCr1q1518rawCaWAy3a35pwOdNLjjqIMjDv6m4P+mNh9HQcw5lvQJRzPKyw
8eL2dIIsyERyodsyI6tvI6FpBOEFVWvuctr0KHs9fyiUVa1oRaL5qD720Dubbv/dJ1joieW1ZTjI
tuKnWJ0iTz88Ug5s9H9Q9BUuQdh+saQphqCB+ob6EFwihKQeuLIO/W+xW9VCV+ac8SQrS1zgHXSt
oo7yhBeDxGOm1A+1eyGxKquim01ShP0Q06VnL5Wyhcv0Q7rIyh7t2Dybsn0kLNHIWiHYiuc2aC23
JLtP6G7jt3Dtbh7LTqBgkDu0mOLVKJDLBOH34g2Rgpxf9mRnNL5N5Yu71+atwFWCBNf3izy3zRsl
VQchQiiqkZCOmeHuy33VgdxA9CCO6D3S4lSo5sCPTgr245wi7OlJ+b5g/+9h4u68CONYmoVFXRLD
/SbqpXHmdphPI0fp+L963HIycvGYNdElpUD8enuBI9qC2G+yxKXfhscmTNgcB7q+9kY+IiDZKXir
MmZfXRYAFBMJKltS/QdZpFQdnOYDTHVfkrV2ItK2aVRnUfPxNAqGawFW87YK0nBgJmi8S/qh4Nri
2FmmceK3TxeSwW3s+sjZuUTeZHNbph3+viU9NwGEqGEdSixwcHapol7LJqTBCikoho4dSauM0sgF
Nswjjo9ExdE0Pl2a0ldxIgVyH57BnbtWQGqnbn9HgCgTi7O8pHxnAw5/+5S0y2p3LFFYynz69I2d
PYgtX7Gj/MIsv24RWlOKBf9HjCquzKuqFP9q+uvX5+1rduuDtq/eWzUaxXTukoBhUbE/uSjLtWq5
/0MwextmJoo1ChZppjQhEV+cA/U4VSQyabKkMnZ9CEhoTEcmLsP6R/T49mWz8bZDdy9xNBHnSQrm
5rFfkEBXjgQjEaUPPSnJTqMy7AGCqEHp//hXPNVtG6my+IVlb1S2wMhOekPL5efgB8hjAN0JBtLQ
loXMmgLFrrZs8XZ6K/lBLOQo38+tIGjDf/H2ckP8co7XseN2OHsJugnBtFm36r4DrvqjKPK+rar2
Gy54E9ayahxI+M47B19Th5O22mnqmecba8NoTIsgQNkVP3XtUr6RWqwU5ptWEBSOTB3K78s8OQ0/
pRuFFJZDYCeTSK2A0Hk7cNcmYa/kC8apURmzKqPDk4v4F6lD4/h74pXz8hgID3NpNLmtYGFHR96T
K7ztKISQLxFeup2g6BoxKQJzCV/RrESJq/5dK/6Fzc+9HB9zBNbe1zYRB1oaQ7kZCqkqChMg8wG1
J9hx5lSMXRebMT9TSQY/FsC3xSyKQt8j6jjp0BfiAAzEr5K25JTlm3JA0dkuOpOgWIINa2OBwUe0
S//gLzs/tGSFvfHfYhe6ysVXcBYIfa+hU0jiyW9keqMMjs+KUKmZSIYF8ctnhZICCTHr9dKGO8MH
oTF+qjJQDZ8QS1PEbvpztlF8a9ChE3vS7hqa2w1Q+WXHQtZK2t4iV01D7cdm9LzYlVxdQKjs5IE+
W2k9J13ZQ5LlvNqVPIDALx4hT7fgjMfRi4w3IqmUHWsLa4VvW6ZZRPLczjZ/XnhnhqCBC09oZHOd
tPlPy88b6JklmiR9I7CmUDRkgsrMvGU2j1zwWuReX2Yf7xBpeTJ9nXhXC58c2+ovu+kcgCi83Vty
B1bZmuvc1CuvyNMu8qYGMNd7PBdg6d+d9gh7EGzIInwptvhvuc0VvyXAHsC2BGj4EkxjoHIkgrpD
1OmlpNvk/1l49M1hdx220h1N+4TA9y2esHar3B0EnH10LdI2dfz4A/qkrBaAi9qwqYS5CBvmuKvB
D6g+28Aclz1N+HlWsBgcQycpa305YYTg53bj+jm/I+JevJ0jDbTZy1v8YKzEEOrm3pzYKEjnR+rz
13nKhqltfOJr6ay8WTF+Bl8RgSBuV2DpRqjQXnAQ/BE5fDO57pH8SCmKQoDtLc+Y1F22LtDLt6Yl
fZ/vAKbK/rbTCQczwrSmjypaRhCnM0NiSq3O7xd5J02mvQLgiPbGe6oaRIChOpk8XiV0VlOdjTqj
Pl/ToQN3Tf9gSgW9g0/bMhP6Im6lpiwemj6slO+z7BKnq1vTjMfpQY1rItN+9PVrN8l2Kl27kYpB
KPxZyLWiKwXXA3RZhAw2n8EYVhySe662VgVFTDtIQYBguEdLihReZ5nBp576f9QFqctxVEErSlFT
nKZstVMB1WXNdFCtn9fGOE/NrMNDQ6smnGGUKvFBySrd3gIDgsVp2/bPD836wTWeaf2i3U0/BDVA
WLllLm8RvpKgcfHtWJ+NhpJk+N720tTuSalOrWojzg8hdg4PgIZvG3Jsm6pgfKd/jKJTsE56o9LJ
oDvGKu53sXgPLxXN+kg17qAomS3j9atV0w6ArBHb7PlJdjMTC2MRhaMuYrzr8lqkIwaouRDjJH0H
IlGpQQlZ0t4AvOEpfH5ByAJK5S7jQftck7Q1q3q3VYF2qi45Gu0Zh/gZi/8fgsVWVzQvgiVrn7YN
+tmZRGu7alYFwO8ST12PYA/VbNuFXH9pxuSym5WyiYx88VclfESW8k/vZYJL3lQo5QHplE1R23vy
B+mdq/5rJv4VKjUEVcRkw0eWgsXniw0tbhSDqLG3F+fbXH/GlMCEmTtQG34buDgNtNLoTTiHH3UD
5B3Od3YkcpgubchrzswrvzTJkiUiv9xx7XK1VKxbQ0gW6Guyatjone/gsoJlRXUqlr3D2KlXAiXw
jGn3tcgriLw00L5btXMFCe7Ixr7HHjRr7Gke2XrlNmrqTyijP0oo9BW3sYOmBrvRXplT4lQtJ6Wl
Ehne5Eg/9JOijsFqk3L+9a7sThhlJ9GxGBU2e28DdrfYsGKIADjM3cMjNMpBrlP1wrqWHntn3NXF
7gBJd9Cj0jMtoQUKwi++tc10sFvYdqvGMHl2G3WsDxWSq8LK0imTKYJOfrqkDgDiAruC0J6uFZ4x
6FmFLXxjJ90+KNKVVwdGvVPXtbm63kjKH/ZKXjwy/9sWAygugT2wKcfOqutndiTQR2fcL+jmvvLt
JVCSswFQT3GQ3IQpYyRmsnjmMca+GNMGFP6g2c61Fopmpz9YXe8Olqq9+dKsp/EjsnF9ZtAIat1h
uHAAutE3fVRDaLG3Ag+0JWWn45lA5clRQB8qzajV2CsNnhirgG+JyUTSfhhxKkaIVi7pFyQLXUQc
CSfy0tY+y9dP5BEjVPezKWQJ6KsmjdJJwvJE5Zwn/sNmbDk2OyzbkdvVTA57OWnXUMrGsI37tbL/
WTub3BlOgIbmZMdgtoCCkYmMAcE6U9nUkGLdfIODS+lvVOGk/4zkZgr5ABE/gI1shZ4BS2mXVAZp
/ZTLYS3PQ6ouScXKFsaZwJnn81HwZ+tUbKGcvWfFtERv8PhFodIaU0IU74gBovM3hN7Uj2uOsK1W
J5wTP25q5vEIi3ckCIfi3GD2B1XCMk7dtnxYywTIOdfN4wNhDAuig0daEkVDUOGr2Lomksf2ZDMu
Zx5aWxSVIipq7jHQoxNfIth8KxlvVyy68T1uSIYfM2dsRy9KyZk1UrD1n6MSyjbnrX5Ab7fj0XpW
ZETENirIQRJ5G19JMWzF63bzA7GgKpQKUJ0aMOjQcrhm4lB/Iu67YvHCq6PtIvHrcMA8Q+ePCUbK
jZurt0PdKwckthy4c8XDOpZRLMcG+QFRUXrTCbDMeJrysfUbK2TdyuKnECwwN8SkT8t6tQyu335h
fDBP1YM9FVxpHnJrqLF0SjONxomjRKGZEP94BL39TcyWNBrS80+kEGBuulNEGfC0EJDnZpU7XqOw
7aqch1Gmze/Y+LC0CqGzPYrR1x5OwbekXpjm7U4V3H+W4H1UEr3k6hrAV7sHYbj+AGL2euhsweCX
lGUyjoTr/L6baZ/CRb9+t6Lc+szQlfEK+ZFsoIiZfLUuvP/Jb3UCR8daJNV5LFh54yvDvra1yZKg
XSSUULkh+0gwS1sG3JR6SXXMy6X7Wgln8VFROC1HAFEMBqv1Lp1W35dhgPIFLqYVgPT//0kCqbKT
3trrolsJuhnSSi1agHp3A1Xs2KNxDhcNdnIi1dNrNEjatEWIQ0T6PORCbTUAmme5A9dGhyL/AARQ
f9KoG9YAUIdZbdzaxjUu4iU5TXJSVhfQe0xZtp987Z0pwq2ZGJQ64mDwRPuZ1MADX7r0ymHye1TJ
KDYb+gkfyleUKbLO7xtiSaP8NhygAWJyXc9W6qCHFKbJA2szyOrIVmjNN/kth+qO1ruy6w5BWWyt
zQPLvkv8HhAUPl/JDR2L6q25XmdyAu7W8X9NRb6BMf9woT6rhQYHSSE3vxQhOr41sLZIDIXDp8nQ
Nd2qjn31VGu6x8t0gzPpvFz71SPHp0BQSaD4xkBSPbXADj924o0N45KelS00DLC06YkwTmE/ovu2
B6/cWvzGu22b2sJdx/npP9y2jZcukDKsTBe2KvZB55gH+1TuFOxpOEyczq9St8kLnyyQpypIXzD7
hDRlcQJBHPTox21MpyAmymwXDvxUwHNZVOCfXk2Dq3ewQMi7lB+Vi2JVHNDLn3uLa1go9+u72YJK
CBRYAommE0Bu2OfQhVepXBwjmnO1ydrTbjOaGFTZd8besibJDbqme1npcgsBQlIO3cGtkjvuOtQY
TADsdYCf26piqrNtisK/J67TQmUSQUAwxE6hH4+fufoEaPi1hrGLIm7mRflHws/8ET1AN6TvwPDd
dDiMByidIih69ZJh9jDYKNoy9408wM3cR5h2qmk3W3TCqjyCQIjEdm4uNcBRljZFE6PsNc4/RVGA
ZqqBxxPaeiUc+Yvk5yQE/cCIdS7DO8k6q+aEKc4IX2HSbqoLMnZPq9V3kThryTFjUr/JKBjz9BK8
AFETyTkVqgfLkZQPtsh19P29qnsTpUOHCBZOPC6QMjvhlRQDbsh7zSag7mkOJJUoTR+/5AJ2yUS1
9MSrnVywA7udaZ2WNfXQ17o5qsDzcdnZsRLgEnQU6o0EpV0NilITQIzDt6FTvo/JB9poiNXCmKcJ
apy+Z23wO6/k/sEuAjD7bP24ispyE+Bv1EKOI+Mpv/1yQJ91I9YSAJztNTXMgPl1FWvw7r/PK3Lc
Iny/LYGrfCbEartwe4PdHc4A6whU60+5XyraRG4ozaxreoIcWq/tZxwbHDzU9IOyhK3mBAJS+0+l
Qx7mk/RUZQ80D3et1gXH9vEK20IddGuHSg52bjVTLWMnYQsN3Xzy4MpRV8vHGrL5J6Spk4ka2g4k
nGPj4K5NnMhBFZsaI38qisnRj/MgTxuZ3t2cUKH0RORqE5nrt4jaJrIO9miMD2+AUVLFGH5pB4Ie
CvsW/cMKYBqPaYBNdjM2v/B7aCqyqhm9ElnwyzefyBQZSY5u6T1TtM3z/82pnhrNWFng2Hm39lWx
xIhkN4NKRm6loRdu0hj04ub2UNdaC+HgaIt3yki8XN+Pj96rn0YkO9wrN0bGn+EHcoWx1TxmYwO5
NstxvfZQ7QUVBRAU2aBUBUNBJ4ZPyHHxdqhK2KpigJj/G8AouUgii20vNSFQm0qcZCRmsmIEu2lD
zOhdFzRO29eiDEp6Th6wCbPcExodZ1eJ8e+BTY8wXp4AwehMsnMLeRrySET9e1OABXaczleJghoA
VH6MUQJjXoADH+siWG1Nn+diLmwCQiMM+zK+kHIBIK1omBOOjtvQL10YfIxNaQM2Ah6bitnZZggc
eZpYV1ATs/ljcia91xlV7XgtiSddK43Y/15llxTPjFfF8/rl7jQHjjR0n6QNptWSNpo5EsOrPI6f
i1lhuEVwIqVPaswqV0WZCDAhSQNlmjvgStPqrcQ4oF+hsFOJ709PwKOK2i5gNxrwwgTxWCI8kfHf
ZChhg3kYX4mZ15JyTVCLkh6VMiesOWe1K5ZdUYpGby29kMDKmO/BkvUrl8+fQa6rKsLeFXxIJLLE
X8Fsyf5Ye4td1fOc82Ilswj+eZYAEBuHJ9hYsm/c1Zz910z06xce1EbQUSXg3R8AxbhMpB+LW/th
MHbleT4KGIjj45ndYDb86XZVXcft6NLQV5zaoLG0Wygh3f0aOuNTRHh4wXKJ7Twjwfn7xH8TChZT
rf34Lb89QPbpIaaGa/7yN4BeapVq1XS4NoX+JtcO+17pjOXeEeVEo6sqdcxj92sf6DicrfYbaoVb
Hw0EXjRKRk6DhIm2FPU6DUHsJ1J5INd0HuAg3lKKvsDY2dRtzG0D7N1E+31M1/++CdLwoC24pNCP
EDkvEwBChxyziaVxNORdni/U7t0gu64/lWbLaVDLxblFsBxf8wFo/ZSL3wPWAB5Z7VjIqbJwAbzn
FDpRy52/Q+ZHQr0zuwEsW7bbujA4jXNOW6/oM4jaNpLc2NXpysSZ8Sjw3EDI2FXjGXuGbcqbpaV4
lUHcRw9o6JruYZDo43HN3WsI+znlY/6XpWE1ANOQq4C2h/uRuse8k5LbiiciOBtOd00NOfnBVwda
8Mf2dV7Kn0s6l9EaFK6bl6rTmEk39Mhl3+YSEFCEiGbKd/nKQ3UoCs2bPSwpSEZLYjK8a6rxJ4HJ
da5AuTXxzsJYimJk0cZZ4Ycia/2oCvs+1kz9Aae1j33DAgVl/nk3BGF/e/FWDKtaIOu2PJvgCtDW
wXVcWaCJP/0t99rvdFSlm3PBMJM527/pzyXEmuN9+gfqmIJyMqtSqYzKhvLH2A3MUDSmpjkUNGv4
GED0aD4cFIdPG6QvVm+uipbp6C+dUS9SmXUyKSVvl4FyqM4rdIM0Ri+4zudWbt42lAoiJ4SwJTiW
Rk6grJHfeR7K8S5ZdZVIalmMWUgRQ7gZaVGlvnqtM5F6Z5FDPOMi0UHMhPot/Xg11eykTc7BH44O
vo+T8EsWm2BKfgz8UKbVQDmjNv9Cf857M+xzqqqUQ6LILQVJl8G7QkYymhaocQmwkvSnh2KeF6l2
V4ZHn8hxz3aJjNTOwFRbc6MZrv/jb0lYFW3C1TBJ5LI63O/r7IHrKLGLoSrJYH6iS8E6dndmTr9t
JRIIOeuamIbnESAHMCQhGRLvIw91BEcjUS3FIV+9ERqdghEoNG44Hs5+0eLresuJKFtUx2c//I94
fUhJ0CS6ImUSxPNHh7FYBoboHIddbOOIpcfk6wOkFfNa+ZkRKhr7IrrvXndg1ztONQ2gJFIRQOJk
Y+QnY30psqMYjJtPIqNmo3+rMDvS7xX4X1OqzxCoFcNkynFj+laxvU4uQeS/+polhccgI9CV15VC
eu4rRVSPKiNlxdow2KNJdPjGuq68wTt+0OxqK27INPh26m3WU1BcQRptyd1i18apurARyAnB+RvH
5v8e5c9CnHi+kQRUULIZTnHGfi9/9etVTKT/RjoORhA7+EpCEVrpAwxz3x2VPJvS5dEcisefWgJ9
82BJsVBjrk1pgiFr+eu+9dSk29dMYaOHSDXgXxUY1opAlfeMxE0qJnO1BA7bq3UDhRq8C1wg1jZD
Jf8fjCn7tmHjWfwGY1yyaxufjrzYO+YgZtwDy2lo1lCD4bPhpT9U000sAilF+1r81X4tGHNYwlCp
XBE9AxMtrsmB8OtfQOmKle+WVaEmVFv8YD4bMh+XjWA0SJUnDf6QsYFchgS728Xa7nK/FbQ+QVmj
hHAjp3ALDq7AV1WX6OMFmrgud/AEiZQzyOnIWArJgXho0Dl1SDRAPOy2oO1qETMwQgTMFR2mbmZr
DhCQlJulmdorniU0LB9iOvdfg7/R82GECAFU54tiB2OdzqpT+7Fngoy36SwHTZh+uoYcxR/gHAt9
DlyTt7tyBoP4gsZSaovLYonLw8awJZnTRz/Y8B2piwPozxqmFfXa3O/5JjBUNXVOOL1+n8qDLRig
jaDxG7upjN1e8juqeovez0j9d8ydOn0l4mjTy/aWBvtdXJpUHOiPx9Q7tKvzoPh8WmoGW3AUkpEq
2JUNAOnslEKVHInFpo0R4m49hucmC3SWJH+3Meb794S6RToDLlk/A1wIUUllRSgSRcav1UVQWqib
00Krz2W1SImYUI1T6X7640Y9pgAtgfBGMs19xKlNtaNz5fNETeAtSESoE9UYvJUlaAM5ZZ2W3ntO
rL0D10PgzqXvix/Qz0KWaWid3OovMEwB23y0LU9KqrXS1s40YpJ/oZM9lr0rhuvefWgz86lQKVKl
A7dyuf3iPWlPqdXo2uK7eFsoBbef+zWhC7EBs1PknlN+41LgF6yxGL9e6H4/JvVTkMLFxyDHmmtr
908Owu6vk9JJVEXAjnmOiWwCw941CFhiZcRr0C9Pt8h26a5B7JFLfRGTb8J+GEPy4GYSszeZhdio
YkAx/FSX9lqW7rl3GDejmz8tITAGN4KKFnNZDlXfNaZ80gMNWbvnWoZEvRk7Mv4xSdD+q4YgJVT0
+HnwQ6oWiAVJrBzIij2PgXHSfSebZ3JFNEZARLBXP0dWilDRnJgI4969N8O+xdjP5q4cnGS37FIH
qP6e1MygkBfrZAytBfmM6ALc4uM8d/CAtSTMY2iBosyTYhcNrfduJVDDAfK574Yh+2JIavoUdg/1
PL1bmUDhtVAXVe5J+/Chw0ITXoTBi/fMMZLdYabkBzJC47wWH8jVjwIfDy/Rz6HT6cKNMFc1wvza
lSnYpGW7veFTgC0h7XVjglk/X+oAudpKhSvw/Xr+Z0g8eac3ZhyFFxPSnShCv5ZCh4PzBWax1V12
mt+oLsMXZre9cAglkWXTDkUmKTZUO99GoeCS3t5CJgvLtB9Nq59xLmpmjH+wkNrrkxKk/QKhwl9M
p8oLn3XAUxpQkFdWTE3iVkPGBcDkhTioeNAH2gIJPF0h1W4t4WLuYuhRqJeoQZ8xv6jkwbIhZHcP
eV0BBWYVdzFjFWLcLgeVkPnB0+29RlsMk9zzUxrQgZ0rWaWQgc3NVONvOuEMgafGDB1Eef60D8a7
fGhgxcRooJbZbl5zlfVc+tvjv/IHUxEpulYNb0lp1UzM+P4rQ/xk/kNTbqeUkrW2JxdPNzZQZVxT
pPOxXyDtJXCdVd57nEfwZIEq5gs/sKksLK0mbMVMCxQyZEKXOArrAyvMV/iNZYYsWpmERjOw42im
5yrfUCzd8784/mz8gbLPNiM0yEHSRx3/XO9L+mfq+AnOGhRqRvXKWv8FvXS24pieNRu+oiJI1gTk
sdvEAcA/rNrNGlqmRE/9IVnjsTeiGubEm2hMwBAaVn5pRzCV39G/aReeY/5EKVWzbE5NIxOT2Ykb
ZFHxlw2NBvNuHJcooeoady5eaaaYzVxDDu8nU6Yj1FCmVqHqtvrFZ54EZWkrVUj0YxkzxeWiirbz
l6PaWLZ8armdfA562fowBPiy4iLfG6AlvmaYjH9xg7f+vDCP6MIfEn2aHteHfCOVm7CQa+yp9EX8
A7xtB1x8UEkk5QyAnpqcUuc+VdlmKHSkflVgJm6T52iT+1wKTwI5sI9O0W3xJ50XDxgLKniV7w3D
ZgV/r5HLuFZ4/EAl4ktwDj86Jgkg25Cl+Bz+SiABFx6l2MMLg19Sn9/vxofm0lH3oW83Hxoqstom
LEvULMZNpsw7oUwbdNlObtMKLPeK6cFqPfFVH72q16PgLWDkpXpAebnAwyzjwnAPqChDwBd/ANQE
ft/Tzn4qCAO/UkAbxyecpThjsSEAYc5/3B43WWAQ4I61TdbaCmeQ43iTiK2S9Og+JDn/bmFiHHMf
XtXomj2SUaR57U312PVK2aQY+R1PchwiL0NEPRfQHUr4E2rqfP0ruUsfoRaVWlzjGAztTyV+2Nfh
rkBn6IlQJA8rgRiPFQLXQhVc3QQHAGpH5zc2CuEpqwio73E9Y5+h91w6wVkgkOunQ1n7fioTEiMO
vGiQuejc9hcWVVFnvpautwfqAmLvelp5ruWpOcbFp516FTS9BRPK9gCXD5bV3T74wZwtVc70I9j0
2/KY48+dpJRdsEobe+nPLkFif9eTgqyurepkhKlxcy9QBY4USd+Aj3PAEV66My9NieTRQwb80efH
gn/Af9nKltqXmHGteTNKlGqhsEsvIt2e40kVaL8LFWwlBDQr+oI3Vk1n5Cp9k9QtixcgsKmkaXWR
oqQIbknNvo9+c5r0cuqPZpQd3sOSQ6W6lxKe4JWFHLXBl00LFr7VV0GjeQtK5+6hxwm9g/JablK4
/79ZfbU1+qfh38l5bfbYXROpaULyTNrtkcZgyeaHmr96UHLveP18TQ9em2xwJeJDKwqzFA8RFAxC
E0wOQFVp5jj0S/v3OTdVDzzL4eY8CaQFXo1G7EzzP8wVRkAGOXs/z72Nh7G8UDkA+Jt8UyrtH5T8
/jEDe/pdZnZPqXD77jglikQNwRbnEupGEa3fOOg0MX96Y9Qc5xT2vnnw0fve5iHarfWi19utj13S
HLP0RwM/Llf/RbegkmSLbMvZsT10ti8JzXFJKAhqCjdDUAFlo1z87akSS68hcPkEzV6qNWhwZLtp
3wPl1yKXouQE92f5OR+EhbaH6je+yp6QhxC58PTCy2C4QwTwjcY4gKBGRgBq1dETiQGYRi2pu2uz
CbHX1PtgbS5CIzwhGxX88QVrZr75HKWqEcXBMncL6wP9dVRIFUeFNxq1QttyfkT1dV8eoM/lJiBG
wnJa6LIzhyEeLxFFbio0WpTQ1ej5ZXU+1hoAyAw6DT1uruE/TUW9hMEl80JJFo7+gQ3//bGijkkt
DvGn++JEKydChFmbwutszvtEWUC+MUSgii8m67zfpzCVMJb1pvvyfAQBBZyyzAcsosDiAPz1s+kq
gJ6RrxT1EqqvGc4TSMrU0VmIrJtrvgbV2wT56oOEqF0+F8s4wRez3TKTjR2Pd8fCvzohsASigCUJ
jPjqHITI4V6QIdNgfMJ1yIEqJnLtpwyHy3jpjYVmcpo1Io4pSUYIPCIDrZ5v70K69WI/+gpg9eyg
3D3cqtNOiJhOm+JVaFwgWw75/bBgPq6E5gbdLCmEGWvhPUzFAPY/v56/qN1IaQ7sQLy6Vvo6I6lr
KrqjRwj5EN5KCAfMuEoThbDkn0w8pcEcai2VotslL3Pu9p9I9at1c+pfLuc0N0fRJ7TCTdOJOXxY
DNQ2ooTnDvbFMYrOY1Vlh3HLmOuSx+0S8t2sAH7Rn9JBB+Qysgx576qtdw9pJzFFGwoG0ZFeTdmD
kj5pG96vKBigm7lSRQ69FCTbxFi/S6D/JwhvIcu4vy0WD5SqBp+usYPCvE6DQBkjUQ3zr3dw7Lda
0MfAPzVFA+9j8QcX3vzG+iUotg8J6A38r2TLmuZXRzefbdH+Q7nC6itE5umbkcxI1JLmdi0jbTlm
BzOIGAFKzsqnC3lTsBszRgDnsA835/2QhowT9JHN0s0XBqiXV2jHBZowLnk3JRJFCcGzNvJ298gD
MOZt/pbsrQcFyKoxkk9cSAbrOBEyC6iZGXWTU4b+x7xRzMR92EilxOvt666GKkS/2/UKFfuVLj9M
0+0Zx7tulbNJKOwX18J3n6imM+zWih8HiONBi2esSvN0OXKUb1JVD3F5t9ppL8UQbHiVzj0Wjv5p
rwYrQebXfzaRMp36mv1tf9UyqIzcVby99yIOELoPw3KC/bw+vu6Dk4hqYbrHHrQO2/RRy2wIxEDS
lCY45mJFUDT2U+KeUG8PKtvsJkUuQEBvoTGVRwtpxAeMmQKoZ3DjsZSTcrbcRLVidanbksMRpHHq
cTtLalKeP6P86EFdrY+4+vdqVMoRB3sRU89JlVDBR+xMDRa1Zqix/w8K8GAj4iJ+33jHzLqdr4nT
3HHapXurM5sjMIdpXN/DnVTi/UU/yKrHMbhyj9qdaBj+VnwP3cUdS5VoPcXLsEGLUG+pltFArhuz
JLqF2BiQB8XnNbATuJlTgzoWbKt5MONxXMNWR12TIinSRilzgj+AIvug0hTd/E4jG2r1/gRD/C+E
MA26Dut+NA7obyHZI3tapTvB8JGSkj/xqT4U8E3KuwYdZapLw9NUwNWF0UTVwg5+riybmBKQxeYH
Tws2gJG33hfSMAZOVikuyrC21PrZPAIz/ahSn2aqwV3C0ms7tZjWuy4SvghT4cN2DpqSVAo+YN1b
P9tgBRj5T0D7GYQWYtX+ZfI3Atoorm6NZWyxUyhRrg8RNJeDViWxCj+JWrZjdMcv0y+Rz3a2jBY/
mH92kJZkTvZtj2zbWM+tUREILpNwNNRDG0GNLb2wVCkyddr9KvtbA7bPsT5GPAYgL9k6O5f9L5H6
4MfiTVkIZ1d4+E0Fma7iJ/yBCc6nc1OqfML8sSDhAgF+6eNiYbQ6K2Xr8kHHAGWoDZXC9vznvkWH
z/7DdVnh3aiGVSYlgq6zBI4+NKiiNOuhGtnMQ2NUJA8dICmbzOgvBf07WxZ8HXqhlHyUXRQWUWxp
eKKshbJcJCK7FU/Dw+7H55BM4IuFY6ChQ4z8RQizYdJdiGDoEz0JcoUWLf8T5VIPw25E4Uk73//5
Kpq5iHopFjwyrw8X/lNqdtHtkCEZpR8k1rQ/KSxPy/HcHel11kjxsC14QcJJ8zHq/9Vre9sNe3A+
b9ZioqIXNx099K9TvHTcuEoJIcHTCivx4Wfo7qhMV+3YRs1iZXrvQ9z+KEXpBWb2zkXDRRiSQr0X
Bz7oNty4jezYZmXEPXNXC8+FHm4EoatkWdPorp9bxkh6waV8/scP+F5eajGA1jRge1p6ErMU5f0B
ITDWY22lSwkqLnSlcx/J9/ynFrbpQhyDBJ8U+HRXsqgUWUh8oORPw6a1kJRBvwxM2FKP0wgMUZ2/
6nTKmEpnJ9ko0JC099n9oQKmbNltxZ8TS6cIm+j+bcAjQQ8fsj6RMypTqxZqtgo/rjTXznEZXqea
dwfdsMuL5bQOlVYpm4uK6vhai39MkR9G9aXFURht6SpVmI5ZW7FRDmJt+sW98ALtddcW3A2SQUpv
5gW9ACZSRpjJDrVO1tE2mMwsQIyNtx1UJm6Px8K2zsNaT6+xk83pyagutD24nMt3/h6mqRp3Ybtp
eT5iPY0W7Kr2BTp71wjCa0/gYXaLQii5h7g6yQdBCE4WS/3q8ynZHDbfXgoNErGqEds75NVgJaUj
VeO2KB5yz8C/hn+0Yp2n9W3UuRaEtimZ5LeTfYMv+R4UUdTXN+ugujAs9LMHeGhqb6vb59RPBhN9
Iqt30f5G/u7akSISvSBI7ZWnHlf8JbQiuYjN62asxRwPwHsmduU6468zmdW1WFO0nnd1zl0OPR/U
yW5p6v+k/pKp2yOLtoVAmkBWXd2egoSufxOZZIbsbpa8W6t+7b/oxVMDqXAB76j6bsWTRNdUVyj5
rABDUkdsRJ/wfbOcaWYWEuXlQ3zm9cT10xQnzil+u+dYYCuEKlRJK4xPLaE716rRIraxPy3CaHfD
p9Lkmg6P+VaK6u8F6KfojL7xTtI6CL2DvQEB7uPotFnrrrZd3KLIwvrbWlk/JaKjypz8LWZ6BfE/
wvqZy85+jxweWCLcqE6tasBp3JVrxM4Sx6r7DOjNOlWMthtNoQfuPSGhtGveTk2Z/DcmNK9cenXk
N17kA01EIsrFQGkbonM2w9XyoE4GJBddIgOuHJ6ATfZrZcHXeTiMC+gFPinshiRmsbIDLq3u9eQu
hmDzfPbpHivjlzTy9uHzuij6It4gj0R2dB1pRAIYE+CPn3OBC8iJKCoC6lAuZPIVWgYAAL2v0eQc
T3BP1fSBCJ/7t8HruP0wLVlg1W6ZrTRneI8Yw9vem8y/XUfoBYgCf/vmg6Z1SSPtnoBny4bUXOfh
X//VxXwCkKF6Zv9aWI+kzWDvytRuVEm7cOCGIetbIASJ84FuAqWUiC1Ew2SLUhKtg+Dk9PbYVbNx
4zdSo3mkJjxvIm7CLiKNIz+q3PA4Nvq4vzE8F2UxJqQQwkifnunr1cO/N+0RHfUQJ1FE2Fzu4RPg
k9cbnsG/RqLME1kr/b0h3cK0wZBAHyRrvueaMFc3tA6pJhCPvV2Vlnx+Rs3ygge9tQCoKBIP7chP
aAncfbQIwNASSrdW4DeA+pGbw2QZNH3Twn0L16SlELDTJsr0317DKstcFBtuSpvrVWM9NmgbMsdM
bR7hxhD0syH26vpIrKSdd3NazKmZ0V9ZxPXpTixkbg67dqhGbNuVqNB4BxvJU6a+FkkdgtsZJfES
2ghB41Ohe3P7KT/vPAaHWe961LAVS6LtE8PfCdKHA3FUXic5O9ZTE0fDE9vfZGwRtGjvNGXp+tb8
G333byyIkJy8e0tlffSgol9MVIOk/f6uZvo1RIzac13nmWVDUMNrAWNY8Cy0zLqly9uDnAAxkLt6
ZihxSsVXjRG3FY0x3LKrPmI2ZgNNS2Gb0PW3gOBRkx0XgooysF1QAbkjK5ZC5z9HhYGKQSDoNdkX
LDTGi9tN8tRowPIjJ+UnQ3wq4eJrAH/AHZS53CEe4RU6/MtcCLADfNEUv7jbnVzJTEPG0+1FaUEA
NxUJ+txdBBD/7Gf91Rbx4IMqIUm66Xv+nihGWv8kFwI6/Da8etDN+y58YXGireOIfHJidEgYwR6S
Su6t4rPFSRMeXRphxKGWBt3Ez786LTeM0dz8SsKW9ZVa+Bwwm5tEpOwWlCBOcnLfDYVBzpk3GI6x
Xv+6mytT7eliip0bLil3G1IWASsl2cr/ettx5f8K5WRL7gZM/Tg5LdNdG6sgVKrqnJqIZBt2GN6E
TfsrpZYF5C9NtBEjZ0JB6D7CY57manc2CD3o5EzHdY0Wf4FWWKBlQk/ZRUIpXqRvDrrdaP1uhcA8
B/Si/yLo+VoEEVqqa+rwsZ8KY4fcLB0cTV5Sts1TSGFp1Y2ZyFIqQBv0uIpoXaezQxuDNXys95dx
7RlteGMCAueQK5OHNoJ9VNUYm5mqENGccXCLQuu2jwexnvmyIEPS7U6S0ZcXTUNbCzVUOgFBarM0
6OG9zUFOVCfQISuhuIxmZ1m1nZ+l6Jdk7dgP65ZlGoaenEDf8ORcT6Th6pujGPAeOXtGqdxDkH7G
gwonIgXKun8jn1THa4l50OFgsGQRo5vZk5UmZgfuOw8pLOZPtlrag95Qp0sJ5p4ZsBmqWSdyUIZt
Ni/HN7wBY97O9SauWTREoX+4JB8QjlVAM2+JOi/auzyqul2iN9VQcREYyU4360NKn66hBperj4Lo
DLASD2jlariZJ3honvy7a2qMSn7joiGRMTz67BELccxLILo4K0Db2qws6jENxxmIPQFjV6PBKWff
NSPh3kguro7y/h37kuQq4/fNErMCTN0dXmIO1YxwZBJhGcoXbhiQw5/8iXCg5vMFPW/gt/7oaYS8
6BsUMSpQIxdAffxoxECm00WLAhlm77TvzwJldZAey7h+Ouz5dowO+EUyvW3C8PIYFP3dprjxUoMr
LkjETNd4FJuKyEAYfCFXxMwfQzduS3hA0GzLccoKUpt/M7xU4pddhnPF/BrhFFdQt6fV0TVLOphS
ydT44jHUnDFuKxBcI7rOBuD1OoFYXZM2m7yl9fmPKZVmSKx97AiTBRU38Lo0NOrtLcLdp/Bh0Y7a
MOywDV4uN0vvkaXZU79EQP/2zd4fG2Zu3LnLRmORiyDSZWboTxkI9OIe/GGCWa8xiV3iiVSlJjw0
7yFXBvTGg1u5XvgPWTodBN6ElqzyyvV2jDOhl1v6UXIS0PC7bERoVq2dk/JueAYweDhIct94Uv9y
qjNbcb5PICV0TkWjsiFEw54ffGLmg3f8Yni46HFoY9tFYK6CPHbekn32RaFjwIKJoEnU8Buyp69J
Qq6CofvZmOQ2sPe5XGb+6C7y6ZpRTiZdBaeXaswBIHcDPtJgMs+XSotjuKzUTSCOZPFrKfwiX1o2
6CIoMyves7029qR6XuZTayQVP7Ag6acPJ/dMlrDz8CTTfn2ejkCgKATsMKRvpEEC2vs40qiEj7ZB
bYtFWfd7GuebSyRFjCBNC7uv71Gne4d/dMrSw91eemelQVdaj3RUm/CmzBjjKF9dIO/dPntMM7r1
X0c76RMgslijQY2ato1MqG5z/BuJ+QWPNXaI6L5ae8koI7UrC+4WDW82XTWSzmbcfLsh8wOSp75N
KIGux5Ouj0gX1ClkN094ytxZ+WwVyPW7OfeRT9FPfuCRqSl2oN/5FnXO6N4EWtVqp0smOV0rPzEY
NAUcBfi54XkwdNYuFlg/fx+GvYCQBgTb3Dt7PbULPgLc0oqbnCx46oWoO+zRQEcx48wMUmxZCrWZ
neM5A8jLOwJXMA4Y1/B3hLbDyMe+/iEjZDRCOIwBt8ZSg6x6ji94QrMHmYNyLLWJuJuFwQlxkQam
rclQ+cFi2nXfxsrwCnZZ1jTpokNTeDo+/1h1fufdjqIkyT83PsSVvrZ8D2iXozvih9sH1mOMc3YD
P85CXyKJHp4Bckea7aXrkVwRRkvMsiYLTsV8uNuI4yY5ma0Mhyk2OQ4crzSO4lX1bCEnFz9KTDNO
d26lFXb4mkBwvwD0lB1vPxqeTDse6Hi7poaXPvJQlRSZi6bvnPYsZVLES550pFUBjadnAdxlu5QY
TnjZU3nstLUnfR4B+DiGFlTWgIT+LSXgV9fmIf43dzO0XlLaPQAXdju4JAyGmu5KvtiKphYeLx+i
d3AHkPGyT6ycJvFLZA6dJsrlC3Np53qs1hfWlxUg7dixF0BuP7Fphrd2fBQ9Bp60aTwjeSMK0PYA
rgXJcRQiokCBca1ZMpyZ//p6V2Mw66Get/oGK84XOQKjlGqByB277SzNr5ZF2jT/zE6T0ocF3JXh
6hK3CB0XQmmZXmlPjlWMJ8BlTHrWPC1+rmdmj0TexM9ye+oMtUJbf1UohBBc8vVXVG7blzO96i4C
xEWxap815YSbvkBfats36IFb6uQ3BwQj+/Gt8+7PWHk+V14d0bCpFrC95i/rxb1p2fe7tWD2sPJh
pQnoaa5btlVXhTqhj60Buc2EHvnCPQve3dYF+6neviTBl0QdkmkzKOUWjR5TztNb50M9JRbm5cqV
c9DsAVr21U8jm4Flut6TLK3Llzbz/DimVfz+rIwLTf4sZ+Yl0JDBiPT32QFtRbnvH1JYgqpc8RZJ
BsDlo2KFFXWQyWZe12b7LTwJmbmqn/GmI/ZG+uKY0yrAXe27jNtRpWIW86cFrN4O8+8k8Be4IJDf
tAMf1kMlsVEFkDKD2nWFdWcEzNaHBagXGq7Ysu5ytCcWpWEHL8dtWplIui/o+SBfV3lG2x0nG/A+
Kuj5wRSA51wjj4zrooGatO/JAMcvAfBUf08jIKevJ93kxnbvo1Ws7zgGw7kgVLsK3J/Ced9azrDj
KKBGRowMKChdeq4G0u4cPjmjrQSoiN0U0kJizqivbfbr74ZgVgmMxHV9Oclsmy4+lw3yyhgoRfZZ
ZZ7LYsi9+DpCf71t1j1FjNRTZYHV8BdrEaw6RAVc06tK5GV433Ar7LNrJdR33qNNDGZW3PwYt+Af
zOeg3JsaNcf8yt+oyelJWd8So0cUxxFG0aDJ1uK4CCpZqkxIZ5ARxuvwJ81gb7uFiLD92KcDZKqt
C9H7pcBSOWF95kjHWoObSZ52IoBCQedoUFy0eAX8qc0bAbW5luTwiy/UsH96nCkplfm5UglXcsuo
rmRSjqQxUkqyP57BjEooZpWLz8Yf7P/OuRotrxDXCeUufLkvhxOKLjqfRr7iAkCo69wZRTI8WMeU
rbC1sX4aplsHolJSgbRBnXPOo7KEnhvxEFcuhgOf9zOnpSBK7cy5TVtbh6pxUaG5ITLkg2ZaQOb7
rdQ+f785cby2uPKS3wowPq8+uexr5NbcpKfkXyenoF1i8nDcr97BvZkVP4QN/g0Xhkt1kLVSar/z
pgHVLQ0fJN9QIbwaqObe3OSrhn1BUNtInCRpAArDe6t9c0Lrk3zxGB6HApuVw730Hj8QkZKjIdVX
fnE8jbtT060xIDzBZ5hw22z2nkjVInTtEaJbgl7k4jpJbptwmxte6fcohvZBx3VgYbCCPpS0tWpK
TatS+xpRNanLMXDWoP9rDD7TCGYnYImfWVJA0H3KuRG1QbBl+eiglq5SbiWqaHi6qCzTYefv1XWJ
FzK5beU92ZfvXozoNn6NjOuCyNvfFum34Giw/AjkuLJXuoojnsDBd/5kzQG6y9fhch41sosfSe/c
k1YGiM2N6+9a1f07TeE07REyTbXqRUjYVzaQoKHxoDxDDrw2Dh11YKJuGB1PmHrhMTm/HLa1Qwog
mu30BdpD4lnYSNbDBXzD6k5JqDCqNUc3fcPGL0tvdWvsGbtYB3QgfmCOs1Dly93KTkGWk20x2ob4
eZHZSQgABKs7OhtFRvtBfEKgBiUKt+XxudPZFCRO3pKaAaOgNEgJLhu8mHRzj0p3rRiPZSNDm0mZ
VK1nwdPZ+gjlvQtvsP0SXucZck/WTZeNmQJyMwMGNWSYvhMTxxbTFQrFGXpv76i/k8KZx/1G5960
ZUZH5au53+oId+fNSL4FbvD1jNut90Ldt7Nidt/t2dUKwt/KUWq+y9rfXr1lVZhwNqpyd0Ynwwly
o92Rt5mY5uJMrn+fTzEjMrEzoQ/7t3FDPv7lX0W1DjD4mOdsShvVEmDqs8r8UGJBSKBtSqj+XrXO
T4v7KS4W1S3agHi8iY4U/2OmPELBEUCPXBVp7CpquGWb8d/JJQIVq9aXgxY+UrVoqsNhx0GdXmvM
vu2MN67+ZaOWjMJ4crp65DQgZTeapJlwmaNazjl6eulxJGjx5QWNkvn+hUFrihYBJjO22/uhq6jr
xJBL/O3QeMvCVsl6JNECKIqY/1MvlOxPDk5IMtzgzZhBlHJqzLkWuW10FdNrDKCiqEX/eUGOpTrP
Wl2cUp6mPLWsCrkvvrLucfNhulU1kQbfph9CfwH40ESB8x9rKd75DBlv6YnUz+KETVHsgTFZspKI
zHtoz4zl5cYFnIz260LzsKtb+3wtfSdB56MnlzeoL77UP1DvpL/bRxWMUvkJmyqfd5UeRM3FKAmm
NdUuWHB/MBnyCWt2HIb7fL3ZIsUxW5mAxLuq+VUNgibnVhtMS5XIBoht9hcK7C7CzvYKJGf1jnTF
XjeMUhGNUI4sYsyko6tKPc46gjaYLYFPGwVU8q0bAXVzrsveaIqu7Jge3fDuNprKQqV1U9ohB4AZ
xIibJOjNqUBjwBKj+FsLCwbQS/nHy/NtaUhyTliUh1HxTAZ6bwWflHFnuYmEbaeRPb2PO6ggmaS1
SFqJDY+kBCJ6WAtOnLp7nNseZ4YKHo0wioiNm7Ya0f6JAEChEnHWc2GgyNP7pB0Hg6jww0E01eoB
UDKCbSBUpu0QZarm9hWmyB90alCLRZaulk8Go27N8WED3w5t3srsclT2fdRU9wN8TUg6e6I/SBYQ
m5k5MHYosytdvzUQfGiWgb/tSgQRWm9s3ltu0Wb/FlkhdfNywfKKfNLZxEcN5iu3bCizgmAe+mi7
ESYU5CKkT5f2zsyYaBmgvaJjakB9M/3cgckiUvtapJpodzIfxHGoCh2/4i6ApxBPg2Ttu9ltNP3z
LWRaENy5vjLY9zbiVFRAUeuYVATutJswZR+goIcjUbozowzO7zkLyOtmmFmgVLl9PdkY4HI5uA5J
sMTz1Sx/wcixKnzLhVCGk0rYvDE8J3K/1+BpcGyzcql87i6u1mSu4Ywxsf+Bk9B0AYGZZ9O5j4I8
fUiOngpIAnyBzlZU6epthdKV6fe+AVaTeU4VcIm1m0CG2RPCK2X7TVXRIkuhKiQMALs13AMDZTTb
+0vreUv9fsutogpOqgi0wpjqHrdeZYdzZ2TjT8JmfCYSamtANxhxIXFKqL74MWui3zNBixo0oXbE
+2VYXe5kdIl+7nv2u7itye9RoilPQWG88ZzkhzmLMRAKBtZ56IPPbn17849pVHGEiqzM/NqzZn1z
AnmPJbpuoD6NZx5AB9wbzhNab9tt4CPgTOwPkRTAH8VP+D309W0h1FcUPoGSGiTGGA7fz0kWMCZD
L2vYA2FBzbujZt4Qoh9ZOBGZx72YsYnI3sDs6b2ORpAW+8TINIXINUmv0UY/tiQORnXEVAV+LfXW
wyELHca5VUq/2rbwa1w+G6yzRvif+Kwu7bw9N2Mzb7cWXOaic1QFXl/NM5yadL8p/FDbUZZwvOvc
M1M99TLh7rxxBzymY7ox5HHbzDElupDkPDB9cyblJDLnuQ8pBVn2Ubb49CrYJALtk6V6Q/XiskNW
Bw2LlJTfOLvxbR4yULJChQzSwkhlGssvN6KZhkb1/XUZ7fJ7Mq3IzFG9QfIQI7nSLDPb+fMGuIEF
UjyxJliEQi3mQb1WVhVvoI6DWpuYZ6N8lk8Mmkc/AqHS/CbG+fUaC/fdC6H60zJgyPOPm+w34LE5
Skz+lYx5M3RmwPnEvEEcBGtvpcheKB9Zmnb2E4i0yWK4FRIrJPXHOGp6AM8hjziN/P38QBOVYCYI
Y8wksedI0gwrWtFDeHlNtmE0Zi5D39KOcJzTRfHLafo/+7u/qf5jtPJ/R5U1C8E6TcnGvPGk0HnK
SYTwyOWlmeYfpbkkEjexbtDXWi6nBp6RFaI7Bkv4XAwaJJGJ1Ty91XK4PXdTywgYnHLkdWboWZT6
nVHChpOTdzI1UQXR4YvCBHXQKNKr4WZ/xsoakSeNj559h6ugpouM1/Y2QqAV5a+xQS0NKde81qta
Q0aVdULCdKiz6/WAFcMj6/nZoeuNRa8SCzIg2H8D1ZI3lMRIyjidUD6UPbqYEK4ilZjfDm/lSvxh
VT+zvR459aZhdCxYFvmHwNkkIY+mM3AfjeFi8huP9qkcbAMJIpdummhmN4uGjNvGiL1+u48rQKfx
xo5RfZ+mUCzkzA/t/y2PwnDVhvKHSzpg/904wuQMGRmTfvOcou6R5vVHcmkzrs9HPwxryXC0Wolw
924YAAcG1zy9nJGhWYnwzU+iAjQyauyLSnrPJ4sBuRW1FuF150GVDJ8fo6Xy4XFu7Uam0h6V9WnW
iG26npEsYf3BCbqQcXN9MALkCXWNO9iM8brBY0xt6t9YPLUxgK1HJ8ljJ9WtiHkv9dkRCR4aefFj
4iWNidzPLvO0koQMbsiWAzShL1qFgDHLU90DQm75sdh0rWL6D4p0VSUnbQALlchSZNthx7dzXePU
7Tbli3uAObL4wVdLrDHq4bxYqUaGVWsqhmlyZ+DsI6aiCfwyw/82INFW7TQtUQySAIWY7kOzukuJ
WRDl5gtHUu07+JlApY0GOvjlFiIaotTqBY80JkcQl8HrLM4idQ1FiD591UnFshdOuwOusSfyoeou
mTheRj5eSpBtl7TEU0gmwPG+Crc576kJvRLE5ymM5yNsZjLz64tw1DcmicH92dS8zq8TubF4gE+s
HVLHockmB+Iscgem4T/QZBzdKvh3q0zsobP6U9NQnxPHs0s7IsNKtKJhELF7X+Bj3zV0s4F6bQ16
mLCVU77+K1utTt+PMbCDwxlYdYm/1+rG6ET/JV5H+9Wl8rDUOcMdHbZF1H3emFAjY/aoTzBzO/SF
N3y3+sXHUca0HcYaHaiZA++Y+QGkGRzqs9KYj82FIGDkoqMNovNzb71fL6kdAU3Vpl8UPNHxsvUm
T9EbQBYLLBCp8gV84O4ZQ47+R6d9P7ZbkQYk6UVnY2FQSLvyb9t2riEyih2nnBso3LMjLYZUqgJ8
C/AVcRGbPMWnY4JfQtWAOvZhc78gPlRi9jUuKCYwG31w2stRkJwplTu0DMKQgQT02mzEIvJJSy77
2cG2eAa6z0AmSflWlNkpndHaSOTxtvG0BORN4HenA1e8pU8m9HsN0azbiPw9ZIJ9ECoW0oqijs11
pr5vlksq185xFNEnLUNtWVRcSPctAPEamqSJT3mZymJgAmiHtbVnSel44X/wFFZlydpdd7m333xU
wu0kZcCyHA9sNaDsS5CeE+tiCl+D4YCgB8mYJUEsstO27wRKiS7QzTgJUZaWDz4D8iWkOrDDa4pn
eBH5hyJgj9LqNA5xYFHDcK9RGn5BxC8TI408guqJ+37H+nCZ5cgmnXkodnBAbcsSa50Mfkj4xxIl
jI6y/Ag49pJfLxKm0zDRqoF4xL3275yGH/pFZkz978vHJncE4wD9vN14c+lQIu1BRKzBI/I2nraX
Ntc5qNRb5+netCaTdMIcv4c329csIpeR5Avf7WnQSTTz4mi94T+xF2yb72VF7iVqsDvjPdlZOf7/
u/WfakJVQinn79XCuyIDcLUeK/Si8+G/Zd1elF7o4auWxnSNy3CSFfxeSTa0MZkjNBW93ms6vTYs
gF27m82wpYTgXX0BQB6jWmngwoqDM0CqoWW9Xx7pfgo78dCKrtNB8K3W8F+Y0J+AbplriUIFw08x
6ut1Y3Q4f0+gRODZ7vDrlJY/Rkz+grvRXjooMMgJhXnafwd5EPvTg/uEZvcxd+bdzNLBp0O/SY73
RlR5sjZnhxX9lm9Vcj1EF7aG07nQVf9Z4nOsxInh+9NwCeQhemNAeyHgXsoJo5cIA4DZQHrAJjwc
DuHrkw/QWcPwW0zjeGERmpKpyP4Fsm1K5grTMSOdIb9NKnNkEijh7EMyIxmZIUBfiWvg6MDtSfIX
JpuTV4kljmYE9G8+40Y8RhJ2YWmwT627Pr3KnjLEnxCt+DdKNuEZSixbEzdSZa4i+Z0IXmM9S2G5
nkfGVn9+WEQgQssijmuXOBGit2lfPubiI+77cctiojGluiR8uGzIYXPgPblzypXgMCRaa2V2PnUy
F5KCnf6ARgh1xVzWeoQTcKWJYL4EUXMG2EtejhS4WZIrzdqpwYVzDGgOkBXj4h/OIAiJB9aJvGPp
26Q6QlLY6Me3QuHWd58dVCHggnRdWKh4t76BUWk0TgPXb7B+bqPl1Q1dE66T7exmQqVc8tWfGN9O
YQ3D/oQ5fr3tCwc8YznYmaLnOoCGR6JY3TGxeu6oCJfOgBvbJf18uVenL9/APQx+qXgyghtGJiHz
4GvHvuAv+eWVNZfYdnnfUMqBkNiI9E5+cO9YuALHQx7NQXVEmUxs1EXxGbpJuEKRXmgkNR0aRcJw
0/LvJr3cd8ndM3pliMK9b5mFqKsoZPTmdfVowiivGEyrPcKTTK4OFygAOoSwlirr1cIRyv6jLYcJ
4laJZSXmLHy9kW0LJI13V7R1pyJAVefULkxKY6oYHHqU+26BsywN/O2wzIsIL5rqyghdDfR+QeOE
luBfxyns1GR3bJoxbRUJOhPTMXqZh9SrJTduPiP+pfm7haJeIKpCYwzaiTssIGiMswKzdJsQCjkj
Db2McAlxOVYc0VLLCRy3gBpk2E/2Dk1ihHXeQs7RK2pN+oqq27RuCwnDhm7BA0EZGvjUq9rH3WwJ
ALJzfFE2nLrxeh1LPBnigMFRjn45m1I34E583baiW036J7pmTx5cuaqxRhe0k3B1g5xg0GnthaWo
hoynyfarfNQBjanzdkEuOlIEC4jNPVIVXZ/8oIPXHjuVfPu/f+jrJTEOfGFdoL3ek2+cOdJIsEEJ
Z6ab9fZYJCoVpwdm9lfdTrcFh7tDT3pOtnsrgBI3UkNI8VTxQW9LT6cvQbdS8XI6AT0v5t37YLN1
I9dGSyD7t8ahrpEqo0tIOwze3o6IxcBjFuy0CRfneurLwW4/MnjF7eBWMW2JSDQ1JSeNmWWWKSuG
GfIcoGD2muADzdU23fJf8oRyg2ZG7hfN6wQz/Y1qFWgGuyRSC8dr/OxrFASBtdTaXKvyUzkYMRoB
e+R44S0JDSYwYqFX+lIh6w+D9MNOItB5npg3mdwWG9YleqAnx5tHpH2oKIqJ07etUZ9iEmwhKq3V
s38yWXnj50PBXZVTSbB+AHeTUoAD4XaqIOCkd8eAfgvbATDaGXSo+/lChT8pHVGhgfoH6nAERDwS
tGf81MM7BGIGJkdRGtEJN01yJJHdXrKOvSshyhoZMk3i99hpGoJLYdmMexcbfUk40GZ/nxo0nCyK
vf5nHaIAY302KR1Dz+UCficVCBdm0+qHaG07aBa3U7LYh1fP4vxEGUdeY4Wvw/T4s/1eh++hwe7g
TgAPjNdNrPgqmUyJJN3CiMQykWY6b5X11ye+6v0C4ONp1N3OTEyfm1EvVZGcamOyQNDHmakDaE0g
eBVQCl9nGAygMSkruk7tzwqcoORerYRZAqnN7AZQgEKDtPApiB/RiHUQp5/ZLCItqau79mX4f7NQ
syRYFHZuVBFjYAWw2TevvfB4u3G5oe20c3YSNE++gRtorWEFED3V5tEnFmpCZrrDNBhl8O1WJSb1
o7S9EsNK16Q9iqhUkx+DF4uuCnXvD9g4HKBP/0A+0M4svjjag6QLhhtX75ZbgPrpRRM8fS/0csPY
OU8Rek0WJOZxOkVHJXZeuKHyD+AeWhvmZKMlca2qW3tpcqAVzAVldtNBYTAdR2WkLonMFz1u79nK
iq2r5qyVHbLPel6yVEEqF2vgR/g8HYkNhqzAx2SEFjDo8H6ULNg9xowKFUv2FwQ3q/kYa4xTknDx
DfhqtXF6bkeNVvKLNqseDnLk+yvPiTOjulPs+Z0fl0VvscaS3yK4brIEMDVlLyZmTIFaEC4r3VRK
mQ7BikxJS+VFooCLQEBMO6yVIA81AGlGwXocGDJ6EA109CXVl8a/7e9IBlRhUzdI65yjsuv70tnk
CAZ7ABVi3V+zkKCPj6hakag3NxqsfEWZSp4iwxF4XO0XqlGpfdeALxhEV0kUzKEMogQuJpPA22vT
GjStoESHwplxXygHGIlouMZb6/5lW3ZDkaVV4rS5UHKcfBaw/UaZO9xL3OPlEFP01spJBp0/ACcO
WWVBcrJiBkvYw6J8ufDoNCbx7UTqTHfLO/JiCOidOCQqDAl0P8FQXZhgk7LX7A4j+TuDGh6zzkGX
yBRIX4XUHcZD2/poLmG5uDEzeILc/SZFEfswouItbmfqMLcIMS1gbWtudSELWLb+kCj6a22r+yw9
G287Oxo/o+IWv3a1wXqJ6ujHjTEdLv9ngXR4XtDdNGVFr9Cfjel3PRgkfjwb9GcFh6iONiwWzYRV
xnTeqPysslbYuc0dyHLxpCJ5hi4JAb+CdNtsAIoxbAwZafK2F0FrUCFPXjQWgaJdLxmUtW2ZASfQ
sfxm5wIL8+K4+mlNneB47ERmHniDZmoQJrfmzSE9b/3L8pL0uqP5LMBhaZpL/xHRvezseAHVpgR4
lMCbzcI0801CiHbuvO20R4PKoBIYppKVqEF0TE3r1cipEifYI1PzdzfKou6amMcqoZ/p0Jp4CtlB
kSfUtNapccsb1aZzEAj1wEaFV4PevvReXEIogiwuvOf4IT/8eTpyE7EWUngPDdj/F2Locqx3nMeR
fJdAqbjdZbuBiCNZNW2KrenWRu+mr1Tuc4i0n3r8WssWVWBXhcIyQcMqj9S20QOsATs6O81aPd2k
gql+u3bLH156/CT02eG8JbyziG8d3k5YE9FoCjYqRQx0ubN09+kcw1ApeXqKGVSqOYZoZvfe1lqX
H8XOuYcSxxSJ+CaS7IALxw1Q3zTHVWd4YwOdF7iY1L70xS07pKN2RMtQyntCG/sxy5RQY9Gwx/yl
Dx8sDAeLFHOTmAsUi+VuZKVJmHNsk3k9Ia+pLZMjCACY5bst6WEy6Um0RRyscgEWDThvcV06f3aT
c2S2YY5MmAgokVqLe17qntCC17HVIlgNK+tXhA05ZsCPNmLo1xTpGoy3wsuvebJwROq0qW8TFHX3
DllFom9M/77WrzSRzyjGTkYum/2RX2LAc4W72XQD6ghvo5lmyaKPdn9eO4q+iOYQLzY2TrjCEE+J
75489e0SrxWPa61tDNUjfx/YDLC7OUcA6Kskd78WEd4M253oj6Qbp+av7QuM39BfIMVpn7dMtsuK
elfip+8OVchwYfLH6MBvTi5d7N638VOQ4sJjPkgnQJk9LigyLKRF6Vbzv6OVkmZETdZFLlrtGkK5
r00zr2qNjmkM9a+TCK0PM+wPj6i1BoTMXkvGhHxDCi/8WvHFiG52cuR7oC8RKBtVRQTRMZE7jIxQ
lh6sc3v+uGmlDzAYPmRRHFzbC9Q2iINvBGiFstIMGHSgZMOokYRwRovef6BCrhNvQGNHB5puB/8u
OJU72XdmKyzpGqlsZkc9atWbD68QxwgVGsyFHo1+fuQSmpK0tcbAVPooBoi37CittS77HsbZyIkw
4Klk1cpdL51dEGdjpNL821iSUQmG80AeC5DXupb2PiZ1lzNxoSQr7NvIwnRwN3CXN86JqqiWHVWG
fYXSXqry3mdbeGfvrXLEiQNXzGHkP4fA9xlybACE37Izq1fSQHmU2+UKEmTQBTHLQRBWXgsQh/Dj
kBEUdkkr0sVNL2G/veB0GRFWn95+0x5M3JjtmQi/o2Lgb9GqOzlz5Vca8J2F3RpBB9ydZ1F/l2fD
GY/Nwc8epyxowUfwOqDgvRpgrlNEas0s6X6SfJLOKpcXyn1qWNCfl0/3B/LcsJn1BIft7CvQoXk6
+cvX1T9N7gdzBeF8cb2XMPycp2XSmydt5QoaM8yqbW5jC3oO5oqKBNRFPqQ/WwHrIb3JIpIhbqZq
kVSo2jWJR22l+eSumycy7qtBIiFxQJd+LABWST8XGnRiMNcbLLS0frPHzkoLaBf6mrwpClcqFeFZ
E+WNTFvGL9DZSNzCyQFTROmvv/RDHZzg0dJbNq7Rn98pafIVJ7id9f+TPSXgMDEcoPBjd0PjAErB
LfggDwdZCpPL7HEDPO1zRiNT/kp2vq3XaeO5oXrhm6I7JpAAhC/da9NklAOS6SYM83QkOM1QYWLA
lfY2ts+Tjpky/yeb2HrrJm0jGHY1oW/4NZuuyZnGyN+7d0FALh1ifT8GDonDs7XuaAZpRE1TgJEN
zlsy3fuuscc0NMbMceMMRDUMlDiTQN7XzxpCxwI1JLvtiex+WlFZnXINE5zJqJRsnASQXeO6UT3Y
27m906nsYw+XeXke1GC+ex7q6CwI3ZWe/SR6nASaAzSqe0kej/pdCAPzodwgmCOruiaRluIWUzwc
h1tlqwni2HV2KLrdMfKXsAwnHn9bNMOK6PeVbWfZZt3W9KrlmaBqLJKruI1aVr33vGk1Qh7HhMjM
xgclWp7UW1pRj/TkTe0l000n+tVRwOEJY9Zys4Y50hoSUgBBok2g+cMN/CvgT6m9D25E359KCbpy
6bFOAPZFL+1ndwlNaVED1sjvev67JFqepkxZwdu+M3h2WXeNsYf270ihBnGsCre2hrLzT+xHuVhd
RUdK+dpnXPHTOpHi2l6XQTWV38mKkDc7G9t5ize2X8OBS9n5tzCfkQ4eVcvd0v1ynBeY1NZzJkI3
TcHd9kxTmG0VARgszRn7gf9li0Bu+HF0c1tiSg+Xr7aiZj4VXgOfvwNoZRYpdS+Q/E3y2ECqTvga
thhgiZmSNV4CDQh1b5UHfmT0IFbJ7M8MWXbXA/g5WcaV/Ld1zhnQzbqJuG6Vr5xgBHsLeOhoBm74
iy41bZq7e5KecnmPcOJ5J/GHC2uPUnsmwzMlZe5wIOOiaX7SAtMtD7+SX9e6qpNp499tijWvmxQ6
W+vjUjr8z8w85EuJeGgVc3GB2oDgOp/dFXLlXWO3wkRxzsfK5WIDNA9Byc2lkO6zk88W7/JiMPYf
WXhfBtebWpNs9ZuBx+/V7/mvJ2l11cn5KUrdfezluoKvEu2rGN7yytSC/HaP19Bhbtdy/0KK+TEI
CxJIH2nQ8H3TZH0Y84sy9oEuFb62NF6NsrEQOS8hXD8dC37l/1yqYMeOCBby4PkgS5l5USVd/jz3
hom47m9APCDRRKE0dlT5NWd7nxNQB9ULHm17Tcmf7Ra1cewcLYRbDULe/+tZqWJ+RANhlTOn4fLc
hcQeDPaJr5qe3pUlrnuHtWnDxtGIMCbxtGC0bQQZfB38xdXZ6X6buujgChEx/ieKKg9z+A63v5NX
Ha3Dbe66RhWGf3s6YlRKgHfQmtevPG1CzvZTB/4+CNw3qSLsapT1gjGkuV3ky7vo77TLLE3McOM8
8w8e96gWUAZFGh4IMEI2rT6bNFF5JiX8SANcNoRaqwnmuilq8JPxS+qolWR/H3CDZ15KClGhr1i0
lTKFTJDygND/HdkQJpi/NRyzGwcczscHQy/ORjZkbEQxpzgr5j9JigqWbowweU/PEuhY7k8tCuu7
mlZKG0VsPOyswApGRpW1dfbomiz7jzwMBmIliWrbtC/Kmd6kHWQ00Qjrnz4YrdeJb4E+RdBl5eva
uizdmgfhNpbjoLARrgmV+M8+A/zX9onJ3JdgDPejtfgT5qOKt7J/43tXIqG0o1dm/OLz5kbLXEmn
ggxX45Z9KQ7qSmNDSuDRR2LLRl3AIuLghCMJCT+yBVLg9ENB37pE4zONsw5PwCShlJ36m1EmZbso
BNy5jVNGzpps0vaG8l9MoR/NPcXsPymwNSa+GdNGgLcRiUCMmUHmY477/QN6rSJ6JsyISfEokQ8b
0ThS9XvwseYKXGozWGxDj1JcgDeI4+whtOeYJPTUcOsiJWyNSOmxWqFu61MeBW/vtCqCXejxMSwg
3NcKyzCtX2jCQjTyYe/jSTu4MEhuBgXg6mfGaV1fN6PvUjGCra39t+ow3TAUR4nDTQVYafCDf5ud
nw32HeyFdCmR5mRCDIVU15zHXVm5KzyW7ocnZoGnA7YC7r2bFOYOg30iTXCsOfzPuXcYsRIH5ypr
ziJ6JyM9N+QyBq9uz8iw4KSDCAr8D1n3oyKIZv+YcOczvyGUl+cs0kB+Ld0trgoyviDwBmb+IPhh
w87Sx0PYs/p/r+dMFGojLIjYW9y/MTZdbq2kAi2ZOJW7MHUyO29goX0d19m1UhCe9H0fR4hyIQqu
kPD8ajEbxmXAbeCeSSdt8jpqbjZMLbSKdPnKdt4mo2DTTU8PsJ824MjX9HGc13eUrpkEZsG+KX9g
LsW+rxLBbIqg72KVP0WLhJNQO5tNIowv2KDL6aDQVSmr0DwtHRh9+pSp00Oc+82xCrkhTZnnvvuA
SZkmPF+zOCWP8CYAV9vUjGZEYabX5m2DmafzwKGe2Jh8Fk40qRRLwr50SW89aQmewWd3p5LOLl3G
/KSVkRzb6hw3Tc2DN90mgEbI4b6Gj6XlKS+6Tn51Ot2FJEbtvJ1/pOoHUCVbxxFP4Ifm+Lb5li34
7PQbre4Rxzb3X7/eIkehdSzx9+JK2rVad+APEXKqP0/MmS8cnnQWP6364cTfXS/fJM66whm3MiZK
f4GWQmn9pdiw0aYeCrjkAlp+Phbzh9+ymLj30SysI+Jw6CLSWaIvtEihwcU0URrfu3LlYoofNCaQ
U/b/dt83JDXjYYG8a4FEFI/MqJmlanZ12Bh0TM0l7BUTHf8DmuepvDfGUyD7OXJ4DQlKgZiNV1Up
LrLaH6xchXOmG+f49xpK0LhesBF08mWriDnNf3qu31J54mGTNbpAYFVE8jaAfUeEo50QOke2nFZI
+V1VzEuN6EEUZbTdJWRNOX7LWNwHp4V9qXTNY6WwpaLUpZAyyAr4inaXolIYx0WJ18KVm8v4xv6L
pkic0icpef/CKKTRqpXcRqww/3OVFH4KJ4rVFPj1muJBvRNHbvb/RNddb6YOXebh9pcqBnaXMqF4
1cf+s4Un14slT/z9BQJT+oZiDrEy/U5ZhiEdLjOHCO7/lMM1UVrX7JQN/fRpQ0HPLQCYI2dgWGd8
CD+gMYvXli7IaC16HkeNwvWUewh2Ldag4LY3Zp+BDTc9ld2rBHeiMSB8UiFrVfmNhyK8ruSBImYs
5Uz+Vlpg4yyePrbfLbNziULDaxM2pzptoPLgFNjUhq1IgVkg5AIyCiQL4eN1ivKmK3YzyV9HK5tb
2u6+i+g22IQTjCoePLh5ROsbQByzeF2U1SMYu7a8PJ3HKaNDZNSHGuJejITXG6s4eGEgEEko4ppy
lePocfO9oHUV5pqMIErDuE6BnJZwnjolfpi8FwVH0yCfkbplYijReTX/uB2RigFb6JtszFA0vefH
eoo1yQX8MZ2AVlVYLfuLeApfZDEM7MpLzDQ81XOPjepp8jhW+Lr5DzsmMlsX3cLscB8ANWtlAc30
gtZODoSpllPDQplBBJgH6qTRjRE64x9uVd7kAJfivvk5IN98NxPYOroX5A7Kb350Irc+mxNT0ufr
7HUh9GsFQqfEjnDgY+Moq/8unymNeeMrMqRtBexnmMSet/098XpC5Yb2WWw3nrjUG+SAPvbvl3sF
KvQfua2GZ/Uw35ifjMRq1FJxqgBmMv6vX7wJx3j+670Ns9KBheuF4FNezpmivqu1bruAkm8J8L74
Pp8STIJo/jB1PEBg9cRfu1Trl0Y6P7f+WfHdhw8TbbqDr15ykZYeIK3B8bAwl3XrH7E8LtkI2VCK
tDW2VRzsP1pfNPEXr2pcL65J1wpguQ9koy+y4So+wTI75xtEpoweBHoaKEL6MfDEatyHzkx1G2XL
UJHPYIkkoLA8wD61N+NBqEWXzCg1H+lJCyh5tuZ9Hg90BjSNw+S1E83pqd6AMt3NzRY+6IXCZJSx
vJW4anGhepjBQ4WgjCEcxwQq8nABpx+HIA0RxfF8Kr04+z7rUSg2G0ZOCl0MTV/UdEMqfG23EiYH
2Eo4Khwoj1O+t0iL1HgjAJkTtKrOvjFT/ZwRUn0H1FRlm9zwq8i2a+YuN0kBQB6MJ2Gk0Sh3T5kH
c3KcrDFHkSlunw4ASh5vTTtBj/on4HVpLbCu7L3QCZc0GuVJsHlh7oll46N36GM5DAIUmFl7MS5A
hV8OVPwvDG+/787ITfX/Hao4MdS0bpTxUhvKIe+Zdv/izmMUnI73eLBEERBBYPqlNxYBLogWW41F
lCkFthho0GDjQq5NR4RznJ68O1I48QYeGjgYtStIPDsR0DlES60LPRbTYZT3Ix7f9ttxrJscHkDQ
OSvgm1ctdbleQwJ5vvnAmLJnDf6CjwCIblx+wDGb9dAHFvJ7JdXf7kjKvYF+HD9zm7r5/piyU85R
LClDv+K/XIcxinM6tYK/A7LFO3lhgBevpg48pm+VtbUDzjWLJDpI4bv3vrQkBTVHT8hr1hNNG5yc
SwxsTy/ZIK9ONV9niKPL8U+oniXdp7T8Ra8XLPBNNeSz6qe58mLaobE6onAFDZ1qb5UkOg/oQP5v
RWh2mcTthT437gXZt+pGRMFlHj9qvPYcNfG/aDasFaXvBmgkOTuhCGngApcgGvQdVsxhlPcS30mF
vNkEnheC+n6ERvSfXil6ffQ1nSjikOtdJDhEOTQBUrCTQMFNx+rKc2dTU1th0yc6leJyNsF4EUoV
aHvIUZdA66BQ5ssEjJp+tdLp2A1XirHld8DYtXsMYfP8vkgsmExVCmCqRqWhKOx0/8crVgcZL6gL
xVcEb3b8i/d8LTZz3YelJQ/P6rlOPbrduyuAc0wlkbZgwdzoAeIC0FX3NBCXx4ycwh5s4qMTkX1t
QU/3bP2AyEU7gPck6HvgG+yHhR4UyUWnNA45D+C14OXnuKmCCgEgBsFIkXsr18+F6pLJJpnvGCPa
vGgnv/MEoy8tQiuD3IJKDZN8AoLXSB2qgBGMeqOyfTPgZK+djr+o7qAU+K1RSjtZl9newfCcNyYf
6crfZ/IP9WNUvYmQ7Aqe/78cnnPw3KAjsQ/H9PL6FrJjRIvbX9DIIgvho+0eugWXoz0GCqkzkT0W
orOkpu2xReGnVJdzUjLoXlMoJkWletJiStnDZstGm6ZpSfWo1cqx9mXFSeMikjpRzTCXrdOvdBHU
JiiayvT7In4M4DR0r3MuO2MeHj0Sj+CZ9tJ0npve2ChR6TaK/GhzHm6ujGFy+PbPjupGQ3NQJlHg
fqkR6DMoGBokdo+okibAR+82IDXx035R0WxnxqGhnyj0K0LQqpGXVDYx5uihlsYCYi1AZzZ93iTX
P5EHNZhy7fmDT6scvCZDxD73l5uqsvWJTbDPaQZ12qoabmHLUvVkAg1yic9B7f1f0XIXh8bjBH5b
DkvIkfGs8l/vDDuf5xAgywS1T2njkjBE/wPa1CILR/dde0Vxb8w105bFSqXYIOYscwSv0e+p9ll7
mUmmIByhzj/N6nwq5kB//dm4t/VMUb3iUKljROkwiKHxT1k9uJFYE6EoCdcgptIiNQgr688emrT+
SZaZulIWLg4XSEdzLIX+5kZ9s4VM0jPRfAx5ajDal0FyyWw6/6WN8ImPmzdiZ3tI/NR2dIWjmqfg
vYYPsEDm7VRZW3GPKPJc21hw4A3054+yzyQCD71R0FS0YBWa68pTEAgjIe6D2VSmFfCmWqh7WnEq
fvxgfIoemc581AjBCGgQHmnmUTOF1YeeljkQGRZw2M0ZjdumJqDNKEET0+iHGSndxhdWd+WNF2FG
nxNY7whSmb5uqgKrOVjSzSJVtr6TvwdYy1/4h6IdezfqURjVdEa2rb4Fgg7Qpr/E7K3mPaN+BvBz
pS8mR9SRy4BTixjyguUqcieKPYvarlsMHGDcGQpfh2yYpVMYf1VRJu0q33rmm4vAfD0c3vSTVRvs
ymqd2QxhEG/5rSHuoNCmdX/w/6wnsbfJFF8RhzTSXWNwHUmXn9S2iOnHstCBUhCfzx4nqR34SgOj
2fM/wirOmZ9kb0mpnO1Gi+BSQau+mkP2B9TqYVu9Q7W4Zd7ZZADq0eglfgnDk/r471V10H+E29zl
+W2DPdn6zcYVbrlQ6nqhXlm8u/6IpGa84aLaml2cMTBnPHITVHcxXddiNim/4LXQPW3PlyhxoY+h
wY69cDvFbSfLaTDVTmKRAw07GJIqk7aE56+TGFBV1IlHglVaKafpEV6QZpgc6UlteoXYRG4mZWSV
4hDadqMglKjzJk+UaT/15IZZBKXfkPGvxhTTDqNbi49mu7n4GzWh5Mtz4T2RXypciF0zuFArZTiF
XgXcJI4v86EPNJPxhTrnP5Bw9/+aIlA6DLukikp0sC4UiOhZLqKxt+MCqgjnBNN9mkF13G6td3Pl
5ZVrqsfilpW/uN75TFSzWQIkBjgv5y6JaJ5/p3Jrb7J0V5NRRk+d3LImjDxx+nTySGsrpSwwgfGt
JEweBX53FiKmHv5tlmGeQoOI9fv5EldtFJisVcHmQ8kkjZSJhqWHQHUq3XxBT8lKSE7FraPDOIY5
tOQs0N6hQEz0xIbkInWRTiAPq8UlA0qyuf84KvOKvnbvJ+mEEi0tEzsa10omRKE2lG7juYYjNDrf
XcU2lf71q3AM5pCo5tIzH/4MHpEmfqFS8NnFzo7jEZZGL8wR63N++UsvlRMBJcloQhCQ3j5jGo9B
VhFLTt3ot0Xu2KiRgnQkkCiduQLlQvI2hc05gQ8pBBajzD8VGWrjrbc258byIb/p/LmV+t6lz6w+
lTgNQO2Xh9db/B0djZfkhX0VHe24i5t6uWZwhn/jDWsfWzA6/ELtxeDNHr2qfzikwGpG7roKlV9f
3G3NOImXA3FUGAFpv2alvs3kVyAugqt04hBF4KhNE+Ggr1an+0XGSDb3O1aNxlglM0y1ajlfzUNT
nKpj5TgODeC8AKo34Xe4gSH/SdESiXhIMJGuvXJevahgFqyUJ5WDjvE+NrKko1W2KGm7+14S4Wts
Ge4PirehUBFubogrtaye1SLR3U8MiLTumz/wJUohPOvSfNYn4zRerbWoSaUcdWMu2ZG78+m1OIhp
pZaLmIJ90n2baX0vciJzAo0gSW3mrBao57gbpHIZMyNcNqoRVaXoesZ4xlHke50BTydNtv68QJV4
9xtNVrKTjKwgevUInKeX+3xG8wi/+KbI+7J4PZ8+bOyAwhHb3o+ocp6saHf5G/cdiqCJlXIQuvUA
ca021jXYmRNBFbZDXHZxEKMVrbgshdte1J3oisG9NT24ZgY+xXxnE3c+c2U0LRavVnCTZ3xYSwhG
5kqzAJipJSY+PGy0RRCUn1R7gYmx6dYSW+y85nCfrYHlajVxwDk5tMpvFii66ws/2kEEpUHqDCW3
BWs2CzKxErvQtkoHGfek0COgr7XzRDfujgsoFTtpY3UgCkkZdXcZU8wMOkWNxPUoHdgQmQdQEzW/
+y2GUeo7gble6OlVsJOgKhxSgwxeAxPOTqW2pNWV17idZoJmpNJXnsgj8MqdPVNajmqeTE4xYkU9
md8sMpoZqKt00IPdiI8pKIFnvqrcPrj3lTOANB3MxcLePuRJXIEm3kAt4nVafeQ+88iVxq+RiS4l
XhXmA+52JimP4PqHr0onbBcNA/ihqsxanTfYggar/0nPCt40TFfn8AgHuqEc15N7fUBJhAGfORhS
lGoovmrpz7Wd9100bUEE/ec0ZZxSxi2B5gftO/vHWnvyCye20l1ODKz+oL3D9VnGbZMaNMThN3Jf
MjlknFzm/F0/aWAZIOTKiThGuvSljK2B3NSVovbOrTcH1Oj0U8yEDuRs9HU81qd+2YWg8Dx15IAj
yfgSWKUKcQsmPb2s3MMtWyYMhTBLZkLcn792nSncxjJLP9BFoqJSFXzqoeRCKFmd1nzpdv53wqiy
OceiCqJRuwW9Qaqcbkcdgfn72ECD7lN+D9Za7vsbqkb+tRh9OXk2aaGWRuWuwhlufkMfsvfUytXy
qy17nG07lw7jXIb9BGGjhV1Uc09ZzhYKicIWtRqlY2GEAdWlpii+IYGzqqfqJb+ZFTXRpXp6m+f1
pp5vYLSzeeBzbrWFiCm9G9XeDLlVgOn3kOABgEERpxWcxAWXcbU5qTttMK9CrfopIpZbtZfLOlkw
GiIMviNX3jAjNmfSOiRP7xfZ2mNZORxIqxCH+hxfiKeRgDfuKXQWyzXcMlSvzlQtViDNRhRE0h+i
JRFWKEWo5cIHczilN5KSnuTx9HoQpYol2z1xoDxdTs5pRl+4LFTzG8PiAEzo8UNpn9QJBTAaRKRT
7UOZMJVUX1NlzsE3SAwxpInkH1HNP0TmZoHawmLE/PFqJRcxrXmWzfA/9jnYxSPVZd5zk3hm4Ina
hNcJlgfr5hlKIgjByNEkV/8VIJryX2krpKWpADHIi8ZI7d2Iu/dcr61+SFHkrELr8LDiLBWkk/ij
DVfPl/ApEP/Ty7dKmkIHTxemIFPSaalsVMF34aq9FfmsRNXaMQZzOGnzJA2BeBJC4EJLn97AL7Ky
PMi4Qzw6jtHfdkr5+0Aacx2vtlew/mmGSYmYyzyp1L376HtW+YKah12py0Ix9WnThnXfk2ONTnX+
Fav+YT63rJyF4ddpeVkPQOwkocDrYI6ZaID30vVHropPOminjf1ZqJjwbiHMeM+j3dHND3oVY3Vb
FW+tWZBmZn9BD3N/uL0m5amt6HhkPpTHqsY8+pPM7tFXkB0+Vs/I0Zg1bbg0s/A0422er6KOW3j1
t7j6loLQ0+WwYgs9c+TGuTfPO2lDKgHi+gqT1gUIigpu3nC+ElX2r1rmAikNNvTMJ9TEypL4Q7vh
5tp3iMo8xW2FO2Ahsv5kXML2itaBdzNpfkAuGAO9/zC9DhJ3Ww9WXQ/Dit5aE7oqILgPWIV64L0t
9VXneSGlZD2cNQSnQWTzfOe9gQ3iRDUrDVlR+Tp2DlIMf7v0M0Lbl4T5eAx5zyxgC8MmSagTQeLs
dWg6Dz+Bxp2snvbui3v0l3OxhTQML8kWv/dHmn/y4k452Da/mxQTrbBvKCpZPu59wEHx35c4BB7J
fb4Amf0S2yg/0RqYE56yOkwTN4imc2eqhstLtk4WtCvvK+mN6y7KYxz2NQRgYpvq7/AXR5c8Tuac
zICOF/0dVVXEx10N4pWV+07YbZFI7QCGN9dZ2jCIHGEceW31kZS4m1wqM6zPxUygPZoE26GKMkWK
G/KIf6sOwwDd/mYn/KPp3ZgzvM5yuAAqzwRqjn9HuYrNhFVrViQjkntExS2Tnc0EQZNhmzKSsHjO
90Hl0vRW2O5YK1efd35DhkusntTIjqh+wUL76uOat6VjyBkACZmWSumytp4mUOHP1VSXy6m5XDfb
ltbDWMhDktH6bxQDBB8a3G/AOkNnJ9NOpESISWzemPqXuVpztnLueNcoPzxRloakrmkMsylm2cYe
ru6pylnniXmwawbJyd1/5LMPn0IDDcbH9jhkX03q8qfgVZG3W0tlvPLRVzyef4HpR432qkyJlEmB
tRUxxC8yZ9iVzHaIebXLKNGwHA5uZ8oRznpwFUC1IFi4cwgI1x72w/7CMd0FJWOVpFx0GSbajdX/
5T95oNH/yb3gTg0PL4+VWYMbazXZItMiBjK/0/jr3nNxo9ougj2C9MhnqKfFNOOr5RYqnyrayN7/
Bs9PxJ5rgvAjYFD+lNU8yd0Ld+4XDNUofSoKvSxWt5uZE6WLZxJ/zCY3nQATfAUJWLbxkY8VK/c0
7RHv1ScW97pA8UnUVnyaAHuFKowrYP/8/QqOpvFvVE7h7R3Kbui3SgCDuDIpe+h07y22QeyAh/qb
aSb9M5NDOU74asBGuKYSoUadZlRodI5stzwzjP7ueJBOM0h7+mr4U9O2OLOiuY/kQNgYStK79g5J
5kY6jTDVf9SOrLA5796v3j0QJxbxIAKH2pi34/pIG2DmNEn7wS/50hnxInVdeB6lroqD9F291WSk
ZlJ5L8JRqNrhUB3IAWyDIf6w5BUuaFARrojzHT5X0Aq9OxvjUeuSAigQ4IXNk2PquTbyQ0vPpKE8
aqRHqHdaegOTf1YrfVO6mmBls0MMrG8ek0sPw6S1M2IcJy03yU5cpRMNSql1IjaKNLn3ZweDOIj9
WQrEHfTLDtjj07b2SSIslqRkYe8yJ5LCsoOYDo2BjrmVd46jR8G5jkJch0zgksbJklXJqRnPnr6L
z16TWz5+kIEZ6XpdY8ebFePW04xYMPLXNyTLCgOridnGjUwyFJbofOE1N73NWQvC/wOdZcFsTD12
czb0+3o1fpu7I7Zq7M7lq8H3AY8+3m0pamE53+aY594y6TNJoZ0bK6WbvxpN+Frm043HWtrxq7Fe
/SMML8hjptAg26Q8xD7qV+9gdN8ti9xSbHcHo1nEKiGX8Lp9CTsRIjhaQ48nViokBEN4pFQndx0X
oE1uL8zO6wkJI4IferdJuzadfx9AARAydDWZMtCEVsZftaXUPmqQXanWTwXoMLTnAGVmHk3vaVae
1CCL1qs/okxfScf1jFpR1y+4dlT+M1KsD+FJ4VhN+qHUB8h6oFc7qwOgVzxY5/U69i3QFdybs+LZ
c0/4g7QMk0HrkfYG4Nghq0gx/eNzLPQLZV+rhGOdCyLcph2M4duWxvb6vizFGnD30594pVe1bUBZ
J2qem947nltdYDKulMaMu9QNcFWzPQSeClWAYZN6xSvNiI/a9UFOYr4xVrICKhHnTin5obJlEomK
O3iahUVLTh0XGJOhXUeqnyXR/xdmn32r76H0QuPi36W4CJVFY99N6+vislgb9dsk6yQKdCIhu+OQ
+Cn2EBhKKB4iKXZKL1zTJxPYTJvtfTfMqOzSDGY9vO9JEI7aFe6N5aN3Ya9/3x5/sNEjUutqJCmF
SaJNHdbYbj6Ef3wpLT42A65ySiWf+lEHyAPpoyc/l9wiO5uSIbevvLIbr6LKOaU9hl3c3UHx2IxC
KYfHxwMoZbCbqA84Oa6MniJD9JMnMbcEEAWwgPYS+JoUn62eUicW8vVB5pWSEpiENv1+ScoT1P+J
kpKPnWVB3zwdIiSJccRTX/2xKEv4vW8klUgZ8PF0ObmiPSqu08fN5QNwwcJj50SrtDK/VDYwtnmB
4RQaNHycuAVhjHAdvjOwoa1hqBjOnU5tOAIjukW6y+C9apbyONhalBnp0EDWaNwvI8ubZeQ8zkB/
uqwItatYYD/00bSlhvDdYQEuKfsqAh+q3NcySgT4S3x99KJEwQQrl8JBYPWmrpWt8ISFx96v4G4T
HuXMMqlQFUrHh4QNbLXjJMV0gmwWVPbvRE7l4sE4cecNRGusShGrHXl4fFjaeN7vn0TnuR696AVO
ncda8w37EjqIQIf3m6GQnA62UbJUwlmks3o+J3WhETS4P3mscURcGPJrewRW1At6of36CUViyiHJ
39hq+5AHiL4OpaBi5t/Z2bAlhEwtNlINUHfmXdh1ELD1nt77DVq8W6txTzl84Nz0F55jsb1/UiDv
PA/AMYw885QN5vYCjaMa0fThex3yFdseanVrTQSh9thlsaODQhOh58Neu43Bcv92/sEf8kTJsqPF
KvS/+lWeLykvczMhW/4a3rfRWtHrW1mAO+Q6w0Jd5B5rx1Hu8GrXSrRJXLPY/6c9EHABHpxEjS4m
3z9JgyWHSpQZT6/Hg3lXUBGOzMVkMsU1Sx8GNC/V0PYSC06rgSfQoDfkaNuyhlhXgPIrFD5GUx5e
48vCo8hyhXMYrwDFjv5gFzsufnvQKQAvhGc1QfZGVxySRuGIEEHc2w29J1V5zJ+W06l/5zSz6U90
B3vBe5c6eXMemyxcheOPNi/samEupbQBoSGqLCMlFRALc7vHPe9q1KishJ6aX4V/poe7WxjKf1Np
TsbSCaKFp5bVGvwj5OUyMd7vFGIhTZhrl+1/49IWY+EeA5E7R8stsL3+k3uTE7M8sHCGQUD2G2nb
s12WQmafpH8HAOHf6X24+HQ3aZqmetx2ZVBvUQlNxXRQ7zZH2Ba3FBAiEMQSwqHi5tMGc+eVGMI3
ImOO8b9kWyl9JiR4bsW+cLC8NQumeVKm2Z1gt/bujqb74zDGIR2V6i/MMipcauUORAhu70MQAwyx
10w7dcUKzDAVHuMOFgT8kAD543SSzhIZilt6UozKh/DakJRl2Km4AcD90VUVdqQmTi/yxXgD4GWi
sBLEDuVvgBhMN32pV8JRsSj9/ELCBerh2Fys04eYwX4nUA5fkX5wG0xwFtWi9+4qRIByxQr5sVGS
nbimnCbl6Q3cGFLtuVgltsRZSYN1vaHcVdFO24y3RsylOxmtzxbds+mzHE0SMiRInzxpi39+dacr
EKu0n1qMIcq0SDR7MPa8b/7WcuU/7fwPJMrNTJPelNYAJ8iEEJJqeNhbz4Ey2XQjc8jbvb8gH/qU
aCorKvXGRC7z+DbHH3+N4+s8ZFEHc7i1Q+E2dIgyBik2rmijWsiwsqWJPc1UBJoseHkdQRvHwfE3
mpM10Dfx6Gk5rn46ns9jAk+LFuq7lVv2ofbGUfKBJWvC7IMbr4jsfC7BURkPsuNiqvLn1CgeEop1
bal3eFNTXJfidiUgtVKYjYfhx9P1+XHidNW1gwqoRfQjgnpE1btY13nTwCvpHVO857srAD+l/E59
370dXhNEUCpjv2DI3mQM1p3cMPScoa0QhIP9mPtIx58BaTSesE5lxKAxTG2MiUIFpKwAsC0WnAen
R54hc0rsbgMMPs06foqsWIh8SRASZ1wbY955sgNtz6xXJcpjgOnCeW7A+tgyp7ahB/kcM2b9OvpY
DsO9i7Jrp9Sy/yvdsKSz+N0DgVICDI6cHVdCbfFKt8lhsXMFXNTokYEcD94f+ygJ1pxrgFUhzt5I
LrzINJeYuErUu0eLZVLg576mmZaOnJIkDl8IDDM668LDOLEC8akZaUZD8z5BRsQf0+bBkk3MNOj5
aEfthT1jE+Dz3OrQKqhG+bQxzB17iEoV1bqtiEBvV6vS2a/F9JgqL5LzZFNlTgn31rbb8kDXGjxk
uMCL6w7Ju5yWiTJJCYgCMtrIhU+YEkD6OGj0V4ja7tmpDjueioJTTBgosw9S2uCSzsheKHku1bJy
R3uyPAhBNPSR7gbYoyUwCDSBUSjxZCvTCrl4KI1AGaVuTOqmO11DMmo/bNghJUa3MIenrGnAOrip
z62Ne5/hewMM2gb9l3i2fWBMJCSPSuwXyYuSoTZdpQTMGbACXFuwFW1zdFQ0bPElbSao39J1SyNJ
dwnEP5qiUWyqwnwAnuiXeIy/ryLwRTpO8X3OCSCfp19d/SmkL+McgwIne5+0VCusMgOr7ju5Wu5/
2nSaBUDimsFPN29nNr5fRyIOJJ89GEiF/IiHC//oqZMzhA84tMgdoxR3tZ0iWq7iny282KsJSFo3
SPxJA8ioweroyMjA68XuAoWuR8Eb3x59xUXHVWwoXqQlXTnv3Sg5L1pPZ4y3Qwk5me9zP78gmg5Y
YyTO/tSTWyNwUd6u1BvlDcJFBEdrkIkWfOiFHq6QmixnX+OY/EA4FLggLdnQDDXo8Z54qsVbmN9B
AXZyjv872Xka3ADeN0/ss/u7DS2K9ogEgEUanbHTY+hCaQWiwNNNEpbqqmec2fphs/IBm+/ZLed/
wwOE3/sjqYZ2niuANR+doiGlXpx90M1g0cwAFWgiLWn31fQ7qHHedyJzmS5EkG0vzrH+lFnovlKF
Kjz/KegcpLnBP44/aQAgujvn/oGBYjk2PZNXpmBfRXVM4HW/QYZRKnn6XCE+pbtRbD1hS6XtYMaK
Of8A6Iy1JPto2Vr3dqG+h9a3bVCXEfjVodmg3j4QVI20QWXJg9A4ublMYq1IYMf3eefg9kdKUrTS
wkEDj0aE6KX77RwowBdd2zIt6oatZMAHSD1kQCLIKWgVVcsxPWNDCKRaFvRGi0Y0+uaUYbvlNmwj
m3dlRFUoXjVJvCH+RVb2ELbLHJWBh+G+ldEHXAhZ3HXLN/QmzqXcbIgBDwAisLj+4zQlUh8+Ev2v
cVOi+yXwqFu4ASBY8WgwhpLPWzjOeBhe3U3gvWzeGQGOust2sLoIubkr87t0//mitzO8+9pp06dP
OOzm7zgAoSgAhctAhOOrjgp4ZMki5A/vEIpmGYXi8TeqVz+gdYSZOlwobu3eOyd2OeIbliZdl+R5
qiNOc1vE0cIHFhQcVv6EvJ0GFPemDnYDvxZ0Swx/eqdFBU1R6Vgu1a4giRPFzQHDEIlm1ubFXlQZ
rX7HkQ4/z144ipxcCG21KQjCl79D5u1y+wjvBTHActb/uEjgy3oZcoGbGcAg/LwDSqXf1r7zI8Xg
WgTXGqZJPFPm4tmYuoW+onlP45KkRXFwybxqs4NkvABtAQs2v9Ym6kwOENZcMFoazk36jORZXe8t
OEDSc3BxyIZt17NFvUxTRyd64VYPZj3MFY3UwL0Fn4j9D7aBr/jlvskte72mF1IdX+gRypCFWOAW
wjZvNHdSnC1kgRREN6YFyTGVW5+j8D42whNHcInrmbcBzXwgz/UoX0sUVEdajlce/rebEzdMla0r
9DR64By8kJLcEKYud4ox0ELbL6d1PbKSYMhiN8O6sPuz0mFSQS1P3VWLKfMsBVN3V1fbeg/rbe7+
gI3+IhP6VaTacYBpzSbZxu0RUP0WyyiRMQDvLYT5ADoWTB+81hIpCszA5LxUvpcKkacDrjlylNV9
zSS9SXlRDF3/Ung4mzwu4Oswh7QeoLNhP+1n/nXAVwXeQb0Cz+TlyUe8v6i6NzFoQEz3mqz2KP43
brTeQNqK1HGSJd8AKlSmF/UQDK5ZoqCzTxdHh/8HiJ2ZPIJj2xhZ64hDQGfpD44oerkezs1quds4
UdBn59oZPDLKnoGt4F3h5QIogFK7QKM5aUbLkGOdUXsP466K+chKeKlpx2XfItTo5Y/K0PYRpRMd
B6X6IxsByChR35xypxiyH/RO962HVsJMUu+ck30Ewdl20O5iLU6HVv3YDURrstLEo0r6+MfGpNhw
o7gaB8A7imrFokLa4D+cr4JUYFx4htXL16AMiNnxQC2xkGUCXxr+2Mpeb94F6bjXdd3Ie5f5AA39
EosscKa/KW/q/xXyP4Nx1ucptYlEP3f8PIr4j7W0e4lVZpJxOdC6JX7WQVH47FxR9ngCFG4da2Y9
uz3qNiebH06303mte23YUVc7n9EOSScAqNrtQ6zSG9GcLNTo8Ct/5dNzNGqZxPA53lG/I5eeFSBW
yVQKvAZcusCIQQTx4pGxpEh1JfAtwMyOLOo3fqjs5go3t0UzDcSIRkCexB9DVSfRVi8oFQPjC/FL
g/4IBTpDCeSaM0PGhoeuC4pCf4ZMyExANL3/rlr8UMEsV8aD3o8H+/x2wQzW97DrtttqQOJ3HWUy
JZGSZCwN0h2uUoKoO8zK0dEQFmtL60d5DZhtx60BqIpTYnjk2Yo66zcIGcat9loPYjsXdb8+byhZ
JZCbLP1oYptJTmOl0lFppgBgUlFeoFZt4763F7E4MSzN47csl9cV76nNGspryW9TWSEfIWpuqYE1
lNQJFUqmvyvw9eMQpzzYsRLtsgVbJ74+jmGlLu8GzSNDzENYSDzQScWTG0plxqUjcDR1M70VMjFh
feyWiQiX+uP3d8vFbDDvgUrs57gD00AglWfkVo8QCELva/69KON74l96G2Wn2q8XxxJazh8lQUxz
BOH01avdHOj5Umds5y61or+yz6ctHDuCzXfIYrrYE8hhVZyFLaManUa318cpmXhnL6hA8juVvwMp
xaQpucS4u7uY0SfJuyDfXIa0vrRpzx5BgiHpLCPdd9ADug7dL7tFAeOOehfqWuKfaV0koxZ+Su3p
yD8OjnPEup8idpm02tmNE/NeG3f4EIsYkCvjbCtjG5B5yCNZAWKlBwJ3f2zfpBV8zs3Y7wMv40pU
hZGbKfmb9D6VCzq/IWTPfVHSY8obfkSgz4ynXGy50GwU9AS7sWI4Awf3+fVvsHX3BoQSDwMMQbNs
Dqc2upnnMSsocijV9Pb9t8JsPhTmH/l22x+2pa8Ew82WghxWxnsRitYnAH84K58ZBh1WxhLNtbv7
nGWGDb03hktU1jYyibhaOvNT8OW0Fegoih8Vi3f5w/cuGpcV549g4lCXM8Q0CQPPzL9SKPiWtjLE
S/1ZHchP8LzpfKxdHnxPDrl3Z65UaHRXb7OgIg9YyQ+J8jS3Xs4wngBvTwelTmQaMhM6sUhM/oOC
+HMb4Wmb9buc9khOg4eu8F8K6hfJ2EyZ8JOpKMMurQ585F4UzmR5Ss5oFv+qzQ9QmnWScI/rjabW
bz/yG9WSXOP4ZkR7EubwA9+2stBgmuBFexBEmZsg+274P4U1YDIwHKWV+GELjp9gOd+AMr18FvwD
purcE+txKHQdWqwTERAQpenJtsA42oSrJa2cry2pudAGuK6QcGIYMyDIiNlXOqw87o2v97lmpBYi
HZ8kKzXCrhgosVpnOClU4XmqTswU7edYM12SB19PzTwzHFJdIBv0oP0Uh1mwR6MpF2mtBI0tPtyT
8Du7JlpVULGrp6aXHZW8Adt1EAQIfcda9sGmK6swSpIcAP2EHEH7DMl4kjWa0MKchWfhS+k9kkw0
HJgdqyz8tM5ERIQnfdELUe6NJEIwj+Gr5U5EiTZDYEbOc0tMGgNxYI0bHgi6MN6aK7849D4oS5+K
eni/Y56EfpGJGqKR8jw6h/0AkAiYp0u8nA2bKbrcu1Hp3mqx1WceCJJzAWWr2e4jAPKjRgulKsRh
hrWKBmUka40ve/1YiE9EYy3Kct8yFxm+oRK5noZsfwYOHepVtafnXYh516XMzryhwc8YLLCwJIHx
CdaIqrnxXUmnQt2FntIaT2MVX5iRu51ubXlU4KXD2K07LLPrQKVtP5CFU/yJ4Jv0PVys8x6Mr/hy
EFQBlKFoC4f0GixSx+Xm/SYzcD/nzl9EtqAtQjOq1fA7nyElQfud6CjR/zSTA723cMjWisMUbJAu
msqbusesX/QhZdPNVT1mhuJeCuqZ6BpDFN3JzTkSPxRQIO/moPQn+Fwn5+rSpgHw7PDuixmpBVA5
vGkdh79qtR7owdg9yOPv3FzOJHdwyR9W+ZqQvNFscUPzk8vVfpHPvMkdFh5uKTlX5I3iMjrDLLxz
7g5Uc9OaIDoQlHr4VnicXR6Kab/Q9NLaZuK/SFKf+uVRfXT1M0iaGXxKKjR86Q7OMutEzpX1Az9v
86SaFS0yt9tAq0tSZbIxEAMTQe4QT3APLFzByXdNHeHtPFtn19H8Vfp0B9opMzCsi68a4ur4RsNw
B9JjmcS9UCLCCv0Yq+7enIRHUIfLE4xPgxnYiQS3oKyVMM5WVfwZMHF9wz+8y9xahQE0APOkXe+/
XcKZePtAQSrQxc2kIdkNEXQwjz3kKgRyAUYkqNzMZmUJovU2ghA3mizu28UYEmHV0ieWAsVAQN4L
ye+bt+emURyAVnQpbXTyMaAu1fSDOWxbO29mOSxw/bOxj3vJvdIhtayMxxaf0tYobFBuq5jsZn7x
W5k3rfFow2QwoRE/KE86zGDEh64NfedQsErGgauyHVkXaO5I6eYxO5Dv+HXz/3/Ynk2PqD7ZZHs3
GMbpq6LZ46af2daGLr86BUfBkjJ4XozcZCU7PlkLo5GuS6/yjDVNDbGy2fCrUgbnOqoc8Uld0bKb
iCwJSuAyskQbgYh4EIGvEbkqHoAZQ5wvEgKqFsPR5agUKe3iVzjNZ6Jh6S1pROIMAfCl5Ua36Arv
Bcf4DJFoBCS2Qo3MCGFPFwAmAUmCcPEUrDXpHrf74dVYyzDiuLqzpSXWAFuw1LdCW7rLl6STOLay
G56VRxXEQd1zqPIWLIPxAHSjsCweJEdvwsZg6mFgFtRRojab0NZI3hizfBUfRPpleDXKFQfRAV+9
PJMET0fiuRaoe1LMU/1VjGibbUOln0gXrGB/mDiOPutZ55h9RwIH9gLKwX+4xHCRgYuu6VHIHUsl
DpLVVodqi3N7BCICOw46AA8TJlxPRwv1uigOrZuP8yV1Bs7LeNqMsYeoZrXAKHt7aAY5VU7phMCs
FTGkNBW6WTMPqRd/jcsMHlpdGvK4tXeiVMOZuMnkVeFjGA2VBeZBvX/mbJ5SOO4Jwf8vOoPqW+pC
q0RObONZLX7gsWu4yCB02CePcmhSx7LGIPjTpZbhxaUFbVsHhz5cAeTwIsQpB+nn3RI7Xa4memFT
s9775VtrYtS4ZnLs4R2iHOCL2vQWrvulY0m3dWZJJt56+coyKVGavGDoVOOsUsX8mKtGFJTseNKL
kIK8unRKEWPM8WoedhI/5vXSN1cwYWz7jaq8eZdr5WnRMXxhqsD9dI04ocupba7Pv/eo3wBsczu3
WmvNw6v4CP6okM7BGQPWxMoy4E9XZcDqzebkdB15orAHmMg8kSypqalg2434nD1CpQuC/OF9/uuu
Az91JTnEC565ocRjall6qNqgdWSpX1nbZIrNEfvREnuii/6z4YTGW5BzSUOB5PTnNnAjW16vTMN1
FGXffYZgOLCVfPcPyCnm3F9XEcniV8gdassyhSalrU+trykyLRMm2uNgWocNNDnfcroX6WnxfNDK
tBsR77judDX0l3LlhJQ9lvTChGyhem1wWQythRcJi7oT+EX0Fkq/fEUbdNKwycl/4LTkUKBf2bFQ
oSbBZ3snHV2/iqSqT8oZwh0kR0+i6zW3nIKp8SlxhH+2AssB4eDxCpE42SxqM44lqniLqkbBg7ON
GFcR+8nglzneF/Yg8Rk5KC+vzyWJF4TMUfazdfjIyo/xg7BwbFcKgEq443/oiJdY/6G09sxNXABD
uzp9p6UGeWrsapoMf2hCsED5LRVCqdLEl9v7kDTIkp9IHBt4z2PiQGQhstfolOua3sJPp6WzI1rg
TnG7nZ/Owakv4MFK4BedvKf4+Pd4Ecuw9QxbSxewhakgKCkDtCISFmSM3uhavKz+iSMvmtaEFBWb
zh0Vu+7KmSp9pxiRywrJB8s4lWVOvwo6WAZWz/ZwyBypiX8VKQSSOv5sv2S9lupXX1YazzUpXV5b
A2XeTETqs6wlcW0Vub1aCrJvnA1a2aqGLxqMdlnY35iuIkI6HzQJDQZbn5vEFHLwrmhnQbpyoeAK
Fm8yCWZ66LG0ykrxOpneKkzH4Mscx1U+93MBiwsazSyGAzV6EJK2b2WeANjO5sjssaAqnt0NlhJZ
j0ZkLVcp14kxUghzMDKJ7zzmr09Bbq7o2G674DqilhnRzg2QtVU8y7hD+q6mTmdUHdlFgfCfMxTe
C1GFDIF+v0XdbXuQcX5XC7Pd/qM3XVWAtCpJUuxDiknAehf93TfTpzMqB26fQsFjvbXlFx+DO8O3
WMXg/LBUj7nZc5ju2X4/uynx61M0jtuYKhpZ6BWi+wyef4XEtZvTAChisRv18Nci6HsgU5/0Oxs+
p1HQsIp4BSZLLDwGAislrv+3o/a1eOVo/RKv+gkYig7Diz6Eetk/s/0EIX0A6JwBY2HL3IhaiCn8
HJi3bM6flRNdtdZt9AzZGJp99Wn1pRqgadBn6LpnNA+onTeQn2dX5mYnsTX4VYY0OOi765ptmMtm
5taC9zpvQja63ABzHQDYnOKdt/sP5kLW4+Kvpo9bUhRtK1tOxiAVf1Dkb/UBM5xv8HtWq5KamX80
c6T0DfxkSRW/VFry2a/eykYrX2x8ocvJubtbzo2fw5RlhXtIxJUguKcP9YFwlAktng9dcqaSJD+a
0aFnqLp7pHbpmEbWWbkvorTlUvkT9Mak99JDFEQmG/VS4bJjb7h48B2+gX2Zyr6QgP6+S3tw1Wh7
T+/xU9Dq8F66HnSWde3XctPvy3QjNqrSdr9wXlzWR7JQDddIhQzJFxchE5Kv3i2A8xiN349LYlTL
tkboU94eMEt7d0BMby1YJBiLwM05YKm30GlAuE/3iGtKry+nilRPreFR/HqPykJxLxgJHTZYyxy8
p2tBAgFF72MuOmNR7MvQrvkpbmlF4M8xq2MYYo+p8QmTjwTJAuMEzkNbxkEvT4466uJldVsluYf0
APXoHhClTpk+09XvsJJX5XGBVMsCH7HCPE4vb1AEeteiMhVguGNrx48S4HFtG5VaanPXGZi42W2F
QB03N5vkpNVEaXfwwFAIQQrMWLohJ96hlXext5uj9Y4wO5gheMu0EqKK11GLnvVKCZJxNL6womX8
5OQZPNozDcbHXhOM0f+HJJrm0RDkTabYNv86O3KV/T5OpMMC/7++x/sSlCCMiCKs9jGXHpsSRVPv
q23O+NVlS/1JW5LL3l+fL9+8SR7Tk7f/IFrd+1Jum0xLQiyJgpKb1xMEVcbmI6DiOJL5xnSHXNjQ
dcEHNyIdP7YG1mVorb03PhUFOfi5gL65pkut5NcFtLAAOch6e8dchK6zWxupI4WxwoJDWkkZidoG
xKAiBCdW9BXngWHQSOpcTwR8KCrO2r9fGO51QwXKj/qrqLyqNg4Dw+EZ6T6Hl9YE+dlnbmO5f30D
aCtCd0IFxFKXzvoMAUHXtLkIs9gL9YEnX6+1KWnddkGNfy1hdWO3IRLcvYgcZ1KJ9Ol3hzlnKvlK
fPDlcHFXmnKqnqCd3UFnU/XTZ4OxBoM1v92fK//q/FqYj80Vzj9QIZLPAmk2KaeITh3vKd0JFgir
H/Z8cHveu08YPu0KbW5Xehw2BQHeRBk/sn5DgrjXgI3qm0A0hx/LeO9LbtJ967zTlhIxVTUQVsBh
WmwoYqNThuAl1D0b0EkFAt9m8vX5hVS7ICVgHXn13GvgyCfeEPzrZPPkzJGT2B1DwObwous0fjrR
s0NRIlfx1yFjzkvR6aAkADhwZVWnKbj7JkPijqgWs5RiYBIrCE3qcdp4r47pADLbfWRcL6N/MhpW
PIRbsdUFB87JpJOwb8gAHEIi1TJoK6H+MCId7D7fel8q8eU0NqpPZH0uInVzgVJCfHPpEV/U4BOx
irgXMzoOPFtio7CncGeiv2natfeZdSZ7SSGMa/G/hD5UxItwREbB0nDvGbvAo18qzu4/sXdBr9iT
W9E8lYPJ/qzOgLOp7TuNNyuJFrS5bIgx589S+l21AwBqkVEHJQ3WGw6oVIhqY/KDvi77W2mCyZHm
0sS4M4SBhzxqkwLz0vgv9p/7yd9owu+ghTDaAQZtDoE0dQAdEYsoalYflYWc3E7wVeL4MP9qtfrV
I8QDpjZOa2E/4494GW9bGKTs8gozusCLeyqZPl5ARe0EPBz63gqVdmgKV34hiDLxjLPeVKeAsHzr
zhbONazHnHRQ8wK7CW4ReqfWzr67h1tQYz49iPgSFQX+6sBGA4AWgonaQXz5eOtHlirzZ3UDtKwa
7fzc7XybaWWa/QGR3FmIwSCh+WOQVfZUDvQhhlPwUSBFLk4Dr2tAAW+oMnI5cR8nBIrNHcnrF2yv
5RkaXv/dnUxwS8xDDAlGln7/Ng1HiyVCCxlE7JOqgDof0D+kNUM/02wmV95NT/UxIzYBgs9d/BPg
/Zl8C1SVgoFmHY04WCMVXu6H+kjcpKUspwRCurOMD3fX0O/RpANhPKtZlYmPRgI4cWYgSnDb+2sm
3hy7NEJmVNu08P4ipJf68XSLFtfXEUNIoId4zk/qUAQWUHBHNJ1TS9N7fj07DIHNhfZ7ARamS6lb
n1UoJtvwLCPdc0JCRpc3InLatXbcUJpdBV+5OsfctwZsiMafXIWRDUC/fTqhD5k4dyrl3pAWdtAU
tInlG8ICMtoS5Tikn6uLfht/z2Ot4AJ1gr5Zk5k0Yd4fQcYmp2P3La7i2ix2oDdcJgaRK/SKeSG1
kmhjya1DPXTB9hVNERGnxJjd/9PphcVQwaZrq3tqc5pkA4vzlmMMYLieLKMhmve3c3KtWMA9aATF
UZupLgJAO3Y9oH8AUSAaYD4S3uw3stxoKKPPmqcfUNne5ueKra3nEeWpNV6Pg+OcZl5TyKEKYyls
7pr6Wd2mPwbVfgV9/mdCe/gypK3/sH8naQCXwVzrpxVL5o4ONgaaxcmFjAKYqq3o/fRFxTEwtRAo
v983Xq7qNpgjg17NpkjJmQwmKRE2LCwQkzJXYS0cQLBm8aIt2ZRiCWEZB7+G0OJncl0ibFUGEwFJ
UeN8buBH9Kd5hEAPSn/Uq0r9Qqhx2sxdn3ia0gK1fRoeLarXHjiKcO4wbL8Uo2vod0wf4lijNL7q
Ul6ne//BM1aXFSUWev/2mMwd9MTwiod56HAJr4V6gRZYADDk2RMFgwsDrtilcWPfWXAmxp5BC6/K
zhxKvNw74HkbFyUGPDmLrtBxkLc/6QQlSDfcT4u02CsvhAGhCEUuAweCOXilR/wA42Z7Fd909fYH
XpgePv72xXf5wg/j85f0PNP1Qg2SjpEE+6s2SquUq8WlpFCnauKd7cWRn0UwsyklWyv03+4t5tR/
8+PIGgAqIaCIm3Iz5hy1m9IXeAvUFVb/kkOWKKKxz3gE1PYmEaviZrpwYwS9mj1OGZpQu9EqR65r
++LQ1f2iOT4pErxO42DHyx4TzR2PK/iLSfrkS0SGYEgRMobeR62qo7JQF+LvUQpUy7NZDj/l3RSy
GqfBdwAV1qDEfBkOIro5E3QISQ8v5VPxLgDSfHdRtMrkL71h6Dodo0UFESZVCE2b97/oT/3RwdNY
Tg77LW8/OnPYYavBtKScK/p/PFNK1wG8Vj81Mncwox528Gl3sl16LyyO5Q7tqNfrR1zhc83UcERf
dz+80bgDsVjNftUGhhL/sBj3k7SWNf0rcQyml/jLLEFibFxD261jibfotpL+L99z7qFfYIpiK0t4
fAyzIjdNL+DQHhbtXleVVxVMklFnhER74REu01xOR5Ig+pI4OTbV5xZaN7p/lQ/B1PGM/e2VkOL1
D0rXH0qiceaBBBrTsh7izjXLBgdRTVxXtIeBk9DZzdkZ8/KbKQzdov0Hoeik/hZJQmQLTn8o+Hzn
il2DmzDLmnq2psOmDZP3ypypB+z0CEkT0tFuCiX2DS3XrrzKsamxqWu7Do2FpPklsNAUwAWfoeIH
K5oxL7M5xqUJzcLj2U8ku040yKDMcmSvWhmb+tTdO1Crvu3OQ+IHViMezJmnyKti3TkxeHUYr+5L
zN6NV5wC0IuMBph4B0MGAaVZFk+wml3ThNL5qrpH5hDuMc7wenZizSmXzD336uU0iwtA9S6n/r4D
3c0mcPgrfTDql+az58s0CPIhlNu/qga4DtU27E04m3L1TcAwT0MMelU3qJHFMHJgvQHoyf9MqDSX
gMFy2ei5g8Z4Zg+w6IMqhSaWDjDRY1ndayBNCkAfHoj6Pf37fS0+DT2jGf+wdRmbNoCaPqz8gFqF
pSqKlZ5vCEgq702mKeX7W94LuMLfcRUJKj3tUeGD8WWNrnY2Ygw74VI5lZ6BZwQpxWxCEO7obH44
Xfnbm2kEfGaCuLO+0OuI3qHGRLzZxlqb1+tSLrJzkyHidi860in/jpZRKq+873henmsB49V8sklB
gXQV5YrP9IqAexDGtiA5RXorQH6DDSKNa9u3slz/gMjP2Av8W5gNsbshotr88TRYhJNYeT5hR1l3
wuWty72l37SWyJQGMQgyPGZ1i7CJSonoS6YaomH7wcvXzNP9qJw+KuU1XUreFXRZwZULGUtaXpdl
U5npfPYnq6508hcI9gXhMQPE3KOnCSQXAZWsxQH77QYFwKUyi5y/na1flTFoz7ajPBcL552CY2lz
ac7HyiooQzaGoalw5RYm1UTFeq7eRgsJFNjpDv3KDJi/XSCrQ7qfStKy/1GEN7qSUokT9268yLB0
/Pgt/uRDCtKFClOhRlWKbhNTWYYuIjtn36v48bk7lCyCaGV4KVcTff2OhmKNXXpG7XVxvxo3rMyR
Vh0nv7jNoNWoi/fSHmosBk1vFbS73Ne0F1rzlL7CP1uLY9X+V3ksjztDRk0DhjzrTbWYd5NCnh1K
aJ3QXEG1fSDR7XOzO0V0azcGcKy6IadepPvPYmijC/KC1nDMIeufVfSYviU/0C37zaQfyHwH7Dsp
UrNt8Z3VSPcy5Y72a2LIAdz5fbuirQkmCk+3taa2cBqMi5T5Z7ldZGgF3eDCgeoOaAG6WKUc/cCp
Hh+8o+AxahiHDaaGNO1GwlU+nU94A8C1+Id6IhFk/EiOWDoL22dIeyA4LKadlJZNjsXcAu/2bByg
yVApkumJu/l8U2gKKd/lmtSi6FmmtqrVedPH0dy5t5wZAmG2nvsBMiW+2K6uTKya8D3DAfC6RuEQ
FQ2DYzW3YLrJwb1SwpArboHP7fFHOHIh95Om7B/JsgiFrz1i++9UPud2+84ptnQ/lMAKH3GQy98e
TdfYDy8YG8leGXtZrvgolMft9nLES9klnyRPNUl6qn417dG6iyd/muwnHe8zz06E5ePcAqAxYOat
/QZxpqtWBL0fna7Sge/qF1Q/UJBM1TRzu2IrjfEEISA92wFnKnEzKA6Fk6qnYUwK5pJh0rbtoy/K
bYKKSWRuRCpibGDf7EhBnh1y7ieT4nmVlPZf1idfFPR4b3sUsY8WykLkubBT9hRiKY3s+0B0xpIB
wmL5RL/oD1xwpez4I7zZNNHPT4Tp2kwABowkU5lZwegQS2jWtsOT4gGwsrpFp9oVS6jBvWZsTYvg
y3wHgStXzcYWWmQSXJjj5xhAd6cltd7jMrceDVHaM6bM1batQ6aEOZcDO/cML13coNTUfESW2kJI
JiNmJxVTBHnYDTG3HClVZ5EZqgdIVA0BgaxP2TmEX6gK+eF3zofOJvp5Y9H16eDgcNLgqAdVhD3a
WCyD6y/utYKdG38Pd99nf7n3hu/S8pxj8SnKHo730Du/loiFuAb3fxSKInT6CzlEXx1WlE1zblxN
bVYi+Qv4vYlReMlaPJirNFyGUXRiBIa1lJlVZD3FcPIpXLxQ3DYXGb1EjEi4T0T35MR3lZXvpCC7
IhoKLX+eHmVi7szWlXApTB+8xkPUHiOO36qk+KudNKTQQJX6+2EFH9TPzJYF4z4m52Rg/oRcW3to
nLmM1CBFHirTnK2AMWYkA1sm7vNF7DmB2gYSI8xEhck8y+IKQe7GIhSilD5FZmW13+auCubcEIEa
QDLBibBmIFroP64feVA/3mefZv5KmxpPGitcs/GWkLBBy+oy4n9tn8hktuYrN5qOQ/7KiU5MZCDy
lth1D9TmzFalhwFEN7E0XNZ/W+iot2Qn20gHkrNT0Xly7QOLSQvfyCkPDrioYMYR8/wd+6l816O7
RyHV81tl6P6IzNkzvlFMnR49B1CFm7pjxoIgQgAi5OPTDHCXWnkn/irpKodjCiQWWSLOEnq39RBd
HSU6dIZmY69gqNjBmsjRHKFT4TDdX1ej8cT7tptftToYq+20tvBYAtA6QWkflh263owzGetdnAUk
V9yhe6+Ex920pu6DmKVi1oWYhBChpWmYcbUCTuEIGs79pUaHd7f5bPH5clJtXJuZf00d0cfz0Yjk
+Y/lqAscJpYYQehlfM8OKgtUy/X7qYKC+KO314xE5lD2vPc7QL7ikV/fwfKDsZrWKen6o23sdbwd
AwcDaqT4lYqZFAzUF74OxmELegMZpa52LDlrEKCVE58IboiDqWzyhaa2RnZJuIxa6TU6sKeJPUjF
nvW+ghlQyQQ1HIyA1jeK16s+/alXzLsxasztAYFwGsFf44UDo4jgOO/jSm3rz1pl2phAFmCNKt/9
fqZNSTTT5dvYt6IpRt8SNrMetVw00hw1CyS+4YBB/XCuXiW8ZcoOHzrPwGpQnq5kNqkwq20eLWMA
orWjfjXnKum5pk/tkMYtCGx5NQw6LMF1XyX9T3k+Wb16+wlKFsiXl8KczCQm0bFUYufvvOE4hnFx
vHySVe4KEmETWYXFmtpKiLduqKClkQBoIwGVZysnhauttzOGajOiVHVLVh+hHGjjuU7hV9IZjolt
YAKmoo3vNcgvkgOaVPCNj+mLqU+/DOCaJvoXfOQzmkq28pK2Fu7kPpdgOEBH4iVfHyQ75X06ej4B
ex1jxdnoR1iQr04Bt4N5sCG5v4bkGXyDYQHryZwAfzyaoworZmu6dtbrkw0yOVRHw7An4u1U5vt1
6f2ujh6jb/7+LjNvkli+VLylLSxQ70+eL5yztUVDXR/SOmD8uvtMSmuslqMFOOwrSSGG/BJzbXB4
F43B7fLR0gZuaSiUdGYV4+GgnIhWw1t29/Ri7E+lyiIqNn4BDE64W3s4ImlJaMM15anGxjwXTwBS
KjQitSrAUxSslGegT2wzpqnQIcn3PP536vTmaeoiS0BKEV0qjCNFFzjOnTRmNuNS7N1JkTUs8JgG
N4MKTsSAsic3+HDmZuemKbJiUEiHqI3bo+q7u5iBfLHEfFxvkhBUwPubIY2/bTGmrYRmeMob/iYH
mbNzgwuuol+2765mQQryKssvkL9jGaXJ/rVDFNEhH5vkbu9cIoAdHL+PLDnOpt6BRIVPJ4nLiU7w
xpaoI0dPtmszO4lbp1QXN50HjOT6bbHjcj1vRoy190RWVlQPMMrUo9XUnN2HPGr5D7i/7r0CMmjB
pms3kOdsn7FGAnr4NDUYkwb7mhRfkjpJnpYU9BOa4IvMOxuLGUtAuy+efDpVYcfw5pIfoxJRK4Nd
K0WFJZxm4ENO9Um9/FCLXsV5jvAibafxERSPMnlK3ZUvMgeXoTgJbREWjRZGhnm+RPvgDDMYJk1W
+NyLRqHwFJDwI1O4FqE6xZh7ht+3JvSZ8/2y40K5KGyCc13MYJUTSTnfbUgEfIpfZ300TGNW0uHo
FlyLdJct8XgR/ZD2qle7PsHfDeb8V4eY4bY1OmIQEAK2u9/J6RALPqF58pGE9P0FlrSoiwC0gPnK
FMtKYnu6oh2Z3LIUCL7oZxI7XKMHJHPw48TjpjWS48WTdAZacbrMcX7OLkd4CiumnAnDvKxrwqFu
AGAdWxqOmv6nLYxppjF0czH6cWmqQiGichLWVc2PrfzLdVSSaetkx1lbh1W+OCUSmXACDpmsP2EA
ggoc2kYohwEzIBkcf9DRLHy8KL+0x4mx1YMK4Y0gOnsRR2arbqLI6dHEtzls6lXLpHu7yv3iquqe
hseqQ4TG+ii1C54Riz/O6DbbznpK4F0/vUh3ZC8SESzoPsbXiVQbhAfqGF7DvruZbl5pZJ7fyZq/
h948aDNOSc/srRk7lArxuyfAtq5E+zo1Ib8PGLVzpElQD6BmfoJQ2wIvYdi3XlMVNxoQg3XSzTNz
c/djjjItNQhPVsdtxJvyNn+rj1IRHv1KLxEc8o58o8uwKbkVXSt7a7YTly5DyXR5AhvS2dswFoWC
y5rLyQOY04XY8lXDkEWgYAiuruXzGoM8U5cSQO2GxU1d/PTdzie2Ez8372HwhbqcDsqoZYI0btnp
Ka81w7NYoew+I0s44rvK5I1Rwq8hPJe70mGTiIo8wQL79sY9sbIB13Guxg+70i4pM4gdeMHSLVxR
YZ566Mr/EfVk7JC2Axo5yMTlwuhJzYQbYhaim9YXvwaYdd3W7SF7J7kCNteghgaCGBRshKWBJaJu
FpGw6xhBAfK24zDvVMFo9ng576dTGzXQzTXm94JKSj/dPAJQtKiJzf1o1va6mPsjhnYhvM8YOcxO
l99pbw/1aatBlftKbDFybKlucY6gfY9wlIBzrabLKYkLKtNB3YZbyWG+HquzWR52bzDv9x1NHf/O
QZcZzWcG2qJp60r1DU11EWojjIKcj5wTfENjGdgSv7UGyMBa0wR15Q7j/WLOef3MwnD8vxOUq7AZ
WJPZNY6YZ9e2+/OqOH6vUCHMDWSpP62yXKfVQDJTGl4na94hg70S8OnP3Jx67Jg+rPBhz6F7eIRB
BjfZssqZeW89KhC8+NCU1SvBpaw09IINSByvlbLcxWwXfJTUWAKMTmBse5Gp5HdQxPJJeJCR4AU5
BnI+/oRPsBfbh2NnPim/CR53MiKbYcBANAzTKbjbXJtOefj+47eLnjKXuex4qYiGJhc/zd8X/5u1
LLpqtJt/oF/N6TlJEZiGMkqesIDp/6GFWPVYLWpfgEFxKOmIMvaXM58d1lKFZoTqtv5EB0scZlmx
7gMUeNB+sOMR7b+ipvZ5T19hn7Zw5uzUkc2jlaGrQ223QOPgpdlfRvCQkfdZsrBCndOXUtwdZfCG
QRFjHBbjyzgUPnGz12f/oLkCqRs6o+8pWq9Dp+9oMReF1h/ubRNHC6D2CxrOjyBGZXOofUKudBnN
XyN5PozrhJ5rSQuRlujZGsFidZDXh6sL41hq1+YoK21Ark2djCRmdBCQUYDTdX9Ky4Dk2X3UgEWs
+ZABm/DcUl6RPI2VheUTSVl+XLpgT0QlRx5HlhFu3Ny2UnCjnGhu+w8TZoUc3qLRNSl/Gm4o6XsP
hhQucmZsQyGWmt1meKPtAuKW+xeisnKh539XPpzkIojcoAnprUFRGWk13IG9TJ47KesEXD0T2Cay
KDctVUa5q399hzIl4ew4+3dDR0O5xBCNjtE/B+RXYWGo1NwUMPyEPXsIbzdQRCW29I62zGX7pICV
8YuWo1S46yMAXREJ1CNwaHnjJlVyiYSA5zNRSKZgJKcwb1TGaxk99qaEj2G3tWagQ0Tuq2oYS3vy
dPvsi4BEEuR2ZhVj4GZf+mvmwsuF6zLMf11Zxh0T91C56gScVTA0bGxSP16u5pb7K8Ir+lQK3OOB
b+moJBCEe3QWLaggw5jahFF43fBX1xPJFil6Iq5ZGSgA/ONHoFiyrW5QL2GZjaielRfDhXacv5/Y
Ur5FIung8sZ3g2Iiz4210lSEgb/AWUlaM4gP5r98jE12P/r4xWQXZsx+n+YHjUd/aFqbtRGh91Zq
cLTUrtZwbIvurf8tzd8yufBoIkBXH8bW9fc6Lz1BXBfprljXMHhJd0vsdnRaD0ZsmwwqyuFIUrwS
3KGbg9dzRlrO2PMhqRBOsuvAdn0mqzMB6fjBIZy0aCRvpWsrnrJuoyOrl5SoOTJMkTpMbbGtHq0t
3RhcQBUduXfhlr0eStRCsUSGQNBJH3qIUHjB9PgCsipk6B4NAdv0NTO8ua4h7j3aQuY5YbTZDYCR
0SJDPBcmyiSNXhbIJ5cCDvw0iivp0Ek4XAnmqX9jmIPA3ZX47VBoJS3gnM/Ne+KMfNKIqVw6yIS1
LyMqNXOgHANZmH95CEkXI61syl+XF7gG21JpgqBmCX9sTMueeQ/wKWC6GT7fQ2Na2QFkUF0PjPwX
6tYPEVrSVUduDkghZCg+DsfEmDyxMzN1Ojuv1eDgag2v5hU6XUUNNSqPqJPTS8MhABKol+NDwZQA
Ib7kJJaPRCe1QwGE7AVfcA0yXYnXRZdJT3rE5zWkY6W9a5RRk3+hVkPKcvdduUcpKEzL+8KphBv2
n6QVhwYBh/j1LpbXcXVzvXQTJiGTEJsiH4rA5HSIpFTh1joxhCOrz4rLPemiHDIpA1J8zKlXvZof
B5+AcgrAMPaDthncHuQio+xKjbH9VVlDsgTy/XPA36cnzU3Ok/T4kaMEQpuLYAw4uYo0a4hTEERk
kDxnohAgusUkPk1rhZrccmBTudd4jtAdpsnISPd4+482J3kJsJ7S/j2GAA07D/RTtNTWi9FAov9u
HT33qvUAH+FjcscXvEmypN9AtN5Uy6LGwOZyT4imMd8Rzxf660fOKU4PLtSI0NS6lrNttwSFOFg5
Kw8ybyAmxBNL2McbpOW5v72rJHLmbL5tiWNn7z0oXKsRglE0YJR0JWbF8Kv1Mc5rz/Gt39sHLPoL
nCTXwsIB9754DLRQn1vW8Z9QoTgvWTbeaN9AoVZOgTCzHBXX5Qh/gAp5jINhFWXzwJZq8iQGzk0F
lgJDJGXYbL2J1WPOHK4MW/+rM+TFsT7e2KubXI6coyFw6AgvON3saLvk7rbRZW7qULV2Hc0Utayq
iGDect/ODKoHGd09kdT3or5xOnyX4z/BmngblDxy4mHmrPwCVoyK46Tp6d21xGI3y6N3Xb1Ue5AL
EquJvqllVBxjccN5AMfm8GkPaMKmmGLt+cetqP8RdOpgpW7rGtlFI3Q9B61nPAvh6nWaTvJdxNrE
wRmeucGoNRnkwo9GaF9ZxHgLL1S8xAccrYx2iVxlhAt1VcA82x37vE9v9W0ZKna86u+Mr+JG0E/C
oaCZ4aetqYhLnJi4OXBqiZruqIIR2kksD7mZnJcAYYGLp9kU7tTbh53hXl94f7PidEPvdc1v+Paj
+rTK4QlcmdIf5guZSeI/2k6ZrovTLOKsa4jvMb82wG8lPsLUQv3GJEBFYGIgfzJOxozhkxFI9vwe
gGp+eiSuECqnk7BT6I6IRZXx5NX0NlFggnRYUeW+U5Y+O7KsKhSRBWlQbVezHd+SLlCMAG689fyi
YJdZUYiNfAKZOTmmL9aq/uMvS8RQHUIqdqKrZ6maVhwcMnApR9Miw9wRQZrG53ZanB90Nr4f1PEZ
+49O+4IHnWszydJdd/akI6n5AX47KG2CkDRTcfvIEjT//EpY2t7HH7Nz9xxLcQv0WL/mqiJ3Q9j8
nkwOUWCUuyzOrxxLfU2u7BIDlGDPo0zSy7t1EKP2Fo10nUU6B5nx7eAxwa70kBim62HCxbw4l7Cv
scng0x8sPWAT1GxrZ+vx9nittDwXIar7NWEMKOhA7VHhm5nk9wSZnaCS0MSBo2KWjAEncLJl9SfL
VrovvfudSoHM73LQvWSjbzsyAHMUCM13rv9G1kUucICSo3DEbvnhi/fatDITjCFl6M72Ij5Hkrmx
BM7P6Ku3yHJu7nfHQSLFra1rQyHxx3GlJ6kElckVSWVttZ48Vce9PPzecR1qzJVxrVT/ooI57W0+
cEh1yNToxd1ZU+xk8rtewkuFLgOgoNA9n5bTHggDKe08yS6Da1/eNZ24mqfvsLxLk96ls79uyFUZ
hktMNvYidgHq0cQj6nri2W3ShF1M10PjybYTGgwVg9kUznzxinrkRwimy211oMDLeSMg/efv4lmV
23LT6NwKiKmvsCTK4ebAKolumNAYFp0dXXK3POz8JMO9fnYrCAMg4OVqlg59S30hOEvitQWOaNf+
MvZXy5zrbvNKmzlqe5Va+q2o/ZEVDqd3lLzQSDl/Y00yBsO9X72CM4OlmJ2UbD3U4GPMLCDRSnV9
8CRChguhlqa8YxgJBqYPiFdmgTHhwtCE7jo4xztwheuXjB0kxDC2cJpJPrbtgZmqoGlGniCCBzyM
kW1SljKvl3B5jca1oBccO0IQSKwATFLV3BKhKwH5eAW3VN0HmlERmHt3Uje0zchBRdX2JcinWWNS
ln/2mYndpuHmexE3PAy5AgHbEfZR8PLmTyhISvpzCI3lniAwdKnr4+kSAg8k6QG0TrsbDXbIE97f
OSi260TIoqzPlVFxm5YgTu1xw/LoFfFHpCUAZmBMkzj+LZHj/8pHdfBXBlxXzxmmJOAxaD7B+hQZ
NjbTRBZo/ARzcnNVPhZ/Jz5C37c/g05by3jl0fyiCjLfyFVDZy2OQzjdcMJaM8iShHDf9HqMrQ3p
ee9jT++kaNlxcIwv7B0k9fLpPCK4/+kehFYsuSYQHYxO/ESb8CjD3x749jtJJrFWc7ySsH3BjrZ/
vja4Ruwzl4IZuIAXJpTATt11CFkWo3J2wY1IM9I5tTaRgiQXxzSYmC99szaaj7vtJjgcxrVIuWpQ
VBoHcA4b+b4kPKs3CV7lAvNCt6GW+cMV8phydLt1guEIpan2YfVZSDu+03U5SyVlc/E4bvNneGmJ
jDaovEcqVI2r3WboFXoO6LLscyD2k2RoQsuhY3dEuRL1CegzAq51HixmSDBi7FY7RjI7kSxKnFfz
4e9eDDmBP1vf9XPFY6pJYuuVpFtcMfYqUSS1wCFna6r5HGSFqTfSOFgFC4IVzOttXGreHEicp+Tc
wgJ5/+D/Imk5Hy2dKkcEoUIBPDUkxWXQQUmLj7F4qD6gxKft2n7pCwdy6riFj4XY07cC9dcFfiZy
7TNPnqhSbYdxfacVY/CxaTeN3tT3RnYpBQP2t0xEe7cURLR/N7nagEvZTQVOeIEFJV2jJ3QqNt6a
AEnqAy0oCMAMhzsCC9zdNpQi4Tm/75TuNYaQ4XrRJGttm/5FI1kWg3DtRhg+GZfy7AtXBADYudYo
IXZSo0f9tJ7gVOVoxJcYLTXTvRkgcRe5ez2T9/LxaOszV8NAdHFEsLKIv3dGDylGZv8lGP3T0o3O
O52J9doTn8lhXAOJJt6l7MhmnjUjaKJNx5bZocIFtQEQp1zN5gvgzKQzk66H9FQ7uVcVKlpjjRPd
vG8Y89KUm5UZ1SwvRBybId9y9XkzUHO1MbfqvSMN2ytoQGfjHwqAkS/W/3Ara9JCgnLINvvDEXYw
xnExrMOaPyz82BHk+0dxDIvEwALUA2Fyze5p3yPKVsf5L3+xmObM+TAvM/dp/KWcDK0yJkUMgQx0
djN+Fr/n6QVbxJWEbTu7053lveBFQLdNhmHJmE0ionhDHDdMoHMkFuh8kYB4eiWO6twYXMmEpmGX
ZKkikjhYN8/Qk0qbg6wae+5STvIfvz1gQ1DjM+Q/epXzPeSOQGXK019lZWr4Ef8dtOYPiczQjLyU
VXHEcCIhpl9qjURMxA2IB33z5ZKKqcWVAf06gOj5RSDNty2/OtTQBXqsWcbrT0HCSIbVCFqqN7Oh
9asVQZ2xH7/SdZaFZBlEVm146B7OluHp8+M1/sxneu1vGHgXM1TeqhOmkQAH/eXyeEfm71k6T8ug
qd4QMAdUJJS0dKOd7E8KpYVcqZAbZ275bqctXi29CMZjPC1uxyQdeq1P6jDJJ/t25XTIuH146lDQ
7q2zBWcT6JSC6n6SSYidCJLsmc1MNuXU0zULOKYuAY/GRh8pwyLLcSIhBgc6uqvnS3ozjiZJvgpZ
3CAXJX54QPwAUMjAXUN8+uLQgpo4VVC0SPVxV5LvBgZ+D3TS+1VsGkteVfDqfNCENQyBGz8+0oWk
mBVw8vPI/YH3S1LOaGIiwETZsj785etSFxUcyODE5RwOHykIDDVUZbK5GhbRQHebTQPBYfn3L9ac
3S5c9PxcugwSq50tV+nCszsxlQYNjxkR+i2FXBgSIIqYFP6VfgVU5EQCvPK6VRojUw6yxhwyK8Y/
MO/He7sFYzNbXw/GxzCwOWCmuPadvksN02bqmASkrEx2H+pOeWuVNDA/8XCV54QnQiEARXSNn5+V
5sCpvu6W22KCFIwcAMIssLiESx2SVo6o7vTM2qnGL8BEO/u63NMhVJJU40TyJ275h4kekTzCxRmk
J7JwlbHV1mSVORrq0CUuESnrlkeF0cjh1n+9ewWe+O3/9Akl/jiLJnkm//04fh7j5G9hPwgwGLQX
R2NZ5l3c7CRQ2RvUrluZeiY/X2TUKmVI2iCMzu4h1YhffF8yEy5vUFwTC0geW0fsYgyQuOoUDwr+
adqXliz50xq9MUokGbLuJ+pFgEgIdVrXOPSABaqNz6sM1Pns7zT9C4hWiwZrG9K72o+O2ZWsdItY
f10PVoKdzxl44Y/cR/aqWMLz06O74f+Wify9C5akLQzZdMpUoYYEmBHVomSeQPv1kc0yhB+qNsx4
s8oGwxGKfObM2zF/Qe7gK1B5ovoY4voSO22Nf4ow2mi2LaMNL0hK3U0Zp3eCm5xof9nQ5yuqW+Fb
fW7dz0zVToksjeuQ6pz+DoZ68DJa0BQzt5bolQ85I4CAj7ubm74L4ayzatnOnCJmMFdfpYu6yNHU
DhAyiOA+3gF1XLwzHL88RtJf7Zz7bE/o6O7M0NdHRx0RiAp+gMAfg0gWE1RtP+2ywS3e3xwUde90
axytwOUZMwIPWMQnF3qqA7UkMn9DWj9ezy2n4YAPB/gu3dyP7ZLPv0Jyy+hgqjcC9VQ/swkr5zBf
OPMNXrm6Bqm/+xg3jvU5q2myZb+fSoT23y6cu6eBd+g/broVEFcIIgHMfSlT9sc7KXHZlYYFI3bi
oIZtPVH06M8AEMCmrjgOi8a2N58wiJ2DPX5dgm/KgdFZ5TsP6EPUb3HaDdoX+uLB2wfkiV6vmdj2
IHJ9ZNTNImTLWISPqLluMASqXebn5ZrzurYwjNCo7SyTKNqANxfYlyOLypZseOeOY1XVNDB+oHY6
HTRaqiN9pCu19Vr+aLQMCca8CSHA9vaTgTkS1zXXMzw6bntKeH+9nUqJjsfE6MAKwfccIfOvh+a6
qMj3MPDpku4ByjCu+uoxlz/1FTuTXNAx0fpVyKtWcela54w56D9BCivcNg6YUe2gZyNKIpOkqkhf
qfISXlw3UaxCmTZG9khsZ3YM8EMv/EkhS/aM+Xgmeb5LsezqLZ1AEd7wMYNfhzxEHt/lNo2nFXXI
yOhZ5hihF3t5ht2OlJn88W7N//RFSgbZbjvwT6SdKVlrDcvPt8OmoRjhp0xVEUILA7ZBB03YEDio
nvhtzFsCi96igrvo0dzrJP1v6bnyrFy9ws2xy+s97tVmj4Gkv6hURCQJm+ziXrADVJLbigUKVmLX
XZkYLAYtaPSVdl6V2DJZl/KKRNOvERffA46r06orYYWOdbuaG0Mz3LdqzYin3PyD7YqO/pARfxRS
4uPTPT64WHbi4+6AY512XVj1E3ODRM1h+O3FtiWP0cU5AJXLQNMmS/k8w7NtoLkbor4/DobN4OLd
75A8nObyBEBQjnoWvezAHW4lpS50dxPYhVJwQihJDHfoHfT+KtI9T8vf3nEOplopwe1l/tUB2Xz2
qyex4+GWVBTdQfiQm1YtNUAOKu1WE5BHolJGS3ScIeEN9TZSbFTJIyCUcWrj2fDidkO8PiKNlhiT
H17R7XhY8j+BSsXei96AvSHNf7+2KEW3xRW+WoPnnxR5m/B10xaW+8WpxhDQD7b9omcVC9vMl01B
FeRjzXkzF+5Sq7AyBHjFzdXdrj1nEFzRqDfJtAwBbjG6/MS4ByVHwEoOV9TfAK4yFb0ZuQBlRE5c
2p+BQwKutO9RHHm/fCTAPi5Oh7U2za/w5o+rDP4XNUZ/waZCClhznVy4CcFabTRQhlazzJIwC2a4
e8P2nVyrvxxgfW/Yb2YRaLbswcirylspYNGTex47z98f3V1yvNSOqsxgGb/WS81tf7IXQckdJCYw
XF59BefRy1h7xUoMzAiFVu1RUxs9Aee9a9qZ+a7oLY5PsKNjOYslrLTMxxbohGqmtoiFG6MyFJs/
t3pZw1bekepiEQa7W4lRi91cH4ZHYGq79iu1SjaRo+OaPOfq1s5AI18BE9QUGmrPEgiTSUVw72Qg
0RtvE58Kc/sYsOqJFdhf/2rkZsnecnQBNzJYPZKP7nVHWBWh9Iqp69B3JT3KfaZRHrV6w5KLAXEY
wQc3ZrSDoM82JYzBPxAeA7p+4DZE3SxFB6Nzx/nl8o6BDSusK+tF9304tZbfeBFNh5aiw1bopay4
xOsEloVUtvNoHXezojqlHLd1sTr99gGsl1tV0uZEJ9sMmAbjPfFyZ7Qm6orDHDzjwFH6hohL+BbV
aYcXZa6YGwiVOB0NbnolCOMAkeuzAi6kk8r4ZqRnvgC0DXsob9zVK6SrOvhqZD8JsbuStD9Eu1iy
2820aHG96mWB1Fr1h+jjIaMsdwaw3lttHnbCpgobdcPC2yWYn5CT56VADZ8NmdJ4GpICv0ybNR9w
PPiAzFUqwC7SqoncZ53lN0uy2CFWZuM5Ag1pbhWnZHWYwo0I5LfZ1Fp/QADQy07kFz0vNhEomhM0
cQu1WuIUqpXA1Eq/eYNm802+h00xyD6W1mR3s5ZRgF6G9iYvDFMmdsVzIIdc6JCAwkOdfrcERt7y
HLdskxkvmLUUX9TF06BEpST2PyQ5UDp6DJoT0qIgE0pg+kVmYtv2gI947PWV1gAaYRAvOfuT9mX0
XG78d0WxNpYSNIhbJYiBAUk+tKlh9Ng8TpX82rYvPR/6V2ynI+KVhZZ7Uj/Sr+/DVXdn0fRSofy1
75TiEWyPhROTTpGD0gslpAj7SP3yZ66AxZz3m9mpaTwIjScHG1tISlszufov9ru/zuiGHtidxSHs
XRZOnlJD7IZQt6QAp88ULLXwJQDTf6exrP2hq4lnhTmTwMh9noapUXF8KO3YcGuDpQxpxV7oG9ku
r6eXdzq4qKwLVrOB0ArVyyqNTqe9dQ7/NRqqjfUUu4Xfzr1bhDj4mAb4OlFlw2XPf2zLMkHxdnWW
aVDwnRPMk2mOYO3ebDEE1y55FJ+Tiy08D0nbaipw0x3raiPF8fyDXPKHVeDgKPXunIhjIv1Zav1y
TC6diK4wct09R0LpfBv09qIkR7+9tBp0KlbxA4CxBQzOKFum7zP+PXaN/3TEC1S/RPG/QQU19o5b
fAhO3rbfM92u6tbvXBV8keCu8w1dv/CF3TwRJuEDB7wsFWOFV+VqzQf97h5Q2t8wv77lC0ZpRPxj
A6iifz+Lca4yNuGz3TCDF/RzrEa0GRY1JtrxZl8/HQvCRFm0c/Nm7igU4SH4CtvgrD48AyGDiw5n
RxV9SLZeIuZS1QR7UoT5aQGbrvoViWWgEtCXV4s1HZpsRF5+OEQtthYi0rkhniQCO9By4HvACmoc
ep4A+dXPiGUP59CHaBvud87IxBJ9KmmV07JMknae5Pp7Y569ph8zKY+UOoOokBOQeN8lQ9cs5DOJ
WBmMEo4gvZpPKrHoKNXMYhMNLSczVjfP2lru9yS7F7w1iPg3RiIuYVXkn3pbhEsPjwxA12LkKX/D
civiK/b7z1ysHKY+PgUaPCg+Z8Qe5G+5gNN6XLYQVOslvoU8D1cniBAqLG9K5dQIjIGEyGokgTLS
KO3sOBNKYnX+Jt+T6FYqbSXRymeLChOR2hJY40qly1tC4/R3xyU/j35ukfTtYe6HLuUHQF8zB36c
At88JknnWPgCB1UQwJlwDr4FfaFO54THHZFPGUPJXV2iwIOvfroiEbp0k1IGY4olxaMji2QFAW9Z
4KQZvw/IFvZ50KarTQsJsyRhdYAtUIlz2L2TX9Eh1RlBCQ9U0tnMNWHvqd6l7PDcKcy09xTJUA8q
xsXy8PJ2aJ06N/Dooa7fiGx2V55X9aibAVHdNvfGNqR0t/da8NVJtFEtrbRJbD4U9cwcPlyx6gyH
hHgzxd93DEgdUl/xjISG/SoMVJRNggEhZbUXxQ6td8l9KA5/3TDsxl2FYoVxhGwwDijAWxZmj9RE
W4rTNk8qJvbkG/T0YdiDUndt3zMsCpodnvct15H4m074kIkEbsLUwe7VvC7KTSkNzw67sE/kn4+N
9tiUjKLnn57b460QZrI25QL0/JWgXjnj0cgyR5RNOdt10n0ZzFxbL/nnVSzSRdMUfo05eMzpJNGR
y1oYQzCJUr388XdZ1sEczht/L8B+jdxfFwMVs6R/KPiN5UJd3BF6M3mm2XQCgjD+diClHynaVrJZ
+gJI5U0iiXjeWTpNLEpMcWOQcD1y+i1yGFap+v/BOg2BruRFxxxQXvINQyCc/c4+L/lBict64END
fLpJYXGgkCifLPunLhdsWmWxWlaVcqvc/9KCkiTlH2YovB46zoZU7nb+c2x8qj/W5gYyPyE2pEfG
u+WPJrwZg9asBJkZN4UlZMrEe/MI3APHBMF+0Wj0jveDmSGc4U+5bmK6CMWNbKeVi9JWz6PoeSo3
KBE1NhFIIpoz2ccmnMwuIYCK3u8rZkAACaeAHO/K3+6hgoxrVnHdrJceQks82t3QvxCdyzdWDuCv
5nEkQ8tSeriwTWAjrU79G0FdeYc5pyoWbr5FbZ4QeO1xp9SJ0L8CE+P5sUxwAueiA4bawPKvwe7J
ps3Ij5ACYTXxJ4CXfI944+63/QvlTTT9F51qk78B7EWovio17NfDY07f5Nzo/PpJHc3cOw7mo/FK
Sdf2CBNANtqr1KVr+Oo7LWqPRL3UuwmFRkPOshyC/25NLtrXN3kStzGdBVSNeZKRD7RxdflTALSn
iGJtWTBfZwA0sacOP5aA5P20g7QVvW5zf5beK7AVUilGOcjiEpXDATYgUPI3XYsAh4XrKvS22UDQ
PxFEL5X132Aw5vLcRn2SRQr6s+BLMBXc0K4nlpBZPCleIJl5culeLiXRJ89pGbQnCazxuPuL6W0O
qSqV2bC06WbOUZ6owiPwPpzTaKvBbnZn4KkIDyJyT2bZCLyiL4PxyU3TlKPWd4iXICwLGOo2npl9
019jLQBxYqJiDBbFcTDbhtJ1l9gcSQY0Uj4G5KE2Bfxa2k3+kq//hbQGDP5wZGR/aWlkzRqS9Kzw
r4xrIY2zRsHeeVFqlkb85NMLbXTmffRqtgj5gJIJqWbazRFsWUsqBuGay/Uuymfx8SLZiKN/X62A
ttzdnmGb5iHRG1I90MSYki74k4NV6iA2D30NGSgvjZ66NWJthozUx+8oNX+cKyHIfTjJ5pZ6F9GU
1NpTxvqbDK9TTOWk6MeTnY+6pdT5qm6xuGm9P0RU0gnXUOtv6GHsABDlqrOiHr2n6EnHpsNDX3p8
wCdevSRODjQhOmwRVDacKd0Db3rE+xyfkFnTc3ZANewvycWcgoGrTUysv7J3vuVBvgR5TZGRokNo
svPMMLREkQVvJfenOAMTiDN4R4NzDWTBNUiB49BYnKppILO6AsK+cUctKE3f8Oy85eQCzl0W04cH
38DikxKvxi7DRVg+VEMO6V5L9G92qNELfJE/VCVoSUBd5I//tLQfZ81Pgw1oB2dyoqM1t4jivPjb
p6fZbxBvsduJYjENjeTX27ZlJex156Yv5uxZ/XWH4QsM53+Q/4IGuXdZHmo/7A85K2d7gKKSCy0r
ARpr7oHE2/xUkB2RUDwOVcm44VYbPj0kJTmz5rbExZEG1Ita1gAEditu1mQfWVBtNZz7wfyMno7r
TJgyioDOv0xPalgzeDuOSW7gtoPpgOc2BcKSmwg3if+6QmS9y77cE2p1w6YG5dsVFhQon/2+Zlco
MrsOvaRzxiy5eq90/nzNKNtcu04g6EEhElFvUHC7lyTFWqpCLcjKJRfALPut2igp8rtds3lRdFBE
BmYIj9e0XnRFUJE1exP/5Sa6gRup3PHpl/E22aEK4Mfq5Fo4PYKwpWJ0GlO7EJzCs6P421y+q0wq
1PUIHeboK2lKjgubeb73L/M0SOp27NwhjgB0zHIv34eyhsFEyF8ogEJgnNRLxLoO5SIhdZfIFlB6
5l668kMk/a4lf7MHlLvdLkF5FGwmGVrrO6oSnhGVkOJhEwIYRyaROHOy6YyX8+tiMCS0N56GPDad
LH67/EC6MzjgkxUZtry2fFv5F2ZUcuwno1dKq8lVYiHCHW1Tf98Fsh8dFoylQG9GUShns3fqcKLh
Yse9yo6OTL6yYhjv04ThWxi1e5oehM97OOA/zIa9aiykcDmS84n7iEWwVs3kny+Op3hOpMabiH2J
WxZFLPpo/hAROlSVD66ocSirPIOEcpmJieSEggJa+FKACirthGZ1v0JYu3yBpGMk6/HKXHMNONyG
Bl1QzwF7rtNj+54mqjCj3C2+Anc+pa1jpHnwWxwlfLJhhO/MrVEOliO06tRU1684hqL88zM9fNN2
8rUWVpFQuKBZig/Xc7PKgKD/HGTjD0E9tjP6l9mOZ94Bx71XJdGIX2bpc2pUfad+t/Luzod+o96c
4fI9/7ea6kquLO7RXQO9dW17BTLZTYMafCpmELFxCRb/mIxBYuDjzBHPjl0nhiRA5eaf8opSjz3y
jkIOijFTxFY5BKVFgR+jDml5kyoi9UXbR0DwDqOR06ofshqMBktqX+vq3tnuXwS5XhMyBd0CYF4d
3axL3Jagk4FBvYC3wUmP5/kFlaxlL2xE1330asOtyeNdC8ztm/IoC2eDJD3HqtaX8sHL2QHya06P
fsEI2U9Q3pxjrOpWo7kSnnsjTqJRUdWKAxmrq7nnXWP2or9Je7nFtVbPK376W97wE1ouBj+xPP2m
fOuxnFnblqpvaTqblflJBtmgFeeY7JRDpqL1I7wyaLsUMHApc3+X4ymUIaqPOO+qNDKCqz8jlPig
7u/NWUQNgidp+x2KPNo93TBC72McXMISRrE0BE80+8joDHCzxYHHXzkeZzmOxodL8LwVMqeTW9OZ
hfyLGImqCftgXDh4PmkJCVsRTdWpKumRVFM6+c3xis1jIu1cCxzGUfV8EzXnSVf3xIjGOI/8dZ14
pTiR+9qHi7obb6Yf1GyRoTKLIdVCOczdEFx27COzNz6btLCiKZ5un2V1ECcPR/KYCI5KTe9RJanD
m3WpneDW6rU3XXS1uaOkgumY3f4Thgx6LTKybId6rarlrqrGpanW/P5SeR0xiZlqGJD4chlGGJYn
ePY6FM4VY2mhemFkA+nqOAh81f2mtSrTZwobKwLBIZEYrcubctegBVHSVoOvCWUJid+e0aSGh611
1XuDrFwiyP0fNCMTR73g9nq3GjivwMtWPjMRYQp/UgLhfmNqI+h0VKR6jLSTXA7wqLQ5bgNs0wc4
JM0i+WjoZOTZxEEJNdThB2xAdnUY4jByOsqrreQ5bG37xk8+edcINzkqC8aSjFXywU7Ho1dn1VO5
ueTWghxLT83PGBxmBxetA76w7xFi0HGKC97+mVunUyzEA31dt30/VteQgXOyhv8jJRNiL0OSZFcl
KCqhvH2icp9oZPFBXIAF7il5AuqphXGf+0dvjTPztdCEwg5cfRiOZAEgTI75rsMx4MIs1I/c9SFU
zuwSoaQ9GAk9FMnc8pcuNjMj4wShfyvnXe92R0JIr+ap9tYN4C5TvwHxTJdb54mNxRs5CEdqP2H7
UUldTBd256VxZCx6jQE+h19jlXGFua2LY5hSQGsbP/kESptwrQDnH7Dw9cv4VxoDKlP9HvetPcXp
T88JhdZY1+jlwnX6gUFsWjC8s82Mk9seEHk7QcBdRll8vzwLHeIgkfYOmbBKuL0RFSP0itlJud+a
fOfi4plhFai1nqbY8qGQ7sJB8RkJi75R4nVW6UVZ9tSCt4lInSLrbVdkmmlvzdaJC67y/wfXu6xr
sSVRbyf5O8v8Kjymgznf/6y/A/0V9qd/EIYxJkjGxNqmFqGATFl6eGUJmKWcNnLGX2mpZ9H+CPp+
0GOr9ZOQwGAQ8bGgTUdwPORegVfM9O3CuBBR/sTDZvlkVzBS0to9HWtpF9uJMgTPXMa1ObkIafgA
001aCNclT9LEfbtXALNZI5HbNZjr2s9QEjW2ccQ77mnZlx4Ve1cLVYaKSFWA7HH0vZ/2m+lCeNf/
NnVwbGI4NLY1B9QAnvlYQ8RPuIoNAY0msJHz5m3sP3quDUjExZwXHsW6JebaGGZyualhEa4K5HWt
vyn3qHcDHb+mLndqzhAFG33z7Z4oJ5yTUqv7hf7YmmdsICiheU3Dt30MmwHfiuzKGG2abe1a9gSe
7Myh7EQxzuZHYEZ/krbz05rhblBXnKDRplJEWqGi9v0yOGzqnghdqCuMnOvpfU24r1aL2ubOFtFP
qYDRt5GMseMjZv/lPWM0DxHwZnG7gRjMVC3fppNq/YiX5fetTPmH+nUta3kR+k5g4tMH0wV8JdeQ
396Ir6NtLXVg+JzPwdHShjcHjfNqQkM3O/1vHO7TUI2U0Uj7yOzpoYV8yoaMsk7WYcwssGqihG+g
t8aiWykeIaHpCO0/idrirJfXPll4zNl8T8kaIV6/tkmkT41NeZi1Ly05/mzoKiQh1K1jiS2vd6Y6
P7ypnmsQHhaCWnYgtPCWdOzX5o541InrnPME7RW2Qs4RMdPExDFatFW6ARGFea0pkZjJUyNUpddD
tkuNQu/sjSJTrmGAk+l2bOImVhPpKSig2yzdVBOCRNqioxJtg/Wh57BBBhREPxDv5evYYuOL3Ugg
9sia85n34o7v+3QmrvUmIxrTegXkdAYYMUq6MFAO/vnpP1YoiSbVa06XGkJQfwj6fni9JP8OuBcY
jJYR3kWh9QJ0thrFnz16EJemUuL179r3ndLJt1vv8kcYW/s/1OvfAJRd0u/3TwO/jdLK9iyAm0lS
Djiu09TSxvD7uRAxxjR2+fdi7i+R/q2EFYgM28lGu60AIO23x0nXzO0ut7pMyHkwILnAvUc44B5U
SpGlIvgv0bZfMV035a5nQHvTKr9/eJefRAMLPYFCqvVGzwF3WSg8W65zqz+4T86XJftfwq54vCKc
BBPaEI9T9KloDACtzByv3S2hHPr7ZTeg2lC/zxmyH7mbSj3qlJMCo6H0tuLwbM/oa7waNVfooqsp
E6ImjB8dXpHtoJHKQebqYPvKNBrgKu9WfSABssurzgZtph5GAvrkGLkBUnD0x9STPKRdK6PNXFGk
YcuCkLf8UFY3lm07OtB4GJP7sUZT6JwCRcrdkgwTKXtUjU5bsc6GddSi9DE82Ce+anQAVcg5UGC6
0RoaAm71NKoKKUe/3k5d4DYTrczoTdpjmqWp9ECAaAESGfOnWTf7PJmN4bfs5y4Yp6FBGPrmodGK
tCUyUoEFSYa06021yu75q1qGPYQm+k67dcMxbECDTSKqQIMbjJkBLqiWPKyHoBelmR0UnH6nt5US
xyHYIXDqPDwhEuFD42b/eA/GMYv65pLnL8vInamyUFqbDMPsk1DCDp6a52sxRk1rRXCOugvTfRvR
cncj9xfv17r2aMpFCl9imWgQ73oD8HFuxyGPhx0DlFCZJTwEhspP3/wKDHbfqtmuPFL5ckNqSTjz
uzYA46ZEzbr7Si89j79/lt1ZY3oScTxDQWaJLaHZCLs6u5zA1mQ225gXAKQplaOSn4OCCFRjbuRt
D2j2Gnfd5TpBRyWy9q1sKCobTV5zy/mz4s59aHasRYRm6e4H5Za0kf1sYXLjM4dAEY3q7x9F3ytk
1Fw+4Xy6uNyVUt4kXED+KE6mGP6DSF7Gnq+i/jN9yGWsWhQKoO5JPe/hDQoprUkcN+Ts50mRBf4/
ZMnjc6TGpXvb5XTKMwKlUrkboFRTXlvcb9/qi74aUDPaN58PqCYxSJD8FyCKe8DsxeDH/Qw9q0fW
63q7FfHy8mhY3xtV3RP82rQukzACAAUcZyqNmehzfNmsO8osLnmKAqJo5Gl6NCpp7u4mHIjyS6N2
8pd3g/NACkmF4VH6SPx+31wTYKiH7DWGLnGqQm8jQcLTDRD3q5XiUct005/aEZpFwAQb849vwjFI
lqJQUGM22kWWTs2qJXGLsYCjWMiti/o4uo2MjbDz/2cxwwXaAgu6OneiEcndhI2/uQ3t2bfSIWRA
iFxb8f7y+2/2fcQ1X7sggmomn0BAabW0UsMHltOCfPMxWhzj+MKniiPhzNMCZkzA+ghwdoDbevSQ
d9mRGa2QUSw//KsgUybKbPZE3wl6rxgrIYFQ7WeKw456V+6cK5KKAOUlMQZ2pi7QTfiYikqDyOyG
iiilmvgXDM0CspsYzSwNJY1YzsviqkBvHOPqpPYVooc7s83IpDDgwkXSmBCuoVUA89l76Vx6Bbpz
H7WhL25uvVmhXM6z+KEKGYxxx9YE48zYp9yTaJon4AJhucR0507Ihk/P/ncyexj4dMG0IaPWbLWT
ug0gmZSBl3rOlg+S/+afroq36HgYd4YMRHCNe7abGeuoPqzC2iMxRqyZ1S8oG11/dXImBX3A6Wuu
9D7TNAijymszBa15IiJLbr2P2xLZzaWD955iox7kXokmIMF08YhLakXNS6z9TUeswhsAlqDsumOu
0aN+sBcdMs5Se0+CBNgcdEmUD+Tfq6lsGeXD59Hc2LbJoQSvqLHv9h/Z5kR8dsaulcJKxBleDOMK
ljGqBWE626hE4wjRBT3TUQmPNxFzSsxd3SCqSXwy4Rv/MPDYso/JAgcoXAXNH0BmhONhownv3qXz
26h4xW0LU8fcxsc8BTfUIrXRCZNAwD2igBla84QBxRyo+/JbpMTfe2E3lxJTRjrVRexNyqYZZehZ
JHBrB1ziBYH/N2yogtZa8owy9bTFbrYUU0CfPrXKl6N90bsaUqx3/k2ZxCsPqymr1c2sxeo8K83x
8vqNrCOKGGGBqEWvl9X8BktrHtLEcDQw7IDZx64RZSxuKOH8/tTuYZZSFddVXJC27VqHR9doyF6D
XUEGwaiRJelj8M3ckv9yzkpjg3QHRw0nPboBqTgSbqKQS58vWY01x3HzpLMhqB9g8HWNTzG5UqgC
s34uKybKwsJtH+4WDTimm+VhQcnQxzQgbUKsI3QoxILWfYmTpTY2HgXCJuQnWzSZb8RH1qNnHgVq
EM7HgKsAKsYrcVHTT7k34p80NICbEmVks6MIluZ7p/UoglyYUgAxAZXj5gTNRR626QiWJvUnhrXw
SESQCzs+0Qa1DpqK4PkyncluBnG6gVvVQGzZHrsO0P0EENjgsKEt03tfjyr5ToSLOO9HGOcTlv7g
3/bgcGo8x0F00HROIW41PWPXMCSjytrgkAxJI+38wJiNh932jetQzzy1ttMnEsElDgsobMO/N/T1
bdYVueaUSlYpRIVonsjeH+A0aoqi4kUphbF/JBS5jWO+HC5mRqpeXH/T/KiFp8WpteVKlUP+VzBS
MFlOHsTtCLE7W7UJv8MBzA06utNtpc78tGGX9NwSTXoSAzUcTGpGbNTT+ST0wFL7J8m6IjBVodK2
hM+eMZBVkBFbTii3OWCL22gdPf3RoxNBOOOBI3F5lOV6J8Fx8TJ5sK7mOMC57rC+T9UvNygSNTPP
MBYTBmgnS9w3aAmhMq4QI+frVTUFxlbO/QeUYFpQfJsvVZiwSwo+md2CHFYVm6zVbDA/xDUe+umc
ZJCZiUSfHzD9vQPvOeUv0X6tDhlqvLlHkZptMdNGb/JgS4aSd7i9suYtl4BmFwi66a5ZkUNyohqI
Z5scJ42yyK7RVV1u0+hO6MnPA52UbRLYXDtQvW/kwCDg24hU1BEOTheEa9uTJsN+5o0uImJQkzdH
6pO+VFraB/UAxZGTTSLGk3COL5MEJRHozacLdNFhFl7wrDsPaBqr9cRXMGknmM4lW8F/7QukylvH
AESfajVlzHB2zL+MvBmSgCIKdTmTZM1kKkz6oj0DGmy2kcHjwchJURcI/7R5Dd1lxxPgYnF3XXJa
DC9WJsTvjZ8W/Z2YZawwpe+7uAfuNfil2ap/vdMuyAcLN3xxclM0c52GSW8Psi0So70mpB+uTYh0
Zt7+bgRChGt45XWHs4n7mBOkg/A1zowsQTx8cnHiSM9vUosIUCxGEAjELcUqB2slOVe295gA3stF
fkaMvipnIthRlEyKHYPQW75nGnbVPC5O1d++2RZCE2Ndfl2Ppd1EkQssSAD3Ps5g7gZHEZFVbzf6
lf8Say87RtenynoyDrZKVC1WiRvtE+obBZtmcn8tjxRxgvc/eDvgO+RtVzqEf7MyA9bqGxPhOWG7
NR2ovLiySxVJk5dqC2Lgl/fItBzBVeGVvx6tAoY79Kscrl8spnoOMe+cTBD8r47YtYgPtDpCfnp9
OKrwE+X37Fs5EyUYSNuBeVMg9nFdJHUne1D4LHU12ArnLBIu4x5FSA8CSpGcY8Co5yp7jnnGE/2i
Mnyn+wJQrJ8+WfRSXaud2xYOVMs7LSmDgSHEUrt9gnPTpXDGlqnD0+TdH2zWp9gYEo2Cggsz4KCR
g7/Z1OyC7vxCOjeGZPVXvAEwjioV6l1Cyeiq9xGYc3aORiAdmA8bbROOyl0ajvJ9FDR6FZWa2EZA
IFYw8kC06m4kdoVnE6Nk8s3N6Vp5sfrQ7mXYIWPF545lqA7lZGqpbERpiikw8VvgOUDdaODTm1oD
R6sL4k16aqnvOVutFroKKb3qzz6TFjEn7ze8u5GweJrfvogXfHfHexRd2WMsXG0ZBIpCAIKI6Cgu
jWn75T+N/z6eEIGvMEXE6Zh+VepPgmiisGGNC/88yq3rR7kYUgtibUIGimFdDhboZL/EPZqiYw9x
NivXryX5gHXwjs9AE+Joy5pxPnRoiWx9pnnNSXqrjBkoo+2GbOZdqchs/W78Y4ML/6Ar1Et0uwKm
qvaOwPUkr/I8XWAjuDN9dLit1pIgep2ZJ/dp8sZ5q+/KAN5+Mj+hL3AQO2QdxBwnPz52nA2NXLfz
K85byf/9Z0qlF5TPu6LcAkhQp/nLDsijTbDXF923btzz6ejMOzfWHcybFVuTwaQVI3BC40glhNx7
usgjl71CnQu1X/nV1X14H+tA8tJZUAAA6uwqRj1bWF1pio97UHrKvhfF6a/sb7/OQ5Tzdg0P76MB
Ol1Bgz/Pw/MLFGmSF2TSIXMv/y8GhYyxksw061AaBdpfWA2EuRJs5DN/AQjlpipMPnlp7NJxVAou
oDYFQMZMbVNnglFAHkuOI0wxp+Y0nedauu0FAyFzjXz+VcG0m8eefDH3hdj9mJ0Cgygcmvgusf0K
lccCQHPd3YqqoL2Ni3zbxpucYTNz0Trkic30TV+QirXwnw6snCy8FquLKjgUimerKosB9x+JcWJj
CY83I2hqokeMMRaF5xPCbdcD8SQpdvv1uud0+9zgvD+aeosxsCXxGEgbGEKtEqKQ8co/lQZqKMpt
itXuL9WfhSYfLTyruOtn/7GZ6dpQLROXzihWD59ib8Jj9xB2lKC7sdsi0SrR2tpTu++5nfqaR/7h
Pe8KxrGOdxdQC77gkWs+dC1OdanwIc6ns/yXzJmqAhMveeBoyNmtl/OHf+JR2Lk6OjMYYkt5gLRN
slEcVMQKleXtcuoOI4PG6q/nD0VGSHqpCLEyDyMaifc8RFswMrxcmhGoV1nBDHv8riH8haDNRmNK
d2DEQyY9CZvtR9vTgBndE9y6eHb+aT3ZoKX+0JPe0rZfIKeYwCdqmvFGZkjgX6LZry2p/JmCQ7hA
M2MoVut/4mX6lAHdDDdW/JAXbC8j+aNlNUFJmT7jX2XhF3BO8CbkP9l/PjAwL0C+70ryCqkD3ViB
OL/LL9foRmk5Rm0NNQirxYHCcGJ/p6Hg0lX3AWu7J/XGKdD8vOKT/kvJCeNA+WeXat2xy7jRx3fP
CIxL9iByYfB7xNexH9KZmYXjqIbHtW0EHBmeNtZQDb24I2uzTtv7zkdFFckag3SNlu09qc1kYvxE
ZRErOkcWJVzgeUhxqnT13uTsYIbaRykoBIQDnC7zd1cb0UbcCDy2RbmXIbnJrFmSe8gsN/rgTspX
HQe6mNLjeei1LTIzrtkl+lmA39mKb5xl21dIgu0X7Ql0vq0Z+0sMaMVyhDu+ZBcPJgaxLgsr3qK9
2Ukw/7tX0D5s0mz2P3F6u/zZHbq4XaFnsvJuAJvGJ8qBGHF2Vr67VSmVBOEfbDNrOibHI8sya92Y
yaOlm4qRRkdIttJ4g4hRLuh/av8cmSudo9PBFMiANfsWVfPGOHhxJ0srYP0FlaVX6jp/g3jE/41S
FdE6S0HY3TUh45nhtEffD/PaktywJg1VPdsHLV7ctVtMZNbhdDyz/h/GcVCvOqC61j63wOLhe/fW
x2rXyz5hupi4VlXNMm2r24ZEfOZQ86vQLJlDD5cvPJQpZD61iPdzKT1paVFUf9GSqFhdQXVTuyf3
NS8FPpeOrTT3V8kaLH/iysAWfrTc6Cy6MDKQ/Wyg+5mSpdu6q3KNIElL5h7xz4wCzlfECcWak6K6
YGS498LkIp61qJm5vlvT8z9XWT796ZAz1CcbV+I+XxwkwVYKlaOY2LY1/OmgwfmrSsbt3BRA03B6
2cyJDeKF1+UH9nV60qKnwp/EDVfkZiRb9wiLOsw9RLYuSgyzsPejXO6wIxnX685tvj6zlRfUmcfI
a2pnMlevXAcuvnkzBBPpglGAt8+8SnlOGEaYtMzKYfUVhAAtiaRKbw6K6fEOJhne7/7Wk8L6JIs6
dNgWfuTn8vHFx18p3fSHOImuKuSCR8Z1ZqwIkO3OVwI30hSzFX4xp/zz54pouAWPcYdxUDYGYBh2
dRosZPk1RH/JAJnFn/PDavX67w3Li1aMu0ms2dWCwLbmIVgfcuIVYPSdnn7UmJVhTdAeCnI2NyXD
eYCimRXGBEXy0MeCHAP5+dCDZLkDWIlKtA79HfU/HwgwtWz4F/2fR+A+mXZ1upZp08fzNGeL2eVQ
/hC492bKrriZUMJJ1dS9uDgPtrBiYIZdGUCU1FqRswg9YDvtQrNE0NcF8ie8MFO/J2j59CiNDKTL
Lr5OmQSimOfon7vLQRlTiQ6Nv8p8SPRO4pFkkvmj1qYVNmTlkw2YK0X7khvIvfZmDOn1IccvTc7P
eH3yVoFNP6whyJrM++jaOT4QNYNy46LOQZ/vzy/9A+c++orKlMoVgAWxlCnF2D0Fj8r+ltwcSMSr
EhAOEHsTL69WgPvSDBb8UPqLUr+nO9mhekFpbzjTdWTIJc/4KcIhQMHfVn1IJV3Kk2yJEViE62o9
aUmDLclNl3sVwrceDkKusVkm8SaM/bE+o8d3pRIMAnecioPfxJoWpc+X2YQtvXnu26NfyHt9bd8f
+QTO8kugBnzcT4R0jMsdijitqzoswVfn61u60ZvqEBENyVt1EBWTDlsySNaN7CBpXdE+om3kFm64
sd6oMX2R0jV5gsBNHbH8dNpKaVQIXLhvbvM6yrarAGKT9OLoIHHKezDkp6XH8JbjtBRejb311rWS
Wn5FVNvOmNnRZZ1WZlsWtuiviiIyBS7RyLe2Tkfjba+vry2jmWgfF5rLNiFUBP/AKbHp7w7B+n5M
14bYv2zdaACc/87KZcCTmqXh3Tx6sNKtHy9dBIv7zS59yTi5yX5TLDz4XwQdQvCC6bswTPNkoiOk
2n9YxKjAE6ecinP6ZtJNAbNIyh6cZDiZA1xF93U2w7TspbeL21EkhTzi0noeB9ic42P2vuX4wcRV
QqR8PxnuAaXEVo5ZMGi732MzdfU0GtTj0qSo5loc7iJu22Gq3bVVwZOKvG+PK7BLfYSbBSUL1VFo
qt4nXrgOZ+zx22S8/xqYSThrrE2TRCpn0R02KfJgNL5UzxWMWnQIRSRysfEJkMlkwBp1ph46R1Bt
mEhpKagF9wMpe84z4xmfarwdDlOnNPVOdGFjei43WdtrMH9EWQA5qHAW6HmebE2VG25JtzQ+eGkk
FayhwFWLw/b45AZJgpAKfTzN6G1MoHnhHz5k8LzLROmgiJOmNzgIh/1svAX5UhlpRndpiN+8+Zh7
nDwtCaeFCDQQfYTF/o+KAF5sLdC3eCPLfGbw9QrOoXN7VLuslpmCZsbUBLGMwh2SufHk6RwmhchK
1mU5LB7iJXLejOkM/ajpucjtZeoNvHUHxST6mk+GjjLPHiZzHXP0NZglUKPAkCweZHEkGqYFx2J8
EYl5t5WCBXLGNnf4Grr561aVOkKW3B+gVeKwhpEJjybv8THB44EpUyVTW5h+IqXw5N4/G/j7s41H
ejrteCrNIWxCtxLyz+IJnPzwdgclR0NZdhfRXTRL5pfwmQ64G2KqXOA/qDohjiPpQS4PPlm5wCSD
QhwHJUut3amoYAhuqRB3UeynQrLFFnvtgzlYWniBBqXZnT74e+vj6d7toPhAqhf374CO/sMm5w4N
egNNs96ZuR3Ct0afeOBJdJzY8/D+Dab14ma1H7NGp6nq4wYt/hy58O4nlKLukrWQM4MLLBDYRcv0
r+Nyl67eG458ygLmUryVl2zsN80AMxvkprco835quBXdz27nP0/ae9lcQGLwH4TM8MSNy4dJTrpK
kEqofxMdyegVrjtTltlfnK8cppkhQSEERhxQfpP1oUSPpk2JsbexcyHb/OHEnABMh1WrcrvZi7b5
MhUQ6otWvP6NttzP5CMvYhcs4zzAa815ErRPh3B6LbG/VT1oghWTx5wvGFosXoyGbAJ3jwJ/5lmK
d3UL8im7c4pz+k7Ke6cOaTTNbaNMujrLUoU+67jIwIn5HW6BybpmsqlgV4w9ZDbWAfEeYE10WKLJ
4kByYxu7heEfR6I8nhAlHbgdPiOB7lU0oeaI8yIUpc0ar+DrntDBP8aR0qjM9cH7SqA0amsd7Isx
xGS85c1dDdVrQ3p75qFYUz0MONLMp02eFFAE2fa5sNycEnlrTFP4HmxXwJLA9/NaoOGPsI6cX7KN
7PXG7gM/BPvo5vu48Ap/QhEe4kaUpnIFdBffIoVksSYX0CxqLy6FFleiaJtHhXSmtJaAw88U0OI3
qUrHEvKmNLw09mBIFsWJEfm7dv/CVHogjUo71986Y8NjaZpyEFKObKx+lDKJ31+Uwp0L5Y55fTSJ
u6xIlv6hdOXWRAfHNHypE5XbVOvqTxvDBKx34Ibyj1dJsDRMLctgn5AmHKIsx7qIkkT1WTcsZL4I
PGuXnsiAQ2ef6Kg0RTj5r5ImGpTU3gcJg0SR+KtuQUl+MnWTaX19/aNgbYLrzD7O+i24XCYNawuK
RulN01xjFCLWYXjQi6BUT70cJ3dEkrXFshh0gm2hw5NR4qMGAJxvPtikBhNViYd/E9YklNA3plD1
2Jb7+qDsYfrCAob6/YGqeXh1Pfx2mDjFIozPKY2XEAic1CbsTGJGA/ew4NLFzIwD/i2gHmpPjblr
GACVEYhU322tQEYbDmhhgMtbu3+0p0FeNM6+q0WNZVG2oGMfKghP3wU7hCuxRdKZn1B/V/qRt1xq
eLTjM6DvXpxSxxFZlrfQT8vQzLa9KgSy2zQ9ZSUDQvuD1/qcaUPea7g3xMac+DXy1kCPUrtgF/l5
Wz/VRt3/rmm8UALT0oTCqLQ1ye+b7mIRkNUKAL81bXHQ2SmOyNzYfcgcaHXnAptkuLchKiSwuxfj
WLgb7bCFXieKVGGQ7ZKuN+sJ2Mu6UJ2tdz70HhQw4zvdiXQdHJSUPcOzl6crYMG4MVzccj8F4OOi
ZuLFVeTCnWAsiCLa9vrqwm0K0Y7Dd+Dnwg01tHq7AOHlikiCMH3T0jVxL9vTmdn4Tm58oBC1pkrA
tfLUJohWzmpgPrhasEC4kPTqdf+ZdfbcxnXbEyr3PIq0w5mH9JM1wnzS7fUOjZez3BtQf4DLoqXZ
DgT/ftjIVHc/0tM/XWPYiiTd5An0iUAImww3Lov3+/BdV3A+cFrpATCKjw/QPlIR5FTKzJAmAglO
zjJ0p7uQ4l43O2tb99bELxZVtPIFhPKxHnvaoFQdPpLEQ3dxnuJvU9qYrsAVtJ2YUC7yinxgXTKd
qIqCmHdv8iYMqboe/iQjUESTjj2mfjLqqzjXL3rSSqCoF8fpueABZatog2bHnaQX4PPuv6DWLhyD
cjcGZVn/ffo3ndBXA88exBr4YMl6xfl0KQczkn2+TZSmo7RMv/AFiPW8cNRbDztCYCfz6GSGFWCL
Mre7E3emFW4FJsygzE/Pti0kdSr2gBfl1BdRw+8Ybzs4kth41KeHZXT6FR78NJuJAF/geZkV2udH
JImvJPKgmBcOaIRFngYroQAf9TEV9IaRBggTRPUk6Kf9BDJ6cQusehie+ivo/bZ5YL8/ZD29OhtX
UQSOBKleAOswi60yLAilQS7Vi1DRRoutl7ZzeY8/nNMb4lH7YvNGUaHBaBgLyIh7hmTSJS3xhL9b
uOznGyrYtg7xzlPbHY84uBwlJrsSzDYWGKF8bvkMBCnb/L3A/+KIUo5fSxLYQpnzJ9P43O/filN/
RmcQBediNshh/k/9o0ltCdZctv1zJxpgUi+3CTFh9V4j4NTLqO40AFSEI5de0YICgtAdPKwRHlcP
A58QHPle1iik22RgMKR9FTA1QjPWcsBf6lDtdCrqsWvr09g6DBGyOVmAeRvBracu+ZGbjoCceA18
YMBLGG6vfVX6YrRVgm73fxCic20zJVjIuAVV/qJlfT7SZGbo4EpA3Bse6Ezs5BWgbxq6+IXGixlk
cCLWpMKzaQdlUZAHCskQnnDKTQec3PVlRXcxi15N4lXMuofMatruRHpd+JnzWk75vjkdj9U8d/mq
/Fc3ulB9zMVcIr0Y8a6PWspER++yKTA0NbXlBDf/GM0byl8EUHGfkU6egjGRrb7VcVYXh/lx/QSM
TzSPWok1NSRDvKHEaEj0Z8zYMYBMjyM0jHNvYoZl3jqFh3PZ6DxidpHUUSQ82TGnlHRjVtOBpHMx
gjf2w6cZuBtMQ4Ssyi4TU4N9kawP903FHXmJdanZSc8oys+Mg0NvoYHPU+7T4dhFhaeO/glK7vZ+
cBmzV9vrxxDM2f1/V+mzQkZytrfgAHmMwjL9G3p708dPtZkZ3ifxBVkQHYVHzQ9THXewYFPXrfhr
ytv9onImm8fvqLN5uhZzYDHfrJ40W/vXN0waGRDbLQ8lB2gC4kNKibF0RFzcPhEh5ZoF624W/w4D
GFDdtrIf2i4MfIcpt8cLK8aTH5iARO7po/ld/g57BnHNzSJ38FVuapm5lFhYBKhvRiJQxAb2Of2c
Z/sX3QMZiGy2bN4FCDXbfyVajzUT8327U+Q9RbNa3+9gOkjZc2Rh72dlcUXEblWjeTQAmwikEd31
izJEfYp/BJCGr6fjx24cPAvu2jU7zgbKTk6bUNkoLglaFI63tP2oyySkwyxUxn6CMNynOjBe3wxh
PzfFQOiec//4WVZRn/BZgqXBDMAqJGcYDIH1TUd7f1hLQMszGYsrFctKB9yIxvRZh4QuL4kBj2wr
mAuj/hcUs7Zdtndn9JPxUqs/yaSHcDUjI1Ag7FbzC7OuCqBLa9YNkHd1C3VUQsF+FycY+iAQN822
KOxoSKaAf49pPSNflNRagxu4aai7SJhgFb2+wiLu7L0xOfM2FFXn8UWB4giQxVy4mbeo6KsZZDE1
1dJAjWUpJhK2RqdpHA22XHZvE8YtKs/PB/7ro92Nqudf1LU7NjHuUDNwGGn7bUO5C2ooLq6aNnEB
a+RdiAi6avhiQDP8NQx9E5pEisDqZJ5r/PGJ4OdUoOD0pJveKqIVZtyZz2zIPqcOI0xLgAkT8iiq
eqLP8WnT90BPvVG0XMfa5YrIonL5hxu2yYApGbkwEYSlL2KsEoRvXYDJTjT3UZrBHqBHx6zTvaF4
RkGPhqQbJj4ZRNtIvFjzM7hp4kZsvciuFsv/Ny8XBTbV8LpEqJIHtNfCQtcqdCVV54u+vUYkCyuz
yM+RGG5xbBR44Ey+guERvAPsY0p3MXVHBJ4nT6GmBwweuKlP70LRyEpfvvQlrsdxL3MunEieFf/R
HiMOen81jd5Oymf5/BD+85c0VvflmpfZg9wMKdzJIxIE1N9T+95Q2z/QkRTxojTEvXpxezkiShMA
GvDIyw0NwJEc/eXxivDpgv+wgCpFhlc4FSPVRJO7YDQXCkOT61een7JEKN6mq3zobbrCmDXxqv7D
rZYoYwDE6cAXYo5Kf5X3b2dDVM16aPGqmeTTwWfPHv9/XvT0cHtN9YFjeHLYQGfalLhMxatmkr3I
QxdhYefXwGvloNeF7b75MPjnw5AN6gdEnyOr0ALKl3AjNxm+6R3dt6L9mX8EhgWe3dQb054QY7kn
5NdHbaEhbpEBpr/4uZdDPXOQg2xHeF1oH9EhTkjyq/t8vTN4khohB52ghIw15Gx10MpXELUXfJE/
WxBJukNTD4tArxZ3c0JfmndlIL7SXOhpybOEnk6dsimIroHpSugXCnIPMCRKKZrr/r9BZHN9Fq3v
AGk08iLjxK2JMuVPMW0Aua0pEpMrpObj5vXTR7U8ZbRX29SkGlfQb5ecjRRYAYhveNVHiNUT4RyZ
MBxoEsULYQaWkrIXkfyvgxfk4DWQzArd1CYGgLBpMRa9DryfDQPA0cEMmTDT8FHMEh5Stp4cz7yj
Dm1fEtlueftwAdnA5azxsgZZtzicGhYzp0pxkvjGAD+xvsqNrWefQmf9f9RZmFfXS/Dd9jvavtHo
8UWGuzXzG3adRVOENXfRivimAqxM4Q8Vs2fkihUd8AWSftPcA4JX3up4TxYAVCAjt1EIkCS+qRUt
BZ/3ebyR1uA2njYrcHJHDEwPh900Bxxm0upeWA95gRxf9odwWsBO4NdOO/KJm5meF96fx6MKohzs
45KKZFz2IzIrNMw85Qvl2PdKVFmLcBqmYkPA8yoaPlU/0K7v8/cjKbJuSf7KABowphmCkkn8Qsoj
HSz9CxqYLXDFd9YaXsK/zXmTAha+NgLna/J2h84vuouOTYzrD1XnnHhp7I2mqsjNVvmPRcxTvxMe
cCAvWq20KDki5oS/GuCkyA4kTzMbjm5Is866gzQpU8YBscjQl7j3+0onKJjU56vi2X4gf/HQDe4k
sS4KuocBCLdPzVRn4Xuo34YhZn09fq2YbGYPPeCN922c9PQZFxCQcraU4ba85KnSNpmY4Sc5ge8i
pUX0hq0fDlb4WsDagnJW3sQQVLAgWRqFies9d19ewkRDxZ4UpAR+RiCtjXvkkWrBNHNuYjxemDMW
D0hUt9kVLPKlirNU2id+SazGbm1Y4I+jcQsAcp71d/4olkanqF+OcjylGjck3ByJJQ8cdGQyppTD
WadwhzTdX3ubtC2BmZWvBFlJHpuQ9VohVTNmUuSSlGFcYkLLhDgiThinCxLS1WU4dhlx0vqRh25d
pZoPod1XgUQhOt2uupw6B8aWp/1EyBdj65cmOuHovluve5oiY9dOmgncl/ll8F4ourzV/3L8gCBD
h7sW8162jXe6wTwyvDs/MUDpZ7a7yCMEj1wtR/Iw3LEo1vCtKi4ntaMkr4l1jEfbkTMv4u6tyCz3
Qx0zdag7jsUo2XeigSp59y9XJ5D8NwUFm+BzPocLh8+SjaKglMinLNK2qY6+AbL6XYKN6tCot0wu
mXNPAqRK+Bn0TJ0krCjNnu4luk3g+NCms0Cqs861aqH7LQ0cBVr/2fL7iVOYPXIRhO+9GDCU1bNF
Dxn3dM9QN1Wx0S31q4+1YYwqErTq96/j81y2gHFPz0mdsM03RGXmGz9J4+g7D+ZoF+28xWV51bzd
ltaoCdYtfjrF/VaTNqd7QdgegdRc32mO1Ob96wukJ0Tyi5FGugb2UN8zR/aU1mg9FDxlb86l7YkD
eBft9Be877FkrnhKAv8zHG+y21w9zXdVngt1vTQrpFGudHl1BIE1W/RRCSOFhkjTsfXX06uOTJMP
imtErzemcDauXldarwG2p7iYS1VL2/TDxWF6FqFWqJ+xRtyUTxiFiQzaDLt3sn4uIy8oUqT9qd2N
Nbvmd0Rd/xvBjCE9XItBiSSpjWUJc4h9UZjVdnOTE8VjxdWIpOfVd6InHywxDGvAVn60yf0GQi/a
C9sZla4G4ZqnDRwd/uBqGND2KdYkWtCAyjD7/7hqVWNVeywYMHDIdhDvmjc9IqLuSkkVF2p029E7
1stKFgxkVsZsgqFZsRCZytrqV/q2KJ21lGM0MTMT4NLzLWb+TyKAR5v6DE7AHCiXA5I7xTDaQ1ug
E4PZ24GI1hB5X/QSb32FG9bqWqUXqP6Fo3W/tCqOMzy39gEZ8MtogZXWnLjg6CI+tPb7seAEdPs5
N1NFLTptXcrAlYb8p65PTS5ThwOovAr8I780Liecl4JKGIC4YOLIYg5T/rloNY11v4j/P9e7CBpq
Fe305PIaXcfrefuDob2Hqr0UjfUzMzHB5ec+WhX3myWeSRd7KaTIpBWezliqh68Cph9eyU/bOfwn
ml3PUvIbsGlzXQy1ewPsa3yoc+qcX6PRToDEWVySmlofpyA8GNOQhp2nh1EiItOdUn6d1GrEhv/C
uRV/HxPz3p6CIWaArUjbcyNR7i7qnqJEf6Z1tjrCwQob0bmulJNPJEcDI7XVCQf++lyZCk/Wq91x
l6S5lIYUOwyrXXl8tISp97UXPqk2qhfu62b8ZBCdIlGk4Euw4rH/dHCT7DDR82a75GbDpQK9VRlh
GCzx4ewbsrAy+MOZu3kYDv9d7N9BAFL07MIql8uTeMc1Uh57zYdAcRIfKEefEhdJQ/3WUfQL8gKE
Gx8kCVMvAVm8054p9GIF/HZkIoencxIVMC/Tprwj8ouhKNA5g9WFUYaeULiK79nex+29RoPfGab3
fuElN0DUedsImeO4Pp+hBT6KXnhlerCIP+L3jd3PX9/xrxe1G98fgMB8uusjSs3yVK2JMgvTHYWI
GztoUEeiOpY9HDGQn4bnwrEKu51uRzZ6usu3w5bn+pABQ41E1l8ozS1/8wDKKofETyKR8Ts6k0wu
ekXsYR5+w3e9T52birTrMO20nGV/yw4nAn2YY7uFi2AAuom42Hu4OCutV36czqHwd1egs5b4djuM
03KksqDJx1dgQSRJt6Hpmdl+KpdlG/ak0/YFcmidn7FqwKO/O5k0zR1X9czn4eCL6wgbmgFb5jTv
a/57VLtINu7c9RvkZVC+C6tgCg/nABqylop+O8HEiAR7UN7xsQ+tkeBIdyg4gMgzO7FhW63x1z8C
TnTEvrfB05WiylncnGTyPFlbMbRvFKgPJFcQKo72xn62ggqcdKLYb4fM6hinaCYVyNMaMfjtF/vK
Bpc1rgalOVeMbMHIpVxzIk1ZCx6lT7udyJxQj7H19jy5T8ogVGOvlnPlvdfZXJWLKBDo0wpxPI5c
e/jmcH1OPBcNneYoZILmG/iutLLkrbfdcEwb1h8lZkyi+9Tc8JxNsK0yitKBc80POux3lx8bAYtm
ZMV5jc1Bed7fk+xE0bVKGz7ds3SsPBmiQ1JmZv+JJSlHymPe3IPvCp5fnnZey3YPrIur29GOcfAK
AFJSIUmk6R1NZhy2B8sgnkREXyzpG0u7dTH3ZhZh8ZcW9pB+4JHY+p71N8VXtHtlTY4DfHNbmOJF
YvcCqWjFM5MXn70QQzjqmRxdzBPpIkK2EF27McLPijmL2SFvuXRAehlurxDxrU8oKTqjhtScrw7O
rSHhGnnWrv6LbsHSZijA49ax++XwEQIMU6fAsUfIUoZGAbGgnOVW0hFHyOzT5WPOpoC7OhKX3ykM
Ke7ObXvTZwg9FY4VAh5JrKQL7K2hcUcewuVvKCwbhm4fIGEYiwoquDDq0ComrKP8FbPxFHCX1PjM
KnzHX4wlRhCvfHnjSxTRoihPbSuvFUJI61A28uvNM4w871abtQANC4JlxM22I1YUoT9xgCJvOnNj
eGS36e/8Oaatn1pMyjFFCmkXA82jG4g/A1dW5lkEVdoJEh7Wy5vYngXgAJq2j1dcdDVcc+EGA0ct
iCuTzeXHZDshSAhQkX3o3S3De/Jou3phRpf4+PIVyK6vwoje+8l1K+LXOTizH0t4BNCeaMG8KWGO
g32xdBnBkPa8VLPG8AXoWqfjqXlQ1O8xRJR/fEFO4bxpDfrlC3QRYw6vd8KBADvpyDcDjBisG8y7
eAif6ozfEWp8c73gYpTYLjPUoY3VoJ9hLVgB7B33QdLOExMEwhigZ68LwoML6dHuHQ4Def2n0o6r
jiIQulXhjhzI5nn/7rBY7WXaCRiXchQr4yx6gJ2PrsCM6Ghj8Z1sgmJeDw/ZTEaqdSQ6fvruaIpH
hu4+ueHiw26ysdc3HVyiEqkazzmKgKRWxg84T1jB+eRL2JGBC+waXnf7BwgtPSpfWyLqFSIBAi3/
LQDa8cBic2WmuYoCZsicZ0vk49X9cA5TrIpBOT1LV8BYX9nnHA5uLrZjFjWo6O0bwi2oEEXsxvPl
o7NNZcdrpDQjY1XJ67NtLg/EH4Q538QKgGc2Unx+XJzW+WPshEAvCsS+FyJ7c3Nluo+I6F2Goank
pOOtONh9JvE7a2TDmlLkAx8EZiMnArP5SPmACcAp2DutM6qxQfYsQwtNP8+L7HiGt8qP0TcvwuVm
b4U/D8Y2yzVnZyDX3YaAmpyCb+NtKtMZJPOk+Ee9UKacbVH7+dfmz/4qIrIdhIGcaHFcD2p1PNWV
OB7TOjVKMsH0Y8fAnAxrSzLF7DTW6yAhHZKlAnn9Qt2nSwyy0qYiztPHQsUivLVSSIjkB4CdkaF6
f3yOyZcTXK8zSXleG3vA68ca726cQTuh/5xxcXGipjutVngoLh6dgwqWr6bPJVVd8xBVHYnWvJ1r
IiFwH3ZPaKM6Wdn/FInLPZKiMdVbWWJZBLumXUIfazLCA+nTGVDQMZv9Wu+WQxxxXbPEAi0Ne5yp
fOP0h816DN3LyfVm7aZosEyuh6Y5udQCCmlE8ECN9yWdziM4/4Y6SZoId4ZBheXFWw+deXUcJLkw
FZ2Nv0Poc0MEqC6woXZ8zlxwVJF8o8JJIA9q+6NJpLhkGnBht7ptQzTBUz8zH2Brub3/hFj5ToGX
HeY1VjxMXo1VGIQvcNlzUgZT83B3os2gMMN/x+/+3Aq4S22l0YwUM1uYqCRS3cSAHEda2J9XozzO
9BAdWXdzUcP3pTQYAO7WHjUTGbPrGFE3YurYzZ8lA31AQPsA/xY7WUf8tdDFUTGd1D4VMCyoV974
31SbQ08siBBu9OlfPTZoc4U8vwd2dluMgoToEOJMt2/0LVKuLpdTFYyzmN9GtvB70bx8aYDLVufe
rJXlh3JFm3VrQHY5eEaFyegohKFAfLFCE8lE2ixvCOEIi/okkIHCTCOPLXmnFCPHUj032QlgANUH
DsWcL0M3I43I2iY8ar7D24G0EQGTCjUVlQ5EhVr7W30v2FdMhgTnGBaQ/BTf4TGRvhURL5min9Ao
kaRdJ7Ogu6YFAazlU6kCDNPJ5p2mRvgR8VbleZ+Toe8cpg5xPowDPQh5/na1nQs+0QeFjR2whPBE
rcpGo60Xpmj5w2Cc4gcWZX3yhfXHnfpDrGfPSnjiu1kWEuLSQJa+TyRXjyB0KKZGv+E8E/pW/qgn
CMVlQUwaUaSIR93sv+FHg1YnJ9XwfT3ymDYefL2R0mL+Me+aZ83Em+rjaTxEtxWkR8Qw4/Nh6sKE
53XMRJefQpqBp+7ipnm1roRCUAK8gAXvdywvKXpKwJWVfs7mUMsbZFeFncElcfN1uNS14xhFw9X1
4gAMWZoV0QHeeKaIS5hJU8GR0Lepy+ydikzJuHTjVMlCS6BLX5U5cODepS2zY6sgSv7U9qRXHWRl
XBjXNU7QFsIsINhUVp3+1+SHt7H0ziU4nZ6gm5hfGYTkLbVzq/PHXsF0tkllyZ7xggiGnbqu6/AR
6ppRa5YbKKouswcqeOJbbcIhUmpcbXLCIryZ/GXPkOMvVU9DIY6EOn/y8BgeIJH+i5cZgtzJAliV
B1jO7piVfYfepEMbWM1ezn6PYWWKQnaX0ThRETCGHvwdHdhdj8lHbdQ1CmfjiqS1/0hwZdWJFDQL
IJJd43f6+vh3sxM31r8JtVjHHQnrhK8KJlu+tM72gW2WfZ4+M0fSBwgq2EVR8rNrKBwee594Dhj6
U2XEjFAM4JvhGo96f0JLVvdIGBo3wggdXxcyNwcedLhbfqnSXdRWHHfTyV9MxbogfKj9sX0xGgz0
u6ShlREJpLoSyBOYbuSwBIbJE9fBqXnxcxNfm/LyqYjzwp/pP0sNrAkOzQXF+B9UYSLPacpxbvoP
8IvTJpfG9VOrfF4XfHJGS1AN5c80sWuZa3LeoLAMb4cNjLFpQxnX4PwHOxzBBI4D6e2E9od/0Vtr
GhvknzTXvvSY9pz7m9CBiMONQyxEu9f+S/lyPUEb8jzSDHLv8XZPOhBkg+pNmObhD/olgqcEr0TL
p7oQ7YVSF+4xGzt4TYhO4/K+QPPQVOe6Psi9qZByYbUMDJdMnhimYu5pXlcCXMEDply09sQq8y11
1vkXUYS6kJ+B8JUEVfuK3nhbGAzLISg/Zo+xPf9GIUE2QFWn/dLj/PsNQW1Tvq/72EDMw690rDzR
YB4nVspmkMuPLWBbs+A6sXwHtAMq/NhUMPhgXLpEO7jLRMcIfPE9qnXVbyNdpdWNKToLWSJWebOq
ARFbnYASJqm4zSOuYdfRRK1XSLWADvmMcBhDYWoM50RrBm5+bbkQh5uD3iA6WIyBkJ495HQrTGLz
ngCy1IGPB4oiWTlr3HbPo7J/GC3oSnMAhLHX2D88dPi8i8xtfrhXPV8i+l/li0PlgtPazQBYLfIJ
wLAthiIyfEH6sM9rgNE+juBn09lIcaT7Xew5CACb3DOwG7ZKVXI6VK2tIjpH0CUR+AeRrDCo/3nP
z6EEwQoCAuGBLsHG1RExsYFrLTEmjGlvDPnIWeVQy9dERxaaJ5PtUAU0pwxLpyvFmO5f0e9m7k1O
Exf311mGGbxENvJ259iszEwbpeIjuvENt0M6g9AieM6orfaMjUD3YY7d1QKgW31xsWkympk4R4mW
r3tYRHkfayCXyk7sfB9WYSzv9hQ08JyrFFsZ9XVYMhYGxzsxg9w0mcVodSoHKTn2vAq4KJTGfYu/
erMA4qX3nMejQPF6Fqgpv3cPArDeCY/ricsj+oAn3XDGmjeaCXgUoMqWY60w2lYuvmR2Z42aqDxW
sAXqGrrgjgrKONU3xnhe4+UogTXVq3sNIU9v6tWli25SjOvQEr2V2/5qVWISMA1M/1+JN5yiYgIC
mzPstSrL2J33+5ZITjIJ5T+3PgRtWwWAkj/g6YP+m0zCEWC0ufz9LuTuSAxg3tv92pMvTRUu099h
L3xwZyOI3Vjff17eliohvqzeX9c8Ruc3y/z5QPBN3UdTMH6AMSseI0CMqn9TNzu0ZlaLja4OM/nt
8w8vaneuhrhktY0zMBL+ArUwF/Qa+wukr7+UjX9EW2Qj/Zj+9iQnS3D8f0QTI0m0gxYBU1mqj0+a
bOVz/+7pg1Emi8HOWdQRyNheAJa63WoMzAGQhs9KaMCtKDojuFRW4PPbDAWcBkeqSR/YqFEhbr6h
8aPTmdUkHmr0DE0SLtpgtM3fbNj12WSCYmYtjrIkE8EdHd3/ZUGYweWOTawWaAyZvdlAU7l4YOLH
wov0bIcaW5++5K37RxqquICeqTZ1dElTKV/hbXsiFzcHgMpAesXPE57xDE5TxSF+rOm8ophon5HB
DfqI7aKTbHVf2LUBUO8bliihxII72Q29DfLgXNOBe0MpO4O3gMJbIxvqPX10MpYTJa8cgYdchEE8
1jfFVrovvD7cFxFQ8PzsVAs/bQuVtJc26GXFW1oX/th3Jct5YPUhrX5/1hRRkX9TI5/uxS6IU0U0
VNI2aPPqKkVQ8IcJtU6qBytg+CmWbbK3+DgqvHVTkDcuuBsXUvx7MKCpjg04MzpLDU27yu6qlrhY
0PHWwrqquqZSNI6j2yW42DWku1lalx8qSTLPjjyzmvWe9zu11NbhKFF5WsqzJnJBANg6zx7E98gD
nzYAd006tmcIKVp6C8aLK1uec2R/gwStubNSzD3QQi7asxFEzn9EQ8CxixARBG0K7opdz7JxwgYc
JOwUZAmP/hYm4jUG0oeERub0Gd76+OJilBopIqPyO7J4sxO66q/K7TqCL/UyVWOaAFE+qPayn2b6
pneCRFXJ5jt5VVeHw+Qkt05zxLUTS1mJqgMuX9PutiTjRIxqksEwn58X/71Xg2XSqQ/JUBzBUkMb
ohXqa1DVW2v5v2yYVfm/33/4d3g+YfpIEAISqmnHv5KVW80gIQODIU1b4dhIRWPB9u2TQ/NHZmRi
fsgq3rUnvFoFdsmCQnNLxKpyjeazSMDsDUO9aokgSp53VJZZ6OgGn56ackukwoC9+y1gwq83I+Su
aNYM4PHECazpu4etwX5IDTZJBj53JwEvTzIqLqvHduptVPgMniztMa/oa+/CxXL6dYpKZfy9sWlX
u4srvVNqjQkcim+CW2Rr8z1pkw7L3ynPNRWe/9akgC4MgP6vO57J8oB57fhvpgA9Ohmj6SDLE72H
PLIH/RPUmAVPws7oBwkdNgGxgm7LFXuRVPr1NJwQHH1hrloPc3NX399FSrGFeYjBlXB0yPW9TWVq
CYf2eC1Qszlb4kOp+alP24UFhcTSMW01YdJGR5KGDz/I85GO8HomkAEZccFIcRuefzpcPMsFB7UR
rypZPNUi4KmB9BOI+RXzkJziWQHvIS6BiqMMdC64jMoaa4Ka18Rz07D7dBS7f1xRAtSK1xIu4J84
Hf/48LbiKicV+29QB+4ycCqvn87aLYkqnMlShiuYau2d0IWdqdwyv2ZSOg2t8pKlkdhtf2kMq2KX
Jd//iUKJC/H5P8L6RwwJ7BWbOb7vshgk8ZtDD88A4DLiDVAvK6iU4+AQ75p44wiCkCJ8eXB3/iOp
JkUYm9nwa3OH4s+qQNe1Dv9HMz4R+qVjOWkCKQlSN9rGIMK7FIY2lyaGx/hHO6FZdbyP4Uj834KG
0WqAfpfHXxTKS2ofWuw7uUZa6FIySg6K4yzl/gqOPYHuu/lAp/QgkMuVSW8TKoXd+CqmbZOj70YT
rJMlEOEvFj+18peKgxUufclktE02NRTfA+qGpi2DI5RwVyfCQdRTPgFCxcJyeAbfnWZtIbQ3f7F5
Bg3xcJc9bG+I8dAk9hOrAxCkIvahCU3CMWC6t6Qz50LTz7GoXYuQ62Ev53db8Lv12/zBus9xCgSd
/v9YyooFo9CpEqp0cO/5os8XYvEAlNwQjuHeSzGPdG1ztiG9RLqGhaaa2JD1PS+HlIccyW6RDCkk
TQ7R/tVJAt6nL0UhRyjajsVa5rrH9pnnnWTqLnwZQcjwrMlsXxngaSoeJ22K7iTpu/zNKkhrYvZb
FWeEYRdcxtiO1RmquxqmSMbxqOvuVVlT1T9x8RLgNVi3xkuDdP7azyUhWs32pJZfXxGQqdQn8+nw
5+iE0r0g4xnk86uHc1j9M3LmSn+Q+kagnxfpO4vAw6apQ4IBx33MvYoZPWykJxiuTma68VO2wE/e
W2PpxAJKMIvJ9DjO5qVwEcIjvM/uFlAA/1+tLitVwVBcj99bmKOFcjG9YycGqoSQ2XUGkdtFStzW
9Aj962b+h/5yGePXNWFDCUlyabKUqANtg2Z4g6NCrzGg+E1U8UXSVkf2XhtRGDsFv0mVT9pBIfK3
W5Rqo6Q4Q/o2hgYDoYPQgEGL6KUbfAotXzeq40g5WxANsfwsf0aUNAwZMMfGnZ6FOzF/W1yqRYVb
e3yQwYH4Oc5Zeke4T/KUY1iKHM1nNpIKPfJfxNlvN3EDMNEwhGYPFBLvtf5dM2j3tCtzSqs1pDsc
Pjnx+cjIfd2eyghNDFsb/NEl60h4HtBtB6OfY9Gr6bcUK4gVF6Y10yHPeKTYxeVk/VMB08PU4Fju
mkIwh2/xwXenuGrh3m77UFpPxldIHUxYg2r0zXN23inyi+AKHlVTy/N5V3vFq2vtZWy42ygdOfOj
ZiKhdFISGtJZHENB/iCg01eJchkWzz2cVHljmb6rxLA0iRCl6+lOb7r1C8onefr8E+Yq5fo7MbFA
73xcSlWDWxlfAJK3ouFySvv9bDX36vxlNmzv90VE3M5g/MLTUzI7QSUGqnY7z+KK7QTxaDGrAbgm
RimvQSGBOeHnc8D6z3hsDKHa/YDC3izQblq83BMgDRoZpiLxcOHFxn+dsM68A+/gpTSMkZz/4CuT
6shz6OJ1NRPaLazhmo2M3aF+6esDTWHiYn954S1IjV7JVXt1AiruCShv/lDIwYAq0O5/yp8hLFnS
F/sUf/dh6q+g1OhyXSNqg39Ina2hXeEU1SQqQ2j3WL9hKj3Pw1TEnj1m0+hFhbxsa8l8KoMMsuvm
c42E3yoWRI0HhQgt1RNfN0Q8Smrm21qMbrNBOHkVB+5Mo/Kt7CU97C9pzXfpVw0Ofig+bFkwsuSb
1iFj9hJh8hwieGRtRtolsYBSSRKo0PCR/PIvxKY6Yu0FavnluJfWJCZPoUDEVk/yd7Qpuj2RNhoW
+hDNzpYH9j+coQ2S+FXxCq4/K0TWfp/twwWBqk+aM58xnbmaeGf734fBRQKwAHTNPYPRR9GVMfCt
yDoNpmFa+y6gdFamJeqA/4u0uTMnH0+lALIZcMpiJsX9yAa1ibPWrWhmd4zjrZQg6tcu9UGc3ARF
b/UVtP6KhurNCGZBooJfddnbdorQa749l1JFNgCoMKAXbB//1HswnZsmatqF3DFt+XEMcazyjfHm
YoAerZPfCmHO19Ko9vLOE99yvrpTkOKEsXljMUqnzEG+SROStquW3zkfe3W0AqzBFDendXci0HsD
oPoprKUthizl2fC+lh3EdwMOT54UZwIFgyPN5QVK86AOy+P4x7j14eA5SVe1WJIbhBInNTAwnrIp
qTZWlNuC2F5OwGnnzUoqNcfPYRht2BgNqGPE168YCnZ+NuZPCMqnxRO5trBVVcgrL1+3M1vood8X
HwEANgCInyG2XuNcnARDmwQk+fJwkbSXPFLOPQMOFfxavuGVf1L9tIfSXYhkfmsZG224ZMfj+oFz
7o8Hepp+XnVyAs2plg4lwURVcUg0J+6VNIIHurBOUKq4ZwtAJjttGHXZBDcOiYGesoVwmjjxY+9Z
fb7EUdCA/O8fe+RLHu69X6E18Hsj3uh/58l2Kag3sTY/4cog5BfQ/Zjo1iz9UJyDK2zBvE/kaceQ
rMspV15vcw7rohhoxEMmMCHIylml7XE4WeBsU8/XLJz2QywrRgtOsxQSuaDkFxjs66zNgsdcU3Ik
+ALP2a2vhRL7a7s344HOhDmMQuph7xI924r2G3Kd/slw20qwbtY959vdXPDO6zU/DJKF1oTXFsXJ
KS66nKohrTg+YD72MhDLnHB6YowDN7XX1fEciZt1ycjho5wbXl7PhmBoad9AOW76tqFJYL28NHV7
YbrYUQYlylFXoPv4q4OWJ8zFeLdpapuaaJ0k25z1Nth5rAI6++VPACkdakfUpKYyjYJH2b0WH+j1
TQKJDfJT8l/6Ev6SoVkhI4/8RJLeVxk8bM8+0WNefYHBdSFGXzX+pk2wD2UIn4hv2/1bJHsD6x3E
3c+mXG2X+xjcpyq68wzFqPxpYE7hRU9iH9OYmZCqfp6N0wTlEnBJvh7n9pONMWqV6nttGEb41/hp
NObCLKy1D3CM7LhD3f/wrtJQwUiOU+rr31Guj7UynwcEhrpCKBV+SxuyxEztiP/qIfAGZxCZMO2k
Ss2/m/JB96XEoFgv/MG/2pMXN9g8luElt3z8NovnSFbRdTNGAXArDgqRUQ3HHAGNYgnKQVXgz8WI
uOC/3eKQB3eAwXn/oGW9utqruRhlLxqA98acxNEXs8gbEnf/tcR7NmbngTqe6IQX86c8NwU9SAKt
x4niL5IVnLrfOpJI+yLqcydE0e174uqlfQ7NqHH/7aIaXFPwUK6oxFXLXLF4ZONR2GuKk//xhSy/
c0zSNm1bQLytbfaLoTmOtO8txYawlVWiDyfqCkepBDZqfufZEdJ4CIYuYw2WAVg9e+R0rposAu45
xNyElZ3EK9qs3OrnnX2yNd32f81NpM6l+I9YD8/nTPoiAH4OoYgq3V/Z8MqppgL97kAv9xDbt1b2
v4BzgNPLsCND31pfdo9AoezXEtw3uMs+7tz7Dcq/zqlW6PcRKUs3YDQb6xx2t2SZCbZNIHLL0HTh
1cRHSMprL9xBNh2Wly9JaIlVKFz62PeY1Rims9HirGhPbqTQpYBhMpFdbnwrWQOioRgxUV8Jb7vM
WGr+vYs+fLF9QYjuO4EUoNgrqxSbDuZuyMDlwqomBR+iCmHqnHhP2Oz9eDyPwzAiyfk7sud9nTDY
px24PolplagkWA6KmHvcUickGzuG8awA1eTzbO+MvSvndIzI4qHpsAGQ9UZPbYp0gycslaihaud3
cD9WnNxDoa3Farm5bYF5VIIYhbaMKW2fbC5iJXouEgGKMIMnomfvKQlbNSpsIzZf/S4P0iP/RkCZ
RyTS0ML3YLpL/32858rikdptSmc0C8yL/wNFLdcP9e9aquewTWgBYvbBTXbuuB8dtDH2w8/InmHW
lSgGTDKdIfW0KlkrfztSb8xYwW5cQml2OSO8Ta2EruNk2GuQ1c7JmhgcV+kdh9kN3UL0UcGSnBmX
Ee/zWNPqsrCl3DHYwII7GwvD1rEnFMO34lZj3r8HR6Et3VRFJDyig6v2qowP+SQec83VqRz/kjo1
yRWW+7S5+u32zn2EwObbighpZSlkS32UI8EnJ3aiLSSXpqs0+fmQHXjvT/myiyJ3B0urzC7kxwDI
3EYhzulK+tjxt34854KJsq31f+nD3L2SQeNMjBGdR0JxJOpi30of/3QVbqroLasSfEwhwQEdfAkq
ofQNHEjKRdQAtiQpzxNyrNPIlrjXzh52BVdpfHVShHNbGVOnHbejebiMwXUUG719AHm60H2jlQsx
g35dli2ArfG1LwiL6eDKsB7yMi1t4Dm3EOIaEj14uuJfxpzEj5DM1r+mRqdt5H7cVulgW/INxhSE
LbFiJLHUac6roOE8R9g8NcYpfZwqqXa8oy2tltNcVMsnAThJL6eR+XGEFXWjfO5QHjQxBx/RvvPe
VE0ozsAWA0oNGjOoxT3NZGvDhOi95YWlI1eV3PltSBIoxXnk/ycykTmPaizxSVExU4XCx0Gbvq93
pRwOaw2B1UjZ9fX0cq6uPyAEMsuS0wHosxo0TSd6QiEcxVsmHnbvjAZn9NBpbzGV5lc7XKosl0ob
eo+MyIMcZct22tSx22HAYBfCP20cr3zPzZrYcDuAc2lhR3CK47+aPnBLQQltpG/5JNfXpHuziYDe
gmqqP8UyZlnReWiQcIQK6l1dOYc8m6HfvH9n6Myfys3jWDlG//8X5+xZMDExXlvF7AaTkh7SHPgD
pnMMZ00Ew32LAPoj8MihJsFYIwYrW1R1h+VzT2nkijqU8DIjHYSlwDhaRVdg4CJrOBA35QFESxLJ
YL3gkron04ptktny34K0dj2uKBfvpkm8JT+oPfNmroV9/mkAzOgXQPxY3M4WA0h+gDBXzKc6On5g
VOaY4ADIWIOeeg0SxJMFCZV9GZtPtBals3KdRaLwW0FGCQK5vxJHexk2uZAMaAIoWEcANwZcpOE+
YJ4YNT2pDxEhlm2uIJ31EBLFNlc4rwW3OOpViWdiUjymyQRfsy53yOdD8Ln3URAEKoU3tNN5pEwr
r57vRL/lYZt1WpCzevoAw1M8NYr1PCnPrASMHG/wSh3oP3JCGG9VzkUG+WfMhVd/kXMYl1QriFdM
Y0+t31PlT/eC9M59joa5pL2HugdGxJC7L6nKzmHyNQMu+P5YMXKC1JB4wQidlNwYoPpV1aybMaSU
JC82OA31ZHJ8KryHZ/4emZ/7etDM5EkhuFfLJB6P7tNquxQmAr9YeAOZwZtrkFQ3zY1D/1KvyY4p
r8sjDlnafxJvYZX1I+d/kNOKpzQKoPYXNONtT/6fXp2CJNP8wEplIpuzL+13lwErzStrrOC50ByO
stWVzpCiajI/StwDx1jtKfLrqDrdn6vjtCX+hWrTrVOvo7uz/uQJ+voDz+2V6mIOWqJp4E9jfECu
2ySlf9TmlDxdJtFesO5H104SBrTDwQSO63AuuygJnSxVrkLuYi3A6213gbtEF4BCO6ShBTJAdUHS
NJEGLn7gckDfeZNL7cbeEjIYgWIzqwToAn5kmbW4Tn1HWWVNHDCdYh7FDjsLvUT9wzrxjgulodGu
k6h4gT4j8dYeCzRZjs7YhZ07670CTrr7Onb6Kx0M6EHhjrICBwR9EiZQriEoWp2jnAkK+hOIgw+x
a9qnZYfva06x+VSWMS2/CnHxR0DMrNBHYU7BAKsGzrnxSc91RW6poKDBY/ztimE7wjqJuH0kZxRO
INu4nknxXy95gc1ozx7rxenlPC6/m4m+q+wrIIH9KUA4XBZ6ADvPpKibex8RQj13OuRTKmZ8H6Ow
TthUWkMbhBg/sQoOLtMVo/kULZlqT/jv4wtuky8ZyMkD/JVLGztJPq01QnxK9LctRaj7ErpwSfpz
YHf15b1ie+ojJiiP1UO2xg4pUpoVrJ56imy24iOL4cwbcW4/+94CkuIynEcTk4JhxZNOJTIqC+Qf
nuTJGKGCsqs2d0OmoXl2cfBvxTQJBDnYYh2BhEUliGjsOVBDhyIfFk/t1RUgA0WOrZ9uSed+icJk
+b6Pl+9kHq/a4KYrvgoF2xQf49ACj20ZnCXB27E1c+2a6pVfEtOUV9MpXsQ/jEhORtmCE4vxfs0B
h+CCYxKqOkd3DBybJ1Z+6NPhb91dsPLD3jw366I1FT1tiaeSA3FPwVA1tjWjidCdEmpGB/6sdRu6
e9ooQsKCXyImXpgLVf+7KF/3KqzznZnDFtK7Ha6lN15zwdQxQmqAq+xlrnb4hhX3OphUJP9jhb7j
5C0eV52+FaMT9KYV8wH5jirPuBFOF3RJSdWPADLDjOjyswUuVCBa2SGeEdLqw5DaYB56WncnpgGQ
55Ge/yOd8ZZSPC7q4WadFZUS8lW13W8+delpfiKwotRf2bGkiainm1CnLuIYF2rtYE8v7g9ryJ0/
cFeq66aWTo3uyTAMeaIaQutiTmcTYWlcHg/Y/YJmNyRp9fE2+DCXG+fH87e/QzLhzV/dBU+wdZFK
FEE6keqldopXdpfzz+T7hRErgFkjZ9nLw0RzuquBJQiTn+0ZnqIZg9vrrpG5KfOYRFcLSG7i+vjt
/o+Rrp7MFBeXbZqNgFqJwHRT94BDl3vsg7IvXK/vgImrmIHFr2dlcfQsGp2Mv2s8x6EOj3n8yPcK
nr2ZKQrDixiXpZ/sMi1zbIFoX4iVPk9vSYtlLZ7TTkYLdeNKZNfSSfTPsYdrLBFGVlV8XfK1EpvX
a90eWrJ6mLrEWbuKRbDWO2GzXRJis5OQN070G+Pzc32ghn/IRTlw68euM547Tdgug4Uu1qDaJD10
Gto0s5cjGFkHlErv0OsBeut3Mak1TyAlqx+W19wR6A5vZuIifqswzA/uCTsbuWmS0FZkz3Q4DIT0
OXWdutJqT+eL9pAEblID08TT/6uzU5ur8YTzlfIT0J7ITizQrNoVZNRZg3YxqAbT3XRca73MyIpG
wDsLlewogUNwBelLmo1fahz3GkRyNtY9xR09iQ1crn2yCicy7vGp/2+z2olMUR1HmjNYA7n9zR7v
7eshzcHpmzkRjh+nUGhwWV6qZWUKtE/B3yIl9lw0iIhT20fApndrdADrqIZWpV+fEz5NaJoAgwqB
+YO14kkR2I6LwVnoWFbwoSdHkUOMQk87+2PPgAxVvi3e2Wek4ku0F7BoGxfqHbtPyZzFB62wp6u6
HYBPS8UE+j2MXm8OhcxEKwr4adzaHxJej8V4dnexfxzJhNp7hUeq6m0jSBPaERCIEQ+M7UpMChod
9gtOYSI71aITHdkv9l64E9NgrkBv8PhC1IUtgjkVybvQtPfooSugwGzgany0rwoCmnz1C6Uhk+7X
9DvP2kPTRXVUh0aViUrUWV/GluL/bHbD1lW4XXQwFymNrPIxIFNPefT4DXqqPsClzkX1K6sM9Unn
j7TgFejuXuntV5mdHE/9wfdU/+IaQ7WY4rr12PJrXJntcy3PHNeLkZn5Io0vu0lzTxZvfIWdeQ/v
UQwTsYZIxVrQPdOJEmOCZ4AIMiHq0PYQFDGrDL5kH79p6mwhGFz8797vvdQfRXsc3kw9Fixj9Wxl
Ho3Ki25xNHb/oJAZQobtm8qOST9RPwODr7zDU370DYIy3gtsvRXbxU5ZrroAjLxUEOl53Ayba4xW
W/4uevpXKC66hjA7bXpJQzEMBkeYttbvR0RC8fmVslxzi07NQAqLoZ9L0BhzM7x70ayB3XfGw7GY
x9A5M0OH7NhwhMXFa4qvFt6MIcTx85wf4HuD0voe0YhRIVfqTNNeKFB8nuSxJAO3hymAqcc3Kpkg
AXrqxN/KH6aI+h+JiAgMiH7Hzob8ZZf+kvjMiKv+EImEfF69YIO0xv0O62HyoVuFEstZflM//bX2
LqzVj58eJyKQcI09hRGob/O8iUu2cJnViqPLfjYnoyw0XdJ9vXTLfRomzL1eCzes04Ss+JFdmuaN
C6PkFMiWmgtLoj7YiorLgJdt80XVFmhcg5x6m4jSRqkouW7ya9nKasIKPHP4ICBSWEiZjRFlK8kO
LdrEcilFYhAxIEvrcbo62QbdtISOvoopipVV/kr1HsJe1STCK0fyDaxQqWZLKTX4dQrDlPZQ3kvL
HMlKNT0G8c5uLsUPBrIDMNdBfgkr+UyyWDBKkoRVYwSI1X0yD9tflUPzDCRMQsveYe+sVAfEdEG6
6iPEUkxOvbmvGc0lwiKBu0uL5yv52VG5kfKAKTB8UMVcyvMgTFWCJFAoW1hAoppXujbb7EwZuxqc
NAL80Bma4UuAo9FMUR0rO7c6lgWhPndiuY3TMzvrXYtJzo6WWlN1HZzoucJenuayM440l8wWWFZS
wcwa3fFAjddeDGw9AnCS+5Aw0bAY43jQJO5JOUDmotVfXRiREcktKG3uutGYQkOkA1PQKutxwx8s
YEi+oa2R6hNm6x9k6gigzgeBy4brsSp/sI+Hfz9Ut2SnCIWcXwSVOBxEsfBRUfd2/96gV1hzOPKa
V6FHNOqK67xZDz3Nl3tJq52vueE2gwZuzWSc/a+qgtTblmOUOFGQvgJeKTpNfftFcJbn0x24Otja
yV/DhHnA5QWewJi+Xmi/pnb+6LpwERDZoJF7AiPiaFMCUBwPssV9FiPnWqtfk07ENDJPtCWD1CmW
cAgwMgIySe3E1lezn2iNVRpcS6VsS39gBra9/Nnj0AeWHlVm87aQuwiJbqyxCFMs5eAsxk1kF1Ij
dO42W5dEtOSzlHZFbC+ZLXBWMH7HW/mSIOGaLHXXKesHf6PzUzgpkqV8Y+ao+GxkJvTQw77tuad0
aTmgwuhrwGmdZ54wCKYYUFT2GBrwG8qoQoR7+2di3yBIxgF/NJTsFSVA/xgF10jH1wzJYAOfrxig
gqRcF5B5ytgRvrW1da5m5JHo88gQFeshWia6FHy1Y1Q3OS4YypVWrtfiF5HEaP89F7lRddzIBfeh
QtcQIvifOhSDC8UM8STs7ceJnA1WpoAYRnyQrVC+K/Rdr8InslUbbUi+EQSmxd3EfJcybt4xN0ZS
F/VkAgW5JmwEdGTSLG1SiooYI5r4+CU9AoozopglS7yZb0j8GHPFrJOpW6ZRlrWuByf3GY3NRjCS
J+l4VXv758z9ft+Mu9YZfje8HcrHvdZmmMp/tb8YFYonwmRS73IHh/cA8i5g+hC40ax/SeaJwW2C
AqCXwoaMXxtTcmqNS70wUf1uw6+qXIjRxqy4r/6V2W3V+XpwxhDBBjQdl6QhRtWKi62dpDh5kfHO
2NuHwCeE1zO6h/xc1lB0FKbW3kA9AqO1PUpRKxE/8vOMHiF7k8s7LRqtQuBuKc8N4Fe36zez4p/n
Y74bFhw9chbduwuvL6yV7s9kWdgx6W0vO4U/ko67XkO/6ns0Cupcy13OV6LaIFmvbIwR6rtKp14I
EYR/GL1A9thh0qyLIYm9h1/saah9n0qsl7MgqXmYgaX4+pHYr176dFNxHPrAZU0cDayUIfgtmEo6
k7Ci9ww1lv6I40ssQGZpMf/qenQbo2C0hmRCGULRQVYeiVBNexomNTK281PdAvHEcU8E3cGnQ/bx
1GKhaaQzH67jVW7r71P6b70G8YXVDncyCZQe0HbRugwfb1fJUgmBcjY1N/3Uf6Wo/cbkWxUug359
DMvVR06nqd4ksq557r4+AmVlRAld0nKnMg4nxZvaF1PYW84w6JdEMKFSi5uHoZKmzEs94yruYuRK
h0AlyLwG+cWaL5j3nNkitM2a8ATwiyeo+BvcbeiDdh3PNbxuTN0u8k32JaHX4Gmz1ypyA9eIsykM
XKotNcUmrd/jgxveWQWZu79cPBy6GXMwLHYjRg9vBhK1ebDftU/W98ec6hUtOEYP2krgXmPaE8dS
/bAUV1CyQovYIPcYpqa6Pxj+TcVHnw7GSr//3tHIOcBaA+Mz4N1Hc5EFNHXouqB2MioCtao7KjVm
6Chq+aU4B0wTvH77tGrUT9Eih7w541MSLfRmtF46Pz2FgMds/ztCSiXBr3dfpgPSyKBjyldx2nSM
MqFMrEqtRk17rptwIJBsiUmesjvVCP/6842CBw8b0LuNu9X7mc1JMmb5gWAdPS9sqL6ADYKYXxeT
rIEOpTkzVAExkv8VP84YIiRjIqvlW1Dn7FeqKRL+H9wQNu7ZZCRyM+c4NoDeFkoNq4y/Tbp0FkSO
nJciC2Os/dUUwnaamfbHRKXmFdr4jNpkWt6NFTj2JugqWIeR7S1+rZfpFQI7yV3kZn7JS9b4MrsM
PGpc3GELYIamvjtHRWNxnf6gtMEBvv4VmhMsXwDZIX0dx2fwtkwNn6Rv0tX1rUWk49GPpAL44gsh
qpjvLWPc3ONu1ZkEtoKZLF+mArURUcR3yJfc9fcCG2DgVUnYIm+vpuv9yhvETEkQ7aBNFqp2e5+Z
cmkmAcv6arbvGCOPGCmFvdOSg7YQrdAeqvm9DjUG2AjDkl5XI74KdS5vT1CS4+GB62uUmQjLeGjo
J4MHPTiYyGvYPt5N9QI6+b0L9UG9Tg3CPuZi/5dVp6ODBRYPxOAi6fUpdlA+XEOmrDmyUYemu3qj
8ENR50ntZtAtC6ZF6CY/bDr1kAVabip+ORvaCkpZnL0sqONsmdeMbk7TnACIIr1yAy+XbbxKvJkU
cya1ORIa+yu0e3+zo7/1oaP4JQh8EX54C1WH3OH+qGdXyKuoX9uaAqmUtCDLeFAnLo4s5IMeq1kK
He2jH+MKz/B4rDxZGXTfeLS6dR8x8I/ZiMU+lRnPE4E5AlaNrQDCdib96vmIpbtgit4EI24ZCMUP
UeIg06n9jWIpN6sfEeZnTwjyyAKPfMWaY2O6cdZzq7+qQN1PAY8g6FWTNz0VSmSzPD1Yv2Yj8/1H
07T060wZzYV8UUIo8PubgsXORTstH/hVhLyCyqailvF8wD+f/Jd1Kgl46zZMvj01c0jx+ev0fsmL
hwm0UDE5QCK9Fb9trbdv+vLU35llUqX90RAC4KsHwAhRetoQDEPdovdJUnT8wYQnYMGosuESiEu3
SSRDKkpou/8z8M2MJ1yBk2+yiYICgtj4d3giUcwwQhycnFRU47KMSLa5TrqWDwyzVtMmBQjW6fKX
gWmkJKi1MkGFDo3h84qjnxlQcE0Yrd8M+7ahpBwk5UJTCko8ENWI/NtCZHketU5TF7Aejv61ajx9
aPpFqnjfZbUHvGjrKG+d65l/g4xweDcOA2j6xtw3gu4XFvXPsrqGyPhQ/RkuJ/zmHwUTPaMhzbXB
M13Mbd9b/b3N/1IwnqyRnHqT9FlVvk8P2mhd7xQZ4rw/j20JBCxS/I2bkdLPFLhSzmjFNqm0YKph
OuTPFo+DyTM+VyAyaneVT5VylyzW6zqUlep85TzvxB8PPuW7gFhPZ1Et9cikJtEttQarERzvQXIj
WbUAgVvPx5Nid6ubDnjPgOqzd8/sap62fYcmjBF5lQTGTPdFc9y365gftJS/peXs26S1QF6h4aKM
6JtxLzfbIpEaa51mfZIY6aycfcc1kit2RsiKi/JPqCQjMI2LWt8FkjtEEkxadlpET6itxq+B1LPq
V+MggvNHpKgJmvBbIa7+KsYI/xLOKkhhPI36TbJ3rS7BKqJC+tBZLHKIWpkHjgz1saIBBGkWltQn
t/7rYBeHVzpggoVV0sH10nNk435f+fGeQ2R7mDXOIYKwWgPC0un18WKlPf5Gw1AOXjbBayasAnCg
wRYrUWe5Zjs6HoEBACOFF5WXyUgPRNTvnbiSzdKT3DSEsC0FdoDSDpAY/qKh9TIeLyUJo9LV//zF
L6KwOZwOExNtpz1BmmhqjUw65gUzNqNG67pqy+jn5Li4qxnlV6rRitW17I0WcVYM2/+uEYkReqmy
NST2+fzSQNvwgDe3vjGKshCJrUTuxOyBDqLLyjDotCmWIukLsu53yhcSV50s/c842994SbI62zfz
UBSvyX+mSu3miKT47vd2tWEiwy2pKG70yefBTgh8wrd4hYb55BtxU9owGMPN/OZsTqjZIxtKMxe6
HBEmwHUv1byLLiSj4jd0V2NSr7cM8wNDSKJIHIDkf9cuvU+ZE7AaGfnAsUKNMOwAXaWBlw2MrWKl
ejKbc/9Q2OC6iayC82QigUNFDBMSjV1ixT4sKCAd+l9ooro8notN2UoQaMAT/UzlXkJyZNm5NDeU
HHUERRJpTRkaTZ7lO57fInCIh/WvUu9wpwRdGMV9jhhzRU5ZxdLTPuHplt1plSRM30340r7xRpLo
TASsgNSPDxRy1jNwk5yJ6jsbBOuNeNAXHUdcoaGs8e22Okg/Yf+lm81Su/frvda5aoTyFjwkH82Q
FN1vUUQfGIM4OalXxenHWcZuXe+3HyUEIEys077Q+OjQ/ZC7kT+pVaoLfpVwhGiFLgaUNYo58lEs
kk0ADygYNULEr5j4A0cLwbPLQW3ux5+tBD6oKdP+OZgQsobymCNW9vJKyp4ZraFxpkFStoqX+oxR
JWvT/DnsaLFFqYLnSXTtSGcH/bIrroDVHCkoSV4QBI4UAe9cJKWn9xRr8hJDwCMWadUAwMpPjbrT
PHS1hoYWswhDWbiBz2zthvRz63mPR1eLaCoFb/cGlIEa/eTi4NxD9pj3Hsex5A9OM5uzAko+S3Kj
IBzbV8EwZ2X8S+RMys9w/lTRcWXxeFuCLLihGaG3Bl/bu5oY1+kgwT5/71h+je18/PqAMsLks7Up
5dYrjHvZd6Q9BvHfOM4mLmpz+0riV3u4AIyYZrAKJPIMspJ/jeSwNH8mSxE3KAN3RnDWm4Z1SXO/
AbNoGBmzYDujb3RqQ8lpTa1b5dHUcAS4We9n8aQLtP+y+CiD0LmdRP/6O03W9f1fAS59pazay0YK
CDCBJ2uiiDFvWIC8ndbyiiOSwiq7DB1hXYTBc2TjzBKJwH6m6OPK0cT2NC+5LnKY0uZAIcJuIIT1
Ao+NoAWIFOz2oLnkrY2SlZK8RrU1Ijs+Cy2VkDGRro4IFp8Qo3mim5dsJiSOCRHwFCeTBriuwAg3
L85KMSked1n2nvjO+o0ofTKeSH6HwWzUMAnK5myQM0Vb0jrj4CkT17eZoLMqgFUJepXNSKRQf3sh
CT4LTpgHUiMu7l8uMXgvxujC+CMjRYv0eq3VueuQiAE6Yb8Z2SKoR8KOdog+b5Z7B0rK8LuY71PD
ldRHXMCvBOzqAHkF+XrwFSqlPbiBnIDxGrJXNNAO6lfPqF31UUFyfpAItrwxuOCpcEmvtapqnlVP
fZ6+xaMuLqPzCIBnIiTb1lWjSP5ezyA6EXe+Ci6HZIzp4o1g5bXDXDdPOofGP5/6HmG3WP+auMHQ
P6VHxuoRwYuyy2+GPJn/UEqQPPSq82dsVoHueGi9sVmJetJZ1CV8cYw8/H7ULoBkieXh0bKtHJVP
HCtgdeRkHt7g/nH782n/z01yNYzjMBkOOINMW8yPMq74MC0YaBC5y5aINiBjYFiycss0ustC5NOt
EpvMB6rFcC5DpL1g5M+8zqEhnWTqkpbrfGFrzmhqERCZEClOVOrJW8m0cNz+8uW4aQaRpcgbeZfO
nUkzyJsqHpQEG1Kwx7wciIFLSzWU2CQIDUx78Ykd0P2Ustvi89Z/ECV0RHZtd+5ygj7jnjrCahjT
NkJxCTLaG6i80uxAGvCxYo2dB8UVAnOO2S8iLcdZgG9D+5o2B1OAtfHN2OhRYnsb7if3sOymGekT
gIHQPUoVxDgYgwsI1aYxgEGPciwrBApo82xB455FPFTvQyQHpvoZ/uqR88NGyGlgHuW+jlFmS46L
J2EU1MI8trI8dTu0rwA5vXBzRncklwutUNDSdbnugckX+emd53SwTws/jUy8nXnJjCm/GNW4T6mI
rTEnjYbgu3zsEsN+uWfliaIcrPGQw0wi8jf44kpngiN+ctX5v+V4jUMjTV1O/SV2dCAwc3hh3BWu
wxHknQAO+968hDZa4baT2QaTVvXgdC1Zi7+3m18ScoxvbttfSTeiSmN/BvbY+DIGQB8KXRSRnlAN
4ViYLz+VWZJi2eP++cl01vMd/ZTCIfcFnQnoRcBMYukbRnb14lcl+1gs8cPKpbBcL48V4OgCm3Ux
JMwzitCF883OGK79eTOEm1/J6q/5JydB31saiw+IurnqKjESbeFnaW7EyLQPIajkgewS6X4B0/on
gIBX0kT50ngKmUk1VGpYO4vVC7TjReRQhG7rtcgXK43fQH+3zUaLAKzsom1Zcl26z0rizQgH6vmD
zj07mEKXaEO/Em7lOzQwQg3duKJ7Ld7OEBptewfpxfeuQqhSKsOMYAXS0Dm8nowMqUHg7TlYAsAc
tWZPwj99iunn1GVivB2DQV8aHJ37UFo4AwwCLT5D7clSoomm53LBy2sJatM/eFD9msamP5pUcRmN
LZHBIEDtoJyv5Q+ldVYauhNJLqUVO4wtpoNvKRgUXd/r1DPR4U16FRyt9QOg+UOXCAf5/jAizbGN
vqzPy+uLRrvEhe/hbhBUSjmIFuC7q4Zm4IFA1MVRcjYpcAMCRboEICbgnMRagvJDKdHHi6M0HLZp
QA4obuEifqU2CK4pZxSWfMtuyenthjkKDsWxdPGeNEX6yHVcEKGPralb0EEzCVSOLa4UuTOfKeFk
8F0gvx+5vWRFnNoi9EMKm3EdVWKL/AVcAf/LIIdqUgCtGZZ+zNIvFlx7Cc5aTEEsMCv5O5uGygWX
XtqdfFeQKrCF7EAEi4clWpNJzVN1eGK3rM63vfzg6OGZ0KscKN8rqzpKEvr5QtVTc+Y5nMPDNU6Z
iZ9RyfSpP1JBb8Xgm1WwZNh28jtl9187jKSggfKmm6Xl7q5j2r17LLZ5Ev1r3uWmrkMvKCmoX00C
ekGImS2BJ9NLCsfL/VsNQOb+tKdZGkeO2H4QtSYlraelF1CszOpg/KseMmHpXq2HmGnej6ZCw4VQ
XPMo5o0cLsJv0QnOrqFWRYk1WXY6a4MDel+6/jZw0gvOXsp260R7h8iy7ZCZNqrzC/Yw7kif41TD
I2ewu5kN2tpTu9WiHL86tdt64GzeW6a1c/NhiTyAWFLmm2EYUpx7IE8+1/5Zn9xTcz1ubTPcBOBq
3XrKrtcFizCGhtGsdC6dSXy3507apaPAnt5OvSkowPz22cKor2wu7pontb1GfAU6M/GqUF/eP/Wv
3rmJBmjg5f633HBUFJehxKBNUcUXihKTQzI8Rh372Pyv22g8f3kTBlDWdlyCtI54GLve0is9LMnk
lsMqNV4iDxg5ZyrlfmKPjQtTybKKDKvZPMi+m5wwXLLRXEiLsF7FgDxYQw0aX/uE/vzlCYbYVdor
6oIt/iJsG/v2IXxhZBYVyvTHTDRBeInhnb+P7F/EloXGmVnNHQ2f3XN6lVE5iuIAvbknLItJapjJ
Rz+MQlv2XJQbIavDXrnoc3doCiPBFdsSs0uWLOnWhqjJK2uuPQMLdQUY8Zzj5jxSaVFMshAsg9Ac
3TsT3JdOlDpiFmU0TUOJmzoHmjYoV/u2h3MVmSKSJJArbW1K5Ubwl0H0b44kvPzWwoqXjmRMNK/s
yUu81nlb3K0X7TIquLCiJow2POTA+spyr5Msnic7Rv5qDHzixlzyFsOei7pyQgBE6Jmr8UW2Rf8Z
hYKp4ZP4H+GcpQoJXv+msnOxs3VN9+Q4goQyVhUgFcrbI1QAJMSkTO/cP/+0ywfDoo6OGxHTnHQ7
kaKnWoJHTU8aYVC94hIOMVZ9xBI+BQHxNueePSP5ma2NhOtz9uZgJeYqi6M23HAY2ZyauQYjEpbV
eJsHvjJCKaT+H7wOGLK3IoP6x/Ry0Kb+WJJReayqEBwwrB323gOsJGcRy6OK9c/zoYOXfRp95A39
oHeq6heQwFdpGKMLcibhudwxGeOx4jX795xZJm2wo7BSmpdcJGVm9RZb621uOI7zijW7mNi3QqT7
I928cmrUnoUtNmECX1SYLZQGLW+pS9RLWtkslPH69nMFNwpQG1ALAEneFkPajtCTMXw4jK9wn+Rh
bMfSMDLkYwybTfJI3OCkpC/w3xkUN9B9+2wE1/iZUJ34thRDnr8RbWJ59iSQofBZKemIabaJnJU6
Wy6Rdv2WZWgPC/hkMwu7oC9I+g4jDC9hJOCVrw402kgYCfLmXN50gSDB4i8h6QK8mhIG8k0jpB3F
1OWtbq1ch9RPFuvfTNAnfZ0xM+aX3x1j3laUTSbi9WeLGLMu41ag/voGtC7HZVQEAYnByt6sBJal
tJZltt5G2uwxWh9AoNRJbiakuFnN7cIVTDsRLBTP3a59crj0S74zERvbRBcLYh+UASHH3CyO7dNV
1mOm68vvDVEGE8onvQyTX7HPIP5jp5HzmdlSPVOAp/pHO292MTXR5PK7q02ygEqycitoKUO3MZsA
r/1erTUWeRzWqgtQYPlNjawX0/8me9SafkUVDenZM1sT2pMICTZ+DUR1c7ZAtu7Z0qOumtZ1ttwZ
tHN9exTCsYssc5g2wQ0Fuw9LxCZkOZKGc0BUUkdQY6aYLPCNkWZxSMn8z6y6hCh8XcUgzMmtM7/m
cPyij4MZmySawx06WdR511IHtm4SYFcL7DM7zPC6Qm8A7R5Q80kc//qrMjKyO0sh6cp2rdXOP15V
jK872uueFCL+QEdMnaDLZlVOo3xTo0ymaGSTS8KN1PUIp3/mAXCkww5rAmCb9kPuOoIWlJgHtf0j
eQT0/7+r5Z64bA5NOasjcAr7LpCUatbaZRzqbwZIgVTKI86pvWijQat1lH6ZZTVG/fm/YgmMJHff
OZUWzx+s9zpscMegQxFC2PiSnmQ2aHHbAZy5pscW/A179uzLOuQpPMbtUUlg3CsndJ17L3wq7HrV
TKc8m0NIfM+HkSiHj0CLh78ZUpjJVz6iYnL1ft2aQZazbAQlsoSp/Ois8lhGGvFsXw5SBPoQZq/a
9iwQ+JxE/7pX8Qq2ljq/C2hc+RyRgDB2KZJTCpIRdkttwLwc16qIffcKTp16dmjTqScJB0O6ycEY
+dWGGV+aT1SWfH4rMZBIrhdkh5fGJ0vSWYXq9Z8IPj3sCb0SawQn2KXp9+Ma2KiFhbKq1cbTTur8
QjTd56UDUcq8UJAhoZ5kvqZ/+j/eB63H/PWWorhx+K1XbLT9/UAER1Xux9/MJi4WsBgNEOa6thdQ
dRHfRx7RDsvCmzPNG7DX3wjYiHD8yskqkxdUduNu6dEWfof4h6/FP28hCP0DyFmWSwL2Abp1d5Ka
mACOkF0/UZQuXwWg06BexPD/zABmLSX1rqLJapwtinKx7DQfhTjOOHmP+up2acQu7DNWGQTpNs1+
MaShLVXQXC8J6k4Nesez8XxAAri9CaSti2Rxx0dsmLS7FY9E2UIH0l9XY8jbp48Q1YYWB9C0slwN
9ksEmYGae1QDZNrwgspwAs5tU6v+2wTDVVyMA/onItndaI29x8YK1i1ZhcT+snfHlYlTG8iFEzLx
OiHoi27u7JyReHarR5dUmRbREl2cBZtvOJUQqDuu18UPZ/U+2sjUX+Yw014w02e4qU4Ih6v5BAVR
J8tEJLQo/37DFNvPnHhCqXi5nqfOyYywvhf2ti61iQjCp950v4fZLJcuLPEBAk5YdY9cdyq3qUfz
3srRDIlKbuuijnGo3GRWMhptDAnP8ElIzddutTKaTtpI6U2ktybB69Ta+dRvSQWTTkpMOoSVAEmL
SJPWAhONGtIOjuTWJvFeaD9Rg3gSy2hS0FRF1wlQlYthoGw5BulwAVZsfLrtW8p+u+Kp8zYZnkNG
W/dg2ewbc4SVXwSgofQs15D7a76B22w4YrDEb9GD3dGXSFeelk+it2DJyaEmfkAlg9oHKcefFShF
J23DabqAHoaatCNkbEngivll6ezd9u4LPzRNzo7oXI8sar1L5EZr/d3b5f1Tknw+ePXOEspqqAcu
4nscSqI27shAneRKAN8Ej6jtXqiouc/9GYhAixt6ek1cLZr5zdrRjjRXQ5TePl+q3dTjGa/bpsRq
w/XFuZTYE+MCgC9yUMJx3W76KuPq0D5E5XoHwJil7TZf8XJxupntKQh0QunzLJivKNoMypx1q5NA
SIpmzMr0pIgS+N72F7LzRDuCmypKhCqhkM/ijjEbnneXhNigbLOVgVNVCKfgSTqH2Tt7JfuAKaqK
bUZYy3dgzc2a79HfwNKTxdJtRCKBE/XfWGTrtyQTsgbg4BRTH57OwPyI6a+7eWqZ8zSX/KQZCE01
fz4pzxpf10GqmWleLCXeW64EaQz1P5LzqKxz2R8PD/1mgKz0eilRFXW16dwSbmhYToL8hdfHRHtp
i8L+/d02dJ3bPk1zwwaRwgyzu3c89CRWCLk2W4XiqTipyv0hnaJb8ET42cbW4+xzidJVdcU3wRQs
JuqSv7aEQ7gWNmBN+IYkDh8ryC7JuolEealzAvDddBY09lCRBYtxIS9B19LvP4fX0glWxzFy0usC
nABhbzqEL1MDyB7M8u8938kG2mtnBXr3fi0FYS9Vj2k3uwaWoNDHOWnzfxmIwMTw0q2OUoElW68y
2+hpBiFd0VtK+VL9ZQ+XgVuV/sMRxXF+GmpaMAbe6FpkubpmrfO0ESNOlxpUz+zOwTyRvrS+0I+I
hb2z+MFRN0gggNkrPF4xyuhPQIYw7Q8tjGJRqgzvgzLhAjoU5HMlgmgq3xwB1HwvOoPhXvVOHSJ9
rvuoXFJ/JyoRIf/QTSLzu6v6shnhF0E2L55S011SlIQIKwKzwfM/bDZln9L51KucazPRIk+nl4b4
dYTzF9vXgEh2SP2NFiZaK3r7PU5ed9Hy6D0c4U+INGBvwF2gPINwecdpBuetEc8YeEuX/l3KWIue
yCFwNztINP+lTf1lwmbp0JSmpwEXFvkUK1AMZIcUaNNRitS//Yf7+YUrfTsJuG9SDNSQqmyxtQDg
kWux1Oidj+hvshGVHOpJFA5yjWTbuvMoFq8YHH4lsktq6klGcNNrZLrLoPulW957QjTYX0BrEiLG
Ac0K6ZhL9Y8251yhrWOsa2UZq6P4d7H2tOR6CaYZP/h6uGJFskiMCLmtYU4IBYyC4LOl9MnQ9OZn
qEjV4RqdWTa4aNiQwDNCE1iN2MyQMZ2Uqzc9n4LyAXwhu24Hqz2tZv2YMIgVT9fWDA3b3eqrXcTu
H5J2kjF5RREyT1yJmJyvaD6UoUC21+2k9GR9wbMOga1cOGVZKeuoDbjaBL9Nb/eo770OJduvE/A9
VLK4FzWn4NiDgNcxon4CLeUoz5RUZh2k/bor6k54zYn0kt6aFAtZ7IDtzETT4TBGc7keG/ARXpKN
LSeItYI+Nuia/g+0xcekP8tI81tSYTtBBH+WzoEFsGuvbytBoQoSpaLWRvrkIOd0xq4ES6g4OrIb
gY3a6l6O6V+hHs9eQ7kB0YnsFb1cYFAah1zZVr74qgw6bxEThtjIEkIreGptXBDbJThYfbhwYfQN
ypwhY6JBiCCsf4GUl3yObkEsgJg2b7GX+ezBTpUMZOYJVpAnmn9sbkR40UqhhG+iTWwu7DH/Gj28
WTQkBdZf65iN8WrlJD75eKNyeUQ0ZAdiEMsDhsQd0G7TX/cZafY9gGrE7t3TyB/u8HCYnzbUAah/
lR8EOTqLhJ/mcEQaa+ofbaKyxY1vGT49Fp+/Ps6J/ViCNqmOaneQ2bgEBNHSDN4Ix0Len4njCzuW
U2ARkSGNeOcnyljTH9ShfQblqpQKyQ0ytrl6tM0kLHLBpPwWUJOto1hJW8+LTYMb8PfP1S2OlnGh
PI5Gd4yPayr87LbK/QP06mMNxfCC9e5ep2qpW3GiUTmvP4qhFToVt6cqcmEKPMQfzfpsmxInjwVp
piKJ8v01h4EpENoiVb8/sv52VpxHdGr5khLY15pnsGrBS+ol0NOrMbFQqxANFZlCAVV8CZGUpkDl
cGyqPjQiD7XOlKCtKfbnndW5jISQ50OhnDGQidmuI6nojmM0DwbwZmkvpLSlVM7NYf2bW348JeWu
7NfDXNWTQDOGk0hKTaG3/gIYGQJKJM+lmNt59tRakd2M1iBaZSsmDyP8tAEygccpWhwpzLE5uNZQ
p6f0/VhQSuvyVFLzCVHN8h6l0cSc1UzYgzUIV3ApORn8v+Ig2+t2yPJj/f+lM47tiIc0txqQH54T
tf1JSLWa/XxPrh44N9CAW6CV+Kp3lsa7NZQRW4wEgNy/OjCsT64UdMZlygVqxpyHgevCPfw9Ir2H
8JjpBcujswvZ0Qhp96tcGr1xGB+v/qM4l8s7NedzZOb/5FzmYtyIkyxiGUJhn7VCsm4TULLW55gp
cKCgC24JBWf5HP5hGeI5D9SK60MsUozC/Ym6NxTQO4qE2RhwDjK8lhJXQoujLg2evYb+n5JId6nT
7QPO4/+QZRjdVigO9UcnuCiYcGCfZBPfidznIRW19FFZLcpIuVhdD6nZtL5OPd/3cO9K/qateBqK
sAZDhbJGs7lPDEN4jESNNsLZG/tsE78rUSpNSYB8VeNLYWoZ803SHv/OKVFKfIMsXFJkn4KSYbfx
APA+w9CcVnQLpSswISKxwUperlu8zeaUXLYDju7lolsiXg14oTr9FWgsJ3rQ9D/hoNb5/1cP+5Dd
DFQWj14cWb7xQRbUWFSUVFZmSLXwxvrVKpxvMnD6oah9+uTCnFw4pJrI4jnX3auvTbOpJf6Mgkac
NmfnzCcrVe3D/uWHaDfxUezdNoj3OWyX2vhybunGGJ4DfDFsb6p3Xn8nmV0ESUzO7zb5NOW4vPkd
KMYod9yEIDItYFshzTyAyW+ndMWAeWt1x7XvNWtMJhDCyqCuObjJN+VFbZc97yBnv58108FRPfqw
B2bjJH8Dzg/uemnhI64tzSJY31006nIXnYvIOATq43S2daPXdR3ESv0DAFbUiyfiGjpIEEb8OAOA
SCqYJam3k3N47gg36KwJGE4F73JYcx7xHRBfHaw/MzsDgGPUarcN7opQGyEeRoefNM4TqihhSknn
YzLEV4BUIl944NAbc6L5N6yWZXA6yi4JQx7CC2FBwSwvtXRBfmC9HZhHKnZn9ZfWYTVd6JzmxP6y
YZss+oq7Tbdc7W5ZRBY2a3HpRoHEmH9Zvm7fbYNtAu2zCt4ZUUN/v724mlZKExe9NhPqK5C7bM+n
TftajpixvTxzWgqibt/D4r1wzU0xQzOlm+4TQApsKqK1iCPnifiqcTp8emF8MG1fAAceSFC7iWwR
jOBP00y0vlJffJeKvgaxyF80wfHhGIY034VGgJnfJtGYc8JJDCRY8di86a7BIVNdmv4WyquqWYYb
Ya2pIi/Q1nyoF7tkADfFWZSXMynu4WdoD4cvCJDW8sVaE9isfipin5miXcQkOnNZVZIWMrr6Uvc3
Abde+yU8anuZ4mMFSiTgfRSlV3PM7z3eVJARVJTr0MPkwjwNLl19tpfHiFFf3prnVWqVCZ25vqot
pTnYtqY8XZf54gvbGOnIW6BtbxsnL+ZAhyiNJSV0Y4PhiU5gt2LPNkdGlsxLRRBb0E8kYu22H+ua
Zoz+n97ASpKxScy4tm10O19i3ZePzU5eZc+q++/SZkbG7A9q46y6/Br2HAEhJuI7beBWvneIs2IB
sowG8+rTxX5KCgyKOL8T5bjMwFNsqPEFdCAsWzp4cmPJBxS2L1Cq1UIsy8AAA6aiw8RSNaVd6omJ
AuijPtewuZEGVaCC/6thZ1K0nXi1fHsmHEAP/HiuKw82pxWafyTu/kuR290X09W2Ys18WkVZTvM7
Af3LeMKhp+URbsSZwLKFXd+pJGEuOQP7vTu0N6dfuGHTFnwi1joV4YC94jAdAhFOPk0eCxlQpHkt
oA4NUk4wFApD5BHDpvkLHVjW3/kwYVKI0jgzTmKrnZ7OWDqvI4VMXiAIFoVf1igKVIwe4DfLyc8B
fi5TfgHUsDrzT7XxDTElFDAsKSAyzML/JsC62RgjaS4Q3rSq98wi+Yl8tNMql+j2jKQZXdnRdwZr
byBEJlgcMt3REe+OshdDzG4Q1QwyIFJNsX1ZFexVArRAV3bY0ApaUGyEHHxkMeBoKoWZgtlD9E+M
phIDDTVxMKYtbWGwtAHUD+mJZwh44sFy6azd07qzprCr1HKP34PKq+Fot+taMbManwcDcjUn98bF
N4a06k5ECrRa/kXF+SOtJR9SE1i1A2lAUUqAPi1cTH0Yzwk9zzSNncn/RF1z1X3QQJHkoCb6Qn4O
QQ437f8d6s/XRZaHpFH6t0BlHPnVA6zmNaoJ57gHXxVjqtJ/ITKMq3lqo63nec5QtIVzQqRkfZ/6
dGKh6bKswsYStgzuB9vLz9nxhLPdaHKMY3/5SHmyG8XjzkQOeFtN3ffrIwNCnGOle+gx5RP8MQSH
VuWotLCwp9zu4mtZP8otAc5VzhXCliKX3UmH6/SvCUAFZmlW8Rx39ly8dydFLEL1o7sGrbnfJbnm
IQ68rTwu4rGZlilkhfzvmF59TXT9LxpsL+N81P/Fy8su1gsaptGkSTwS7MfOBz4zMuKC4Sh24VTd
xXjFD4ExuZWlgsMzlaHYF0IVqyKq8g8zRmPxnL2iTsPrD8vc3kUUfMVm4PfcjtEnHDHAyLwwKGUF
Uj9819u+x7Gakkn6lf9lLw8Rk7Sj+vuD8iQPCU6QdGiS+Xf417W7+MTVpLd9SmNyMyecVyejq40/
1/vwbFS8df17l9h4KupW/x5MoQWBqeF8t9wgQF43cFhWkNIsrgnZ62eJdjOIOD4kv2aTHTK3NDWm
DLxRuigk9EanmrEVL5cZ/wXXvgUIC5paDMCL+mSh4vA52wuRWkhGqOp5K3XDD7ui/Dn2NsU5K4wr
pEJ//Bo9c91Osmf0SLdf/ljaDHmCB8SS4U6TwzN4XG6cD4frfqN3NgH9cbXguurTVGUsle/v5t6T
Q+tQY98robXe6cIZZS8VO1KGIlb/iZTOAba90SXeV7ukeTcWzKhRK73OQEaceUowx/627PO+6JFT
DOYgvgBsfkRPPt07lYAQQf7RvMSITlUxRXy6aXvgd/ZjAamMrs4h+TS23+t17ThnCd5BZx2/eBZM
4JBClv9t3+MoY361T2ooKJLtXO5CCPRm26FKOilpnxiSpEx1hzVMDJnDEICpe9QeA7vd2yO4v6vs
dxeJqlKV9/GwTN1/dQ052eKDgoDDw9zPPdDNdD2CvA3EF1DIAHyvwQZZixRYoTaSacsuSHGrpise
DrUpL0CqNCJMHI+Cg/nRGDquOdAhmdybIlBvmwGU9wWhJwRM0FF+OLfgQdh8kMHoNI9N1PyZTeOr
yNSbU4CDq6XalBIhcs39n8k6gtc0UGKc2SDQAicdRqma8yqBuiR3/W8aDN+u75V/1cD+p/Sb2VxB
mZNfzn3Hs18O9VqmZ06sOBXNNnS+L0BqBJZTQY6FeUhiripQ918pORWGgexGD65gZofMN17sE/tZ
w7XZpWuWD1ExdiuubGjhHxnh1xRilmyo23FnYTha8j/D/yyM3XBazI0q9UArKZpjTFLVrgCBethu
odKuA0xGG5+ikSJpsgFvxKpe1MIEtHtJCYmCzRry5F5uQ+yAHZ1NON3yGEg5xmUtJ/K+2KI9YAhW
x9tUjncGae5SVAaJ1yp4EBH1GVIHKH1SrFx/LEP4XIwQAQTK/J982NxifwSCUBmP01ErNj1JHE/c
NZyNpRvMX8bOOw2YziG12/Nc+It4zyZCuL+Hy4a7Ul2H+cyF3XaXMLWDgOFq3Og+sLhlxSXuVHNu
iyS1meQ7TE/gMdLENl8WinP+tQv8ewdY2+mNhvsV1dBMiiLIE/V6Bczc3BuZHTZL7MquEk5yMpX2
z0Sr55wAy8FtfXqd6p+taq1jdjIUVMQPk8ETzCp+WS86QPzateiz1box9PTzm3qdNRPtRzMdLk41
wAu3kwwb/oLrRQIzWGpsyupwz/3lcCWV9qTWKRzq+XClxQlsXyfeL1g0TkpkE3+aVfY0SOwflfmY
cFG6b5t74TLhbuKV8hncYvWC7guVZpfU5wu3onQ/WJ6ahWrdRZKyYCRjFG59oLK9ZOjEjEb7ZoQ1
V08dHDnNHt+/4klzCDkrshyzacHa6An6TGyyWD3VJ6SOsYq2H4Tb7VGb9QiPUlQyG6EXpECr4dEG
kwGBGMNF4QfREA4GQYdpTH9mORQLNxM2/sS+wM5cWfcXRR4LHMWGBY2tpXKDQRNDSKJo4IV0Gam/
Fabf31eLd/HWrPLwacXoj5+qnP2IRajblm+g5rvBPynIIeWdNw8OgVFjQK8JaiN+IlzJT/K5zvqN
udwH2zHOqxPOhw0ZCnKUfd7uaZVW0gGBG9dvTn5qM0JRcIGlvIv9GpQh/ba1hsfSdOGQD/wB553M
HPASGWm45nrSTfXM9sPkVuAFEMxADKKENTuY4208NpCayXplFbBbNQUb1yISHS7Y2xinXBIsPbu2
30XO76YCNm7EtsAzCLD2w8JhnKucg89xy14u5bZFQ/560DINl8rj1IeLaGbH6mtPsO2olfuc73Vn
4iOAAExTGfyZ/Eq5EtUS/Npvbi1jY33hVKXsX/d+VWQjUzAnWr55WNlEVQnXVVvvJVaREL457U7g
+fPa85d/IH3uftE+GBSXGDRQTNY9GPoPr1NT/YceaeQAYh00uO0UMFuJWcfIUGwqe/gKi26kj7zY
lGgywVUw6ITs10BJMfMComQeZt6nYEfBdkMtbZldmj7+SR+BdmUL1R+JFyfRYbm6rSxfSzdkGUwv
depXDKMiFQ1s5VKalBeGzIudKPZ4eA1bfcb2d+pAMQqo3qA9upyOa3MUcm9oXZRuDI0qP5xtjI44
tB/MZhegWOfBq3mk4gdyqlyrHfs7JqsCDxbzF0NjZVo2nY+Rwr6W76ssyUBZhblyPFvZmfE4zBgL
rUdYzv4kURWEM0Fqm2TpF+6xR9nJ86Ctzik55tE4lNhMIpEtYQgIU9TDF7srXJA/p38pzI08WzVW
fa9m3WjyifYVcAadC+qJwf3acBYS2eflbijlg++UYN0g6eDP7QqA7LtDjKNUbZ80uf/GwhhKf26m
lAem6QwgzkQiPsRn8CbTJWJoIE4MZq5J8O2U/q3kjb9Nwv4EoteS0g2kIuDPjM3WsfnS/xqU3fM+
tKQNnLzyfAR+qU2+fmrxgkMA4iw0vU1LAVwPZjYfc3JsE4vI2XTDSaVN0KPKTD5AipcgmsbhNUNp
aLXfJe/Xg0aBHT6rxBsDV8ZHzqvBwYLAoDa/5Rm4YqDZtR2M7+aGj1bT9w3RCLwnUERHttHR75ia
gzTrYehtxXGhn6r+gp5CTvx4aX2OcbofWuIMAVDTFpPuQuvV442uXqG3e3eImxOo27mLA+luWvMe
2NHmkAwKKezrROhXaaWHQgNEA95/E1mMyEd3Tqbtlzc7Ee8Rj9cZC/1LeZEw/WcCAQcx80nv/bYp
tui9FO2Buh3rocMkM6RWlVAsAKyN8WvaBOnCf8gRUgJeSLErEY/PH5Kr+vZ24FuZYUmpT8nN/FdE
wi2tKbV8PxnzErhuqxLOOg51Xqk9z6jo2pN0crQvZbs8tsfhSfm7bvaHJGc1vKqqvUQMKO1zbfqQ
+CzV4z3Wcst35N42U5H3nQbPpRLJwzPb4s38YdOXwnzWTYqGrq7WmdUifA+S6iINa/eNHxNxGjph
F0Rkrdimtjnn0AxFucSntZzPANdCwglzkVAZHf2/rOt0jCDBfx++nEC8gZ7y9hB6WchG6QIqhPx/
P+kZt2TYmPJ0jDw4TOAQw3kh9w2hhs8/sfJfeJCMZsqVDr9iiLysgWPGFLx51L1BVCHwtVRADroC
mSu8ilC/JF53VkVWpFzKVdnH5caSnn5awfrtLfDaAm7zodsBoIbxnG1//Ak135nyOE/4qembBa93
AMyqLdb7yvGAIbTWzZkd5l3b74YEqbHzifhQHz1Nbd9+bN/ABKHji5x3ng9dx4fWKnKFFiA2KVtw
ya0q+7W0HThbDTluvIxfxWaxRDkO6JnEfJ7wrmCMHAMgPVBjMynlXwE6YSM2knWERSdQkuCeL/nL
MWNUu73y6hxl1BwjdWrMjidxUa+ib7EGBASDXxuvJ1mv7qAb12oBou+UdUl4mS6iLNZGq0TGlhCs
kTZAEOhK6Kjd1/dzFYL1TFt7MkA3ejI8mZT6R7CVVr9Rqv84+cKNeGPelN6STKLVTMMNFcDK/935
FFJPD/qK4QREA5o/onYlc1OtaJA/k3DY8YKdGW1lzuJXNQnsMKzb4eCDT6ZdXatJBNHkkW5iq8RJ
VUxCbnD8wPljcipwkoLDN1FtMzYsZ2kS60IohTPgvLvd4QCGdbUbA12O95ejJkxtfCyI8kp0VaOd
3t1n8n7cpWGkpWU8fSDICM5LRoCyruH2YgHZfWtr1yCr6l2RczHY4tDxRUCL1C4EisE8dj5hC5Cl
54s+hUnuGFeElS5jiGQgDLE6opxx6bePK5mXBGLkgC7Nfm/eoXyDjDNXg08V3g7Fz0dvYiFqHPxV
+pnl+sXSGGj8I7oUUnvMzHmCwsj09Mt4aG+Rf9KXAf9UtS8IeMpuOGZviIaxiiDrDWvFNkamFEvQ
3XhfYImN2WMFOqKmRrh9JMxGk6smvLDwfgrGkDuLVEfssVuY5cNr3kn5+15jnNSGn9dZRWJbLiwV
LSItzE9lYU0gDyTFoDm7pIFsLt9kW7QdcW6nVawb/mNO9E067t9SySyErDLrHczz8AhItW8cIhed
VDPrKh8gOrVpPZ/u/BLQ4OPGBK8YzbPMFc3bATKUaPqQfpkWIw5EfltdboBt2oECCbWPda4hBmde
TqKOr4J5ChVOIAj4oIBLOZlSzGtjZsJyuYRF1vDjz/qtO68oYRlh60jfAHHustCDRzKcbgoJz0ga
/XPAlhbRc0+o5s3iJx1+up0KJki6jNRdF2z0XoIqdGa+hAr2Kz6d28FnbWNEaIC+miIhol068I1m
LSS8G7FXfdK07jwNGDYyAvEuhlXByYzA01l9N5JmAV+ivZeb4pGo7S1IZ3a8VW2JIAcxBmnm9P7/
gmkMTUoh0ZnRyEgvWEhLmIcDUKTu/KaGLO1uHtv6x3caFaF2piejgU2aqk9mQnjCteva0EheVPeo
fv8w3nhENmiNwr+EY0DdVhYEqpJi6IZICZ4QgHoUxUCp+2iyfI0YWKhROcKSOUBVrbHDEc2BHY2S
dOQqoG4YgOhgZGzEAkO3zk+5SHYfeW+UDQwqGLjoh4XLIAGKCCDk/x9As4H80F+Yw2tdJwmrhO7c
6Z1vd7SkpZF0wjEXYkh8kVzHrKgyZi6WzzOq+G7UYSYe7IotxX12wbmBd68wBWaFOW5Ea577t0IX
6KwFw3bJmhPfGwie6PjBhbbrpX6fDGAEX0aFhx74SfDVMWneBegndud2T/Ep3Uaw5l95WNoBhMpK
7NC+DbLI29JC/9y8IQ81/Kfb9OkJ2EmwxjpzFbJ0lMyGm9YQp3JjMnoqyaduF2Gx674NDEAYjgJU
k0Ovip6j7/xwbkrFQ3BB4flj7rhMuYGke/GTfqeWU5qE5buBVrQaewPDsc9oktOwPbaHKqKF9k30
hQVmX4S863f6GLIv33fmei3TylGR9Ibo95xoZLcDdRwmJh5GLy3Z4p6GKs9GKw2xAZEoJ5fttrhn
vW60D859aOsfVXvX1jyooYIxCQ9ZKKY47ekZU3525FpFWTGSVApBVS+W4L36/LVx0BOcq9EkyLod
OdUgwRRVi13L1HaxdqPvR8X5Uo54JY8wYiAYAES76EtaxHggDtaNi5SQkQFUSP29HSgwKzhOJ+V9
vqz2H0H2fMJhRJr84o28yRDojtTYzjU8bkgeYrfBnC9Yf1Bfcu2nGnQZTIiOMDyu5DTZsiffCJSh
zDShXpAOFGnqF0+UcrGNAmD39b14lHaxj3sxHT6uD16VzRtNyjEnsDWSoi5z4yFjYVk44n9dYzhT
A0f4Iw1cgf4O+VrVCTXo2A6VOCVdQK+Z9uEnnMj2vLe1ZwCbk8xm8vEsG9Zpt+ayW/0km5sshcYo
lwBdJeg6Eo0BadDreduBQTwo/gsRHC7LDeU9fWloBY/WnRyoEW46BSh3X/KvpH0huC53jzYAPYW4
5wE0ovqbwk0lRQmc7sy6IaZ5jaXl4NxpoMA6p3mUu/zAZj7juKTmBU44dmE/ZWHQYKMYzJf0KF94
JllE9Iby39vaLGBZA1gWvLhJgdOvoVCF7csu4cAjMTTHCfxYTCiI4jFuyz2th43nAkmaLZUT8Gmo
gjr/0Efk1ZkYSpdrzKkcLqYa1o5MiiiMhLiYG/vJtp9ZflyKfPTroeE/feuteOGq6svVrNkbaf7Q
xFWHFKAm3EwhFclQM2Z6JhI9tE7YTki4M3WW8J4WdxTdG0lTkZZqoqjqpAzg+wtfLCZIwjxTj9Wp
fPteMxqBT43PdRt8nOAyi6jdB2c2uqIm1itvujLYfaIntnVgwRYapUjiMcgZRRKUhWbT3I/t38U9
/Hk9EwJJBEuK0tTFT5lrwPqTfS6huHjJRM8c6G4hZYS5P8R7aV74SukqW20OnDS0Ho0MH+y2liD5
aZzNhoVXJNNt0sbDvEKkHuQju0ZU/vvbZlJIlVzvZYtaWWLjlZTh41EAmYwwJ+6gEwMnfUlaBmCO
KONQUEON392CeKJJciSbfVruwEwS7h/YQNWO52P/MZAw9IKxztIwrfFMNGd7uKDJmLZbyO0PRk50
mBQdCpaOjJ0j4clClYt5mdBFCK2NpKdrlWngt2kTSWOJGqcjkX1i79FxOxcirMcQNZwEZy3ijLYV
vFpADoh/SmEVXiU+kLT4ADxGzSv8OdA/LM5JExZzyCkFTNixJnNUx1SrnHcQ4t06iCJXUi9Iebkx
nS74a67nW4HfGGY6fRee9qn5DbzonyTBOO8Vugrtm8kFDzT77W6JIssPogadMsgB25xA6BSqZQn2
qIkFApx2oheeG2ygUUAy2IHFPxtbYRyXyHTqQ7XJAPl6/eV3onIhk0zfkP4frA5YDJVXMBJ/Q0Po
5DT0I6S6bnkkOE4wUBlYu0dRWftqqIbJsCJO0Utn+/dFGrIr3TMEjlks6rf5/+o3hgkYHqnHIpMN
oqBUSGKYELEfI7Nn16B0qVtDEGBaSOqN84XNLojYqVD3EapZdCJhhbvPN0O1tzy6z1JqQwuI+0/c
zyxLx0+ahKdrbQyaKL71VmLyhcINpbmhF9GClifYt+0NlMAv6uKok0XO0JknLyK46p765/jTQrXn
NdrejLnYeowmgaE9AgN0ucX/Qs7LLwo2ryi5NNJFPS3xd3aXbSTR6jUkKwgYjyC9atB7KSdKFSwY
8JIpWjEyWo9052rlbWsSm+QUFbJvxBKdNrapM5w8T13QNR2fy7ZIdLnwsdcoyvNHimt7ANuc+I9F
PSYX9lHJQNDs//e50g9QEuXMG4Ky8MGtfhjZQSCgjbRYENicT4prQNyBGyNCRHIB5XedlerDfUsJ
2oydUBx8+hClOV5G2UUAsaXVqEE925dDss5dYBDYUoAvHHVz8eEAXkz3OUiOo8HSxSqvv8vGOPrn
/44BBDZ8hQY0UhpZO5TbvhCj2U1ll2VIhBvtmoW2hlDaEVx2mQ53y2xwHL9ZSZgnIbF99tGkUSRo
IetfcM3Trff7W1DbAhnQgFFrfMi/rLSITS60xGfsTif90Ptm70m13qMUzFeulMwcC6kODlZb9uST
rog+yJwftSjbfV/Pw0XLMAIzMo45DH/f/jiXdIdiUG8HjArK2qEeuUNEfvqn4B0G3rYCm3xWnlDn
//Zib1YceMrEMJ+Nf/DILID1cS21aSRpjzFN+ZZ6vkaa88cnZuxzCV71bRLBFeF2DIacg6t+XD0b
PaeI0ZJzPSMNw/4q4ScI4WffZFt+Q7sEzrchHBf2PcYflXHpbdreac/sKt5VKADO7SSSdTpxDSqZ
g6wFwSEq2INdanDJ6gqCNJqX7A4RSqBsr6MpTJO+La1XchVSvK3SPF0xnZH5D3/o2XdyHMMiVmCb
nn2ZS3X/51HosCkNpTT6d3Vzi1+ZDEELkMSvbk+OxnYdRXZ7baZ/tVxWOpU0Nd76iqs8FKUEOhqi
yqG2PUlGiMXP4QFBURZElVOmLF3Vo6N0figYigZ3PwTb7O4zvIgVaPDXyAQDeT1DOYqDD5mi+AuG
eymupMZ6KqpL6tVvN8lIvEbuEX2/7nrv9XRGZGS8EPfgDRXpgfRGOzS3jjbUikyL7HRnTVjHDETR
IBsWUUgi84LyZHXWU7007/Kvh1QvvWfH1SxeLvxb0yi0tqdbtJboJVjqDD6wyE7/Ci1GwaWuhxrJ
+N+FLPt8dLOXnk1XsKhYQS4DucdEi9Ru52+z7VyopygvgUyPSNhcdB5kKGZKUdLx6QtxVyoJQ3HH
OMqzyPk2TK6e+o+AJSl4G/24aw17zAv1XT/d5VtsAvwDLbBRmAMCU83Zdx9eeTiK3eSGdXItk7Bj
xy1tojZnqxhvAbuvYysVJKWBM5AmrEyZyF0P5YP6wINYJDQYvnygWn3Xvep+EQ7xeDUDwwEjA1fL
5HvFIBXSOz4DzMOgND14tiHndUTMiK1wlRgZ3G47v5xN6G9XVe47KhaylpNE1GeMncQQHyxKdYtn
y461bwgP+xPhBwlIEW52WITWf1mVQni7wBQMboNU+dbVAqUMrwxtdOkjDjJ846SI5/5L9O2Z1RD4
RecGXfZhD6zM5gMuLH1VcVSI8YF7gAtdrY39XUrOwt2ZDqDQPAyo30zseb05XhntiB099xt9XCSL
e2/FGy9ZEq1cyKumT/KYrDlx4lRnGiwf3HMCX0yvxsAYsjLw1RjhJPOOq84d5mfZam/9EqLosvbb
s1Hb5JmheImwG2Cj7r5kJzsyRmYMWJiVfd7vHA0TVwWqQI/Gvl7lJUSpUF7YvgwxscSStNOxPXDF
vIMLCxVZM2ivIBJ8sUW3PcB/rb9WgPDmHo5m/NHseSo65OiE6kl0VJblJd8jOO/fxUWsM6o5xGka
lubcmPAhvxupFSQA/f8dBKpi4YandnJ62o/DZCMVrkal/j2HKvEFojavIBOON8gfVrMksprUr+Ov
pO+qzeM2CBjiD+7gLPsD7Sn+UM+axDh9R5U66pKO/Go0VtpQkJhTaQTeHg8g4rOZahK+Pi1JWf/Q
Z3dQbONm25GtA1rRh9x2nLz5XffHFb2Twb3ixb9AENIdg55B7om3095ooe3ORAXdZ8xA49d1PBEZ
BRKepG3k5JnjkGAwL1vpb1lGnU+OkYd/oH1akY7V4vfK+Dk00dfIxPyCa/LHEEnwd3+jEYbRDlQs
77dghOgiB+49+UlhchxhH5MnhNJteTwOc05cTawKLBGbuLzzhW1rXwMr2qInlWOvU3cuevLd04LA
q6S+x1KPxUEg5/I4boDtk0r9j0cMGKfXMKoJ/pBGNNvNHqB4stfhxIiBjnnE5MMksb6Bb2/R6qVN
KJfuMlXacL196T+T9/Q2ZJN4gK0AvSWDJuLmVEPRPWL07N4/oOlFicPYKgf2iqR5XDQ/vlJkI4Ux
vDOK9R6jlc1CX6oDqcEUZGyV26ys8nLi+JCvdwWQBmmtM2p0ic8GdVauify9YyEsus+smRXCLy42
kdCbovCohuBtnrqQJlup1icOYMklW6yj6p6+7I1LfVlaPLWasFpi7YFvnbAT/a8YTfA1xyxmv6yT
YW38nqfevvjJS6B6T2/Kg+o5yhrVXAGQY+NcFjBpvHGeomAkRvg4Z5a+j1/pt2cuyXTqMP6KFJgq
8bNMXlxd7gGjQxUrOSW6rn7+nW819F+InFl4eB4Dr+aJ7+tsqu69sguQRbbiTv1EMomRxoX+LLPA
rU1DHnZDAXrO1gEdpWZGENJh5h0nC3xU2/fvQVn/r8r3WO9fGJuvxDFCELhkJFc1QsMs2wn6mfJn
XjC+Fsytyr/Ywz9Bfq6xXPiQ1noohZhoE7tv3YRni1qhw4QYp7DpiUzJcfF9GuqLuMIC/zDQMo8K
2QCOST8J1mbJrl6VdcG69qp9rUFBNeN73L0e77yqqdHuQYz0B5+m0ysVjTD6MwXdgkE9iuua+yBa
PKbL6x0PEL5KJfDevRfB6nmI6xbLRotXaYxNMICHp5wLT7Iw2KaSFLzepVVN8XsCp0r2EW5+lPOh
ovmaVzRs8+DXshSfsSHt+TWlAOBw6K8/gg6xoSc2D/M4+WGn+FU4hSCsKOZIF/jTN9s4HLCgTw8w
UFTMqZfZ303DrO4c2qjfqYVAf2/2eQcjwjR68wfpQSBgZR4Jpslk3/sNj6giSEyAffaVSuPGyns7
v4jIpAb+0YBbB2iqUggTJQ3Fwwp3SfVhKdcFPPORuT+X3nwI9Y415uRlcyn8WrhQWY7aY+1bQTmR
F5G9KKW/3vTrT9MnHmkNFDZwnMOMyMH1+G+PWBKnEXs7AuVbJbQG177VPZjGP3t4dqV/Yrbv6e4q
cOCm6M0zpOMzC75/gqct/lDcg8fQ6icqYKvc35aEfyd0r4sZ1BF3aNVVsUZ2u/iVD+7YISFygwAT
N+sqj5ps4fRXfp3aoXzPQuIg7UhbWp9k0YHiRqKecLWPsMEcjgOJFuv2eyB/JJEXX2AddtwbLJgi
GR9x98wsGaaeLyd4JQH3WBC9w+EPL4lyca8cpR8LPgWkrCs8IpIElSLqECxNYH1mLsH9x9K0y0be
C9NO3yuaKSGHxCay3GS/dB7vs3NMv9wDFijngdDhR4mgbyG6e7Fdby9WZmDKAbi2ja+6EN4sXkPR
dS/GIlre1IQ7JI9lZBvKe56Wx31ZhfIQweijY225BFXsHJQju94BNWpwz1Qo/ydjyMAgfah0NqXV
bv+aICY6FJvSWe0JLaISLWFn9sioXkFSla35N6fi9Mp+8JXzOVZBYqMe82XghAPcSxvt2ND3jyJI
C80sw/ye++Q7zF5K7b9sA5ssDyhDvAWG2Zt96F4UxjZICys1cFZFzPkXIAoDSZX+9j8ywoY6tueM
eGMs/E9MNs6r0HUX8HM6TkhA6lvMsvPaf3ff5NSplPKcFZnYAorzi4meL/VhHa30te5eS5g0zZh6
8GH4X0Xhfb71UqBqpmUWyKqbfusMNhjwkXr+x3dZlYr5HJBSWSsEouQ2DrsgDg5kb6ED0dCLlxcQ
7mmMsbOQym06csceZ0bpkbBdbickzV9iAto2Rr/9ZzQtNRr/4+2UDzmnNVAG6bTXe3JCIGxF7jG4
I/kfrv15YYN2wn6IX38INgpk3tsb58UcI8YJJ3FwcxTeBNqxQNAqxLT0jq3sSAUThFQhNjJZlfLp
d/vDJiUst2xdA20uCAU4uvBxrfkwDvWAHCUb8DNdNENJ3RNphWyk4itLK1RFh6/IN9luPv5heegE
DBkBSuCh4k9CyWZZsc2UwAK+6IgajXB5FA5RH62gMF6J2qMwsFX6xmZV0hpVmECYJwzO3a/FZoJs
TNECGHKUPFEbyd2btu8aEvb2wAaCa7HmPMlKgzDOFv8ujNNJrD2l5Aq25WBtiKPjp7L7pjX6xzQ8
oWcoU8WKRn4S1VFdErE9m1IPc5vBHmJAvtYdxbm45Uo96fREUiK0piUK0jT6Why+W2w1QxwIETLt
68cHjBTMtXJ5V1D1x21FjfdCGF5b0SnBaU10+cs/EzjGcnyWQ7+8KI2zhJCbqboQ6RuvHbjLEFiJ
6bETJreyYqLcN6sa27u8p5QEdw+Iohpj3/c98gxR1Mnu8xKTxWvlUG0gOcY/rGY+paM7MQIBwL2G
DS0QJkB/yf5LcNO0i3EtsG/N5T1q68GB08jo1hDwCkg7vIGSa3WlhsbaQevrSTOOmPE6oCY2QjjV
+kBolZ7ZxZ9c1jIJ1DWPgygo3qRI7txC/YTYi5UDPCDOS7xtV6LLBjED2drDMRVOclsha4viIVcn
49sfBWA7efwIM6WrN3XZ+ofb4DsCq6a4cdQ6FXxYIeubuxGNzT/J8nlAo6eoycr7poVW23i7P06h
2Km1ZJ8tmyP6S/Hz/8gL2ZGruoEzAnmhF9/9P7cfZMM28iciWQ6KAclQTkRjUxu6UbCVpaRMyxas
ayTfmKrKn/CPdohbQ8jVP/NLftPLkFUQDoISVoiLNx9D8xM+3kQGLEV5xkxlYN16dYTpLUVCScMX
JZHC1dhONI2SSX7yFAWjivDa6rUtpNyJ1G1425XBvwscKIZ4EZcmWcC0i06D1ZcDKT2q97AGHLrW
6cB8eOpourcaBs3u62IyKaxQAyxfL1EZXYC6xWuqKw29h27jHzXMlHc/aa0MaD04OW6O6hG47+p9
5NUKb7i9x9lOggNr8NynGD9b7E0KGfTFzplh2wjcNksr7NnMHuWxFd0vVO2iXIcXWhBbydShrhXg
EghOj8qSsTJYw6QsWZhIL8Gd8BDhPZaTldmTqB1LyygHlcxIdsiHCyHPOMh10GKQOBVg4Tbk6T+l
aeU/7ycHQ00WtNS/BkrCs2ErO93HkLvHqktuQy3+JpeoLbD1ecH98oJeCijQ5j8wXFt55ml+UpGo
DJHpsBe01fQaF/ogr5+d2xstJQ6we0qqrmXrm0zHcU6Dpz2jMmRqUjNJ/oB9YCcDtUvocsC6ESdp
oSrgWwtWl//748XQvHUWvRzT79Hipa9jfw0UVch8IrV+9BY6ADT4Rb0OTs3PyXVmv3pKlE2tcd4n
A1jU7g5WPPilb+kvNN0Ub5rgvEe3xIqvkFp8m+fQeX0vU/sVt1Cfx2ICMX7mbhxMhnnt5weXM7jx
re+xaZqTr61JH6JtiyEj1ZNzeV2+hDGf+96UKcSLRTXk0OlJwosQb6M2LnXAbI+t6pFm3/EVyxTJ
YCAbiKOyMng66V1iqP8ihJa572Dg6GTnt413jrV+vEh0GJnPanW7SNqG2b1zqKk2aSLKKS/DXGFG
o/Q/HNYOjYeNaFstToxGTLQ2o/lXQjYtPFSz8+uThjLu7rnNeXIAwRzt+DtNkizPOc9TCoUUpBCL
x5GiIvEOaOnD4MBsF7jSrm5bqgys6FAR76Od8neP8aEiYh1ARsX21OSwsFc1y+0ro2Njlrzh/g7A
j48zA14m2n47xFOyGlQW8WkGpVMJvRZathv5zqVSG2J382pedRwSPsfsAl8tmkl6tOPDkfYmUXq2
+6UhmSMO+zY99UJUFFnb7XgbZpjfnRgSA+R5l+3emXJDwv+pzxRZByalY1nNbm0H92x8NznXObDa
WJUyQwhog9AW3VZCpAtytdJQlOaZudWFE5m+5ggZIDlNA0Kx6Bd5MOm5WOCziTd2Xy7xkTo1L4pj
7NDj4Wdnqr1FGMVv7H0J5ugosQVubTnrfjCwi5KM6bkQRrAl0nGmgumwAv+oru4pg+mkdrK4DB14
lICIQi6FBG1x/YFn0jS95uAH9EOx8/6c/BQeAmLI3QkNAMSEQyRQ7uKSMVuiZXjbVHLt/JupkdSJ
0hD40ecvpgVwuBC8iihPcwMOQ4irOUDtHNNVri/ROwu5f15+TjMoAp/7iiVgqFnLRCl7pOE94eUi
8HViEhsTvluV27VIKJcBJxfUWrGpLmyAXlgGPwwkojLl7ERF7E6H+9nWf0VGsXHEy3Bn7aT5MOOt
nL57/heI6EHqNEGWVSGUZrTjHPkrTTkOPFFhFSdhxdKN9+0jChabzUJ/FW4U26iOXySUnxOqs2me
c7LiSqebrUCBxDkiMQVW4SCYKTbtDSr40z4RxUU3QZf9FqZWy9O7GXHwjcLOUWv9ZZAWNLVRidaG
eAtJfzL3XXbtCcG8/j1aDUbuc2K8O1wsqCdFEbUODG5Mh/ZM8sTFG9przaTXzLILIM6O2k4/jPq6
A20eh/94znFJDXzUpzoZSu/eduP5pinddfifJKVHmouq4FKOodFzVFSH2I9pYjL+HI9Wp+d4uZTa
rapleZ8aNFKcYJevfaZnXubSPLm+xD++y1iQKuhmq3WmtUGgV93RXXLVX04W6Fh/SQfFt1Ud2JOH
45vo8cz/4jpQAG3zB+oEcmjIra97/9+ylTAuErYdLc+Us+wV25a79TljBNB9buXOAKnLaOBrtjUG
Nd+q/hsTq/l4eC5/n0t+3TIw8a3/gDNWozUzsHN3bQ+3I2NFY7LYbDx0FkxxPCOMsehuglAkDJ6c
W3SC/pI1kqgCxb2/FqzH7Yai3SRnwBtHv6QbnXQ0524KdBrVf4BrHny1uekG3x+4D+prjYFdhRze
rrYIj1wKWiavuMnpnb8woYSygNu0oFQVolH6rY2Ap4IQ/SWcq6uKQLv/h07sS00EKRLo08Lzn20q
tG0OBYrifjf00yjuQ3l/jsGixLRnF69VXNY6lUWTiht8Z9BIlxNfnBYeM/lgu7QC8Mi9TVO5U63a
YNISql+ThnJvQCqB3YHcYTeuOU8vQjYfmBWzw9hTE1WN8sqJHmyN0je6I4vdUymHVw4w4JAxJSeS
q86wvTGuMfv94ZFD2GlvW29lTkIT/XNAW+pBVs0Qgho8AlJ4R1hyg6MbtLbbgUxv1iuV4vo5EEDz
evizr0JOcw/UjlF31cITx9Z/W/iWVZo8nyJdU1UU89x0q2r3eg2oNTvAdHtCKaIfMIxh469UKu4+
Y2rHWTWnBcKPewGEipt8a2zxjbJJNguru1eYTJuI5lanO03Wc9Wc38cDxlYK66WGKiZ3WYPfcRcq
vII+it/I/7EpNNkHCA7415t2QZ5IXBArxXVkwX7LgT5e51UYg0QQTUu+5Fw76CPtQuXv0z02CYyU
kQ6BggQGL/VE2Ru3aWl3X4vk/8w74WVuTucJfIwUxuQf0ZmWhrbruaG2mdnzWph87LfbYYOYCKZk
KQcmAACXUrbsNFQsWHBHK8hH/FAM9aZemmsdCIfxqQolhq9Yn/vaWuECoBVUqkcVolxquAHLFoPB
NKqmhlENYnLoQktIhriJ7KA1Fj8y5JSg8FFfhB0x9yKr+Hkj766E+zwQvwfJq+WHqQEjEqeiiutf
e5CF+uKVwcAO4grIIp2DO97jaCULBlAlbdvl9NhNDOiyg3e6vTTYsGwSZmd3qvNKa6TKZyNdasJi
K0je7P7NS4WgFKg+50d9ESDcCNZYxrmWJkatn2X0OTWWZpYBRFhs4NvdAdeln5AU8m42SaRTpUGX
li9pGcyjt8lfl/XamJU/OxuJ87K5/n4zn8FdOI2JtfU6T+GnBSjHnTCh1uHMAfuWLFNh0smeKRoi
EUJ2PqfgneKLWQIgjPC3jxzDSiR6ArMS/8wxoWE9LfCJnXhlm31oy17KPw7/Otnq+i0Iw6m2z7Q8
L6vp2Ki8ww+3hGI2l47xvNGY5mvVobyZLoaUHlngqn/N8M5q6HhVCqY1fae2L1RdatespSmFhUqD
tQpNBI8f2pghGI7hYVfFUqtKa6B2iMnymzf+8CmLElsPCEU9pIAvnNai0mKpZjovz69GLR2q2Mi3
/lL22O21yfS/kv/FiH+5LPoc2pJmmfb9/DRMOSk6p92eCLxd9gq6ArdqXOH2+PmgRmggb/mCT2wP
lnrWdMz5ADawiBxba4La4ElI4VGKepLyeGI9/i8SXt5Yk9D0gPN0zghWzgr5SnI6e1MTCGVs7zRh
nrOT74+dw4MITi5aXNbGYVNiQxXld5xKFfx9mjPQAH/+2w6kKMZWqFc+UGPeWQ+FtYp65KX6tCvv
fpqy9m+hc1YKeOL8S5ZqBbZGqPrGd7CjiXsaOvlSOwpygGberlCW+N4YbTnvIUGYvUe1Y17Z9TTS
cborXU9WOiC3pD7OGW+JxYpJV9Gmy0Yxwhed+J5n8XiIRESjB8wjAnQM+3n7wHdiFco179z6EyTh
bo4UUFV9g317FvmoWyZY6VAIp+5upypTx/gZfwPlc/5bBuVW5qfRvdvT9OoskySHIEUTL5qk4mTI
hDGhkrINWNIe1v6cO51IzvWDCU+EEUzADi1D6LlbhMK5FWyWWDisZTVKq1THAwIDcRJZ26uRiyel
wqmmeiKqOxGrxSzrdcuCsecnb1E3EVmtfXB5we9lkMq09emgO5RzWzIe+6Wwx8uWrWtqsuGg9GHq
A0v3dHoO5Z7NIF0IPPhfL9JIkM9cvGKLq/44UHbKP1J7P5k4ra0WW6GHXP1rVuTT9DOCnYqqUS1j
VrFSNHEQ+Y1kINbKgyLSx3b6bAGol5zfW+NTFRDIMoRGa0S6eFPfHf3keCcfd5N6K8XMhKFgdli3
IKE5hq7De5CXv6l9NYgQIb1UWJ+ce0ShXiXoFKcbNr9tyWnGY3GFElOmMBbl/FiUz4eAeYeFfIT1
wM1WL8YoI2bxAyG0HPI/KNI04+mN4eKmhHzNXxfMNrHqJTUtSySeHLwbRJOF/ZjlFDb1WZCUTjpk
B+6z5f7l7qbvLxJoyPsrhn0bADcTNlhxvQvWCvyQgLIGARYNHx4pid4VFRFl4W3d59lKKDU1O/BX
ITyl1dhme1BPa1kWvHNSnWEZMTHxK+t7Yra4E/9PHKXlRcBClnaFRy14+t1ku3eklvge9ygDxSiQ
dINkrWb8JS6Ky14owc/QAj6jW/+a/zOuyrszVrsyDJ3uJ5TiZkh+nYMQQm+y4rbuOu1Tp0/nFsAo
CPC9jp+IhGsSWoLa/B6YThELIQHICTXjghZqKDCJuPMntQ44gALi/kLceSd03p49APtFvJY/p/Cx
1dGpvOposd8EpIy+S7AQ/oaaBj3zgDf4520aScGwwOnZBCHcv9gzlYZc1ll17hXzx20jwbwioo3c
dEChgVJya/ZW/Vtcy4Hdk4z4PYjwj5fUbKQIE7ZzAhEFN7dLG/YLBjMgSBiF/eG+yqRXupSexp9T
goimxXSS998vZwN++z8ptQX6zk1XanVPMlD6R2C9M8KRPYGyzFvuDAeWonCjgAevufbdwYnLYBQ5
nI85geasTfoZJDRsmCU2lSR9+SI6wdAz0qyxlSfkqZ+yeguC6waLHfXZzZUyZPu8iNt3qvcnAHk0
QGQJF6zHwj0FR3DeLBKsS5N3yacJApnViFk9p+c2wjjRvCxyVpXBF/Ok9lwcNBFmkvyZ58iNuW48
LTghIq/RBWGcEdC/L5E0B8OG53yYecIdykzUrBlaxcFVFnZ/YtL8W0uDKQLyV3Un8kzdQKlkp2BE
vGK5hxaQx9gO/iMOqRQ/k0Zb1vTvAX86OXgXanOaA/YMl2ox9Tu4PLPuvRMPjPkgOOIGBMuNm6W8
ZV70gX0CyXi0Q29xTqRdSjBmikRsY9SI7Zv2QKkrA14GCfrwcYWzxr6Lx2ObKy8M6S5brNSteF+j
3hpbz8qhulSaB7Y6vCg0ys0bCQo11xM++a4yjiU8RT1pC4zkw6IK8MoiYGCv3njIRTMWBujpjTVz
fhQ2h32b4aKVtinlg176/fBddbir7en8VnQH4vY82RYpKPVHg4rQIGthJtWxif8HDN9bMKEDUTZ4
IKHAH7Rkwu0WF38kgVxiIjZioyLDP7Co0js8jOE1noBHvk6031GmJGB0u9SGd+q8GbXDcNj3MFrC
8GYarAWVVneixrfSWo0Dea9kb1vbxvslWU7eQfN4LpC8PVoo730uuMOvQQqkV+nRnSa2WxsQZCkU
YQh5vTjnY44OXvAFcdJnY6SZmim/Lc7OiJ+R3M08+lu4irIPRUscEJGyZbWLuktMwpwG1g3GCAxj
dtuLGKO2L/T8OpTakTNZ1u7c3SMWgOLEL6CXW9lra436/WvqGPdgAU/E+7PAr0vPxjbG9D/nFo9B
Dnpa9L6cWbHdyY93CfG9ZLMY8IlP86Tr1RpFIcKNsCW3MLpEl9NfrtDjqlYmCKC9FX2vWnCIDZtO
OQ8du72xikjFKpLKQ/8I3n8GN8r2AcqtE6ezUuw5BKnYoqOT0WwhTxndYsynXzfqK18XPv/KkMnc
rXuHYTFGCSeHwD6sOgzDswsSak3XBWxL+rtj6tPxh3puh9t18ayhztlATlJGcCvgS5wvpn5JZ02s
k659a+Pegc+wq0VsGRZd5vRj0ddHcyOgLAmHY+UJsl2VvoSPb4p01mRouUBFOJCx1He3/FTHQ6Up
QfpuehsHsJymTMal3ywkQizlHZbfkgy95LHKJwYDqrsbdqlALbhAL4kLnnPe3S8UMETPr4em+Rf/
a0T+Y1vv4wHvE+hkgy2BdzPpX4YpEPabhluz79cGNXD4nTPnsMVXFFyTbOCjWmSNCmricQyoNAsr
X2AS13LyxOxxWWgy+9/Zwx85aqsl2kmkh1n/5Di8UBo9ouixROlYpj3+iyxvMz2rg056p0eo+IrO
lZ/wppmAlY7N6iOVV7RKoTfejbDX67Aee+lrOq0+k//Mfa/zI63mJd8aIxd0khQeJXLZyocgvC4M
wrDR1BluhRAF19/7291WjlYUlmblVKo/L4IPM3Xpo2PMOGZoTz7xVWf8dWC24PrIDm7LuxxeFGMp
h7NgUJM7Twhzvdoh0PNYZjL3qa1vvumvQr5bcf3Zq4ZUY08E5A1+/i+OIB4HPP+QpOuQwpsaShYu
NkM2nPxfDcHtZHrq/YlLoHrTKmwksBg8it9T72B5ns2BNkC4PQsSzFUB80h6sK4bXTCfYI+rK6jn
mnsAS3zHTv1zIGG83fmOqt68xVrDXt2CX/2+ZKvbOBApfJ6n/9TS4StNjFEyj57imksIhuFewxwK
lMK3AztNh3azHyupuCWYlSc3P+6pPnKKVmxYQMrtAIneeXtATrQn9TVnlaycg/YHTLMeBd2tgN2R
BQ5HBtn6buaPl3j+Owdi+lOyt/NekW6OjhWYiso1RR2nPREY5/ODS22cIDbNmbR+MN/m8QZiRAVx
vhOaYQrnkxSGwR+Tw1L1pPK/TKHRGZqVvDoIw5A7Uub/pTpMHjC4gb12Cgv7/Pm780tf+DK/Y0XQ
ygbGrplPECUrjMc1lW8dNCS+LU2o63n3GwuXTIbZhfewRmifAYJE63jLjL/qfp8fDxOsPWxcz6Bk
kzQ/KFvrH/4kov99hGLdRb1WgXC2gOYMGjoMYk8hhr+jO/kz/FqTc6QRobjqjqxuRIqJlJk+EZ/f
/oW5ZNATy57ARXxH4HCkeLuWLm218vzFwVWse2rnsNTWrHOer68qGtJ2LBjjCemo2vhVRd2vWe6J
59Yp7jg5k9Cquuq96e2YDTdY2owplGRQ02yrqET1YRbi7nB4HNwURsShc6JUqxPol+8JUO1mgcS4
Fe9UY7uLkGzswxJQ+CsbyuXMaPiFvan7QdJ1Z3M5mkeULQEroiv322aXu0O4Vi7+0R+QPiaM3TqA
8VOl7iiTuALOTimb4+Msts+0RB5HpbzIGBE2ofrQ4jpLrUTFph7VekZElvb1wwUEQfPI4Cdr5ZEO
fRetWPYsz46LuWLtxsaxMdz0s63JBzulzwr7TAQR2F7NnbYfUanL7NU1OX/VxLU+590RkzU1BPjj
28hLSAh+LowyAE6IAyaDLazk+YJ0IhGSM1z2YSKLh3oKeLlHk4XnUpnZ769lkvYBpmENLc1K5poi
Tbifv9aIyTiAkuBepW9IVLgvP88V3PsbCuNalxmEJI5kyJqneUU+7cR/0RpllMq2uC8IPYMuLP49
i5wraDiD8TH6mwTDJPPo/fpNCbirUUON/bN6E6pwxY1WKZc2zeBUgDZeNIZiVsXf7QtJql7nO0py
CycWCBmwrVyW8j/xzlwYZRSsvTjiSL36sxnwRfrZ6GAsY2v9RwBz9F+zNPGrNkQc9yjV0NpE1of3
olXuKkg47+cs423ok8BQITupAke3qiyAdlkh7krvghqhMI+QhU+2/fmGd8D5pKQOJgU3X0qlkTxl
X4CVPtLE0UOhBA5RAc6qn9fqWFk71PjEfAeDZY0je7pYEnVPe8nqlj21gw0AlRyQf9MQF6NaRgTV
8JRMq0IiIWKQss/BTIPezDL7MUYSKPFDMddO1on7vR5EuvIBEpWl4H6c1iPZql5dR89YN49qQdRq
EjqknU71j+e6kpn3B8ZO2HhRxScXj//Ua4E8cAOVdnjF5jBQKeAKQfvPqE0mBguCq8Eb3yrWCqh1
2aZV1VXjtg+KU5l+OgXrKJfpCcXz1l3ZEx02YsWJxjMHtF1lnzcglwGPycdwmJ/6Qu34Ey3elCjQ
Ff76dnhi4pm8GVOw++ZgXmF9aUnryktyXi68Qz9wV1orCcoBVOAumInO0sQ6rkphW6/TPSuLljdG
EhX7syKVtrhZh+z2Ir9GV1kmuSppyQUvSYZUqHZnSV5mEdPqCPWtmPVVvTpiQXPLpw1NcrHQvueR
riNjRevLhhk6ei/biAzXR0UZlFqmZhEFlLsjK5UATzzjojK2zFU0MGBKl6r+0kzSvhSk9DkVtUOu
r0pYSv+2iweSj6rKAX8FAWo/VZ91/cR2XXjDD1C/zulPjkRNglBCLplT5tVcT7md7fSpAGw6DaV9
1q44ouaiYNyAwzSWDWkC8hnCEwXv5n0uAiCYAx3dq0Ma22kUf1YBrFDJuPrgUu9+krJjQ2+BNh9R
Wpf1rEoQpV3JZLy8wepIDK+sUROLbAR1+6/XGcX4UxymlzGYRFfMk724dA/+bk8GmE2+rcnleaqd
aP/v35ADvyQsn3U+b8ZGLaZjZqg+DJykqc+m0mfK9QeKv+8RSoGNFbB7klRCo7Klpk6/zPy+S5hl
1aJCQkje/ueub9oe/3wk7Q92eIo7yJZ12zC9GIUQnUGdJlX+vhWjj5LtIljieiRdSlc4Aohdf9t7
r0vbbY8rrU7onV7hvtMnHaqW1OsnEK6ADC91MisJiLx5UYml7VoKgfOMMNQLxkfqOg94ldus6eDB
8rDdwjM3WnQtK4WxGs1WHq0YyEl7tnB3fkjWNv1r0+qc4q5b2ElBCOIPEXLk6TB0+134SMAqDfq7
ziXzNoYTLMWwdrL5rYLTr8j7xaysVOhl2JOIlXDVZ/2Rea60AEMTZrjIZHDtx9mMlSmxGPC9k4G/
sOE7736ucrxnyJer38FQUmKcNfQQpn9kPI6S7Z4X/FVXfwgMgqlD5ZsPMF4YsLN+u0l/0UZUTMvu
CCPFE2tzpWd9zNPFWtEg/nSTmWGVY0D7w9x1anfRAzgE54Lq/9CwzsWT4WQ4I6zh1/lktc+ym0+4
iq1LUGyn3M2cbwszgHj+WXIGFeCLdmXfgUpEGoWfTQDzyy5uN1cFrBSSOsXPdyVzNw4Xln+kiSJN
3/sChUa1PFrE9gCMVoUC0oXGWvJEdM8ZGITd+FHmodrZ2yHN1fa1PT6OUolQv37ktCRtL0+AAqbs
Oe4WaUra4AnEEGk41StMVwJ4eHBr6QOQ1eK+KyLCLqGFsCMZTwF9U/I8UUPSx7/ZUpBD8JbQXpi2
TemqxqplvKsUFMvbm/C8Gwq34178ry8kNj41N7ML1k5FhMB0FTOE4vex8LfvoWpj9zVDFWuwTQAj
McXFV9Uu1kpZpToNfM2A3LpGCjsBEa2XhQaELzByhoWzrukv5sASZyKK7G/5l8ZiStWzZFglta88
d2pN4XSpDiHfdt3wnFvLv7rXmHONIA9H15km7eIbQ1eK7DdSoZbahbCeUeh8IbSmE6CAP2W0j90U
BTjWcMHHoWJ62LDAuROP6PFhnJWbTd/NWStFjD4TEqlZ/2XzLYFhPQFgO5r97mPXSqm8YnqemJlk
dERI9tkn3u0HhVon4rudr0+U37nfMby6BUTj2Z1/XLgd3Gph1hJSZS9IMHNTi3hT/1vFLr0wGjW+
NTO+xFY2xiXXraeTTHlvMTIoghS0VqYO9Yw+P8qPV2tls+SfOVyEU/qFaNb6XiQsh+wtsBnidEZT
V9YzPp+JKJPUaTkBfgWCJXwaR02qUlt5EObrDGR8j1Rl0RrkOxEIiL02+7NJ+vHy2DM9Q/32tVFu
hcFMm+073+93oDvB5PXjfVdUkWjKpPQ6Bsk1yOywIp5Msd3v2LAYSW6nWj60iuJEYieyIowB/Juk
RcYsjgTR2iGXCCkqkNZKwJepomEP9rqqkdYUZZu2MyBvltkbW9zYP+Fu7QX9MAHFbroSC1GjpHYW
fPvi3I6uJvZRADoZLAt2D4XtA1me2tgLqWi8/WHE5rmY/vC/JTloJ+mV171nI2Gba8gq1ReM3AgC
oVjsKMvGToQLYkR3Wbx4XvvQAfCS97WGHZHCgBVi4MovqoNraxFcPEkOCcb9XhT7liPK1vVawpSb
baPfDZBdTREAi66GPzjFgRf1V2RczFILgMv9xqxZHPaSKKrsvv4aWmEEIV97cggd4tvnmuYYA/F3
PhGm3Lf3gTcoZielQoosLn5RMDvMij+C1sHYefbeXqFx+5Tw6qOsir3qtHXYuTbov7GbUoln3Z7h
gwf9imhJrGIobQWp+87EGoYEQDIJXbssLwgh6LkT3jtIubHjeY2yTZb/vUnWZx+KaHGb1mGRQuUq
KT0oHFfLPITlu3ehBeFbLnh5CkK8V2gVz5DmFkgXZ3kzjlI1b2IQuaZ2qlSqmBsLy1ue7QqTSgUL
S8sVzmEyKySqGz3I5SrRELed2te7gnjA6ChiAFdxz6BFPukHrIfIrDyITXRHifwZyBqjo1gb5CY8
Wf91hqTE0sbMMJKv7sT/zMiLZcR0KMxTZoUnIYiz6pTQAyXscVeRMiPcWcQcKBtw8v+XMP93Ulp7
+04R69w3sPmgtBldAZIJIAGi/8q0UvIm1p5SHqFB0s+jXCcYlXcp7P6juo2gPu6hKFF0OgKjK6q0
SyxP/Bjlwy1Fuaf9W/Js2PctJ0yLEllAj5wXhv32I964JEafq4sHHmyB8CQAV+MjekMg7IZCAKfB
U1a+04f3nqON3/nG6hd5BgIrH4U/Eg/27fTinxmBz1l9thF5pUYGR7exZTIOlriPhSTxa34cKHHJ
7QSZpvIGaGnJHTUUvc2ZtH/nudoLqkcwgJuQHwksvjD+aAoOVrr5J27cMOlobgVqgI3UNI9Tn0XR
Z9sbVPlB9pEuUS6c3zYfbQpLrGt74zLldKv9QSK3VFdTPGYrczgsAojscTReq1pM1Ac6XQlL9XMC
e1OF/7mSRrwHvBomxhfRqLI9V3BBoO/7XcrJMpIyXiHZW1olpdX2q9sDJKuRDaDNstjblFi8hFHG
vvoS0GQHXIGcBlKK+kC439eYTxbgsJSjFqQbDjzY/hqK5Y7/E+QkyF5v9d2xvAMfPdLBTGCZMQJg
aCsu5FGPOv/pUuaSaQARksBAMcWQCE1khK63078cfNRetq3HETNTD7ka8LNM3AN1FNaJMOKcH2f3
zCtedTvbAStYkQFeZdZNSqlN6EbL6hJfdzmpZxn9CW1c9ydOTeYiCSmQrKBIHQHO7elqIAW1cnby
taXu0XPuUw8cT8y2zgUa5XR6N2ctPVGOFlPPvl7May7K5EzKudKekwvG7NPpk62tOKiugkVwLc12
y8zoUC/5jRnuqmtMRHR0HKZS0PBpZdIyPwnSBlaKLByo8LpbcV6u5+sQv7Y/GkSZaBWtUHViUclc
/YkKStllPyhzoRVs5xAjpwd4lA4d1byykG3XbFQMLz6xKnSJoOUPc5l0IjvbXHoztIiUmlgCusEU
wo21oS8mVtwqLB2QDaedIauzxJxEug6JTsW7Wo7vHklyZDOYiF27pK3xcxHr/WNstRdWwcYyGL0f
x1zGlLvDMCgjmvBgxfQnjkoyvk8zr+jCJk2sqy+EHY+4o7FoNqEP8j/n23lxqnguv6Xk9ds1hLIy
43rY6MCI0vONT62Yworf2fYXPGHbkghbEAznVaBhShJy/RHDAAJGsK/eKvR/YZaEejBz5oWY8WXY
uznkkjEO2My9QlSPkBciLGXTDDDqCVC9c25fkGAWNyxUdU3mKSZCcg3KCgMjwsPYFj44Z76CeH7K
X2+Rf6WhBAXkqKU2k9JT0aDu7JgF0rN7BwtgA4UvQvy2oYt3YSvgpxBjwyynJgMI/7656eDiEpV6
wtrVMxwSO7/x77Ou1HWjs9voBfCz0BaalEtqHxeK6eXNP4j9eNwIynTJgzUqUlO2oDvK/BPmyJGt
+6aNVDXv4EKLPPmY8PVF3o/hfZWYN9x2WxQz+ajASSYk4U9clfLpbRvWeVvs9COI00+LMlO+E8Z2
lO2iRTgOls/icj6fY+FForyWNWLCoHyHq/4Nk+j7DFVBVawRC5cE0n4dUGkZvYSNxLh2JQz/10pp
ozTFxFaxTZNZSRkpKlYdU9rtcDwyQ2CSA4+Qb+5ulKUKRnvxR61evEcQp9TQMlN+oz7EpcDA9cW9
D+31/0nHW3Z451QzniGIOUsawxFiSn6asJDpfGY7CMX9Ngi16ZRPQKaB11yBV8J4JTusYgHoQO7R
vVLq+v032+UIcVi3O/cbJpZ/H3FWidlPAFCj+seIoSS/NNs+HwAmnexzPiYDVZ/MYdK7uLzseXVr
n0lbHsMvWHgsATzePyA+flDMHo7hS1CepkLxA/EEaUZSzPZTwURwnSdU6xjRRJLVtDAo6HqGkCUb
GI767q8tWsEcnR0sKx2dDysKOawPBoHQxswE0sgTGffjHkT97a+lgNjp2HWsgq/0JO1pu1zJYAD6
2P4WxX3AYB14zV6ilNAnzqciMCojNbfkHMDlfGXcaSzDztOF4vkaGrWuncOKoO/QI8INhuUWY+Zj
NHgQBlXiPGr0M+v/TJflN5PI4amlEoYXk8pS9DcoWlT3Q9gOYu1OX9CriqLfcD1ximrU8q3u7db0
aV7XzeCyi1VCY2a230/v0kqewM84yvjdoR/AnmZQeV7nocLXi9ghjQmh9Dduuj4RfzlkvhpdVtOe
wvWLMH9QwOZlhNMV0ctZFi0ylhfKS+Ca3l2u2aDD3pt0oCWCHgVx4sjP3uvMQ71hlW/er3yzNefw
jQTi5QkTbmBlSMzbnOPn5ipVsh+UrCQcCrNuZEalMxuWEiS3Mw5Eb2ahLBd7O8ogyj0vg6fJFnd0
28VDw6p2b/yfQOLlAVlA91IxsuL+8OgHWK4XPv7Mr9nZlaiEs9PNhpiuXp+sfqMC4BsnaNE4WqVA
3qyBiDwv8+PU9fbV6W3L8mvWS3ApPbVaH9LvHomxkjdWF5RfNHpZ3oTnEa4zIsXVhQGUSuUzxWl0
TjM1wO2LelpOW2cFhe65g08EvdexLSdfZWMSCSsH1N6Z+Qzhxe6kdH0t9soYr5q0ztnpwGVIlIjB
wUljTeFxoetD2njgUeC3L0TZ4omt7DMjDcVkqivKoRlTMr6aFlBPp1TlUT58YozQYvG2DLwSi3Sp
ww5gjxXjoEX0+RXP6a71GExGwUohwvHk3MspeTuO+1E8sgKz3LzdG1+J8wqhjQ1uEQj9QFzCR70u
IO2uzcCjceS61wYLLEQ/PiFedBLeHp77XprazV8VCgFmX3yhymbxenBCDeDXnaOwRx1DfjApxHvg
6mzS3xMxkUNW9M9dJdN+mR2rSlYYYj5DmuvPSOyZSiV2/pQ08dQw9rk8e2yOvtRqqkpB22v5B55+
vk/5wRmGP6OKrM4xY2YwMa5BSFTQFyEKAAUv/VIS6Fr6cy7w6q5Va4VRix21sFSuXh1Uz0J09YUX
DTkisSV9+Rrq2Gh8EfR7gjzBTqZ4N4aFdDFWvmCCoYOOyedrheQyH63arOdQqj0tT8ogFYeF13a+
71VotGmgqKT2GQCp+PDaWyH+Jo51lzZ4GFdCIbb+qyow3jpJoZWIc96F1uZsZsS5d7Oyr6gInJMT
uMXBx5W0WSHevMeERg6Pt7oqxQIrvdUVPCjh8xr5gGOPbHYfBg0BPuejPU/y7AuvtL+MG8nbgNR8
q8tlt69obQtiaLS8u7k0zDoynhwoH+Z32TitpOnMNpHYqjMvp9jNQyiQl7Qw72pdxu6XAfYmnteL
iXPxHzdmCkveGf3b01kDejp4HHfhvZ3+xYwa8j9g+cRzXISxE+FQUQWoPSUgJ5k1sWdGJsrphT6B
o/Mt2udaD8qMJ+5C6Ef3kdl7DadNuvgb8rhv9DhK3jiA8ZiQdfJmM8+kOoHRGmxgDhsApys2hAGm
pf22fqEbYI5cPAkflGC+ECCXJjSZE7pLooKJ6VZekBtHExAdo2aGW6AFD7hkAZVOLar1TUBaK3bC
dApZDqyFT6a8OVipZEQu7hADA1S2xKPJSQRcRR9TMio7Ybn6hfN5C7FsGlcGGGaEt+oI7S/FMyxB
fIMGrd1wwKWuEdtkjxuHbCL4YejVMiI53JtKKk8FxKjVqEqVonIRwqxmFuKvns/6wQyRCEHxDwnk
cFV2SPsO5NCBo5RFZyVrHYGxnFJ/LXhHHfRU3wuROR8ic2H2gQ5UwQjGqPYJyOViRLvh8vmkL9QH
M84DctzRLzXV3iIm9qY7URSmu4KOXqOgup8pFuRmu35TzM6//+wk+YtwQF3OsTr7kVriaPcnxWn3
+zTa/L8cWh6GG58CYmKn8CfWMVHhSpSenyLdvXPVd6Qi737ijos1vLJ9yxmEXsrwYVoV3tEC2+Yl
qPeY7HaBngGOOkD96iNYCKXPPWRCDyUYULpz3c9jljBQGNgwjdl2o29E9Vi7oH3gcSEHPZwTY5Lb
xmxRON68tM4mp9088N2CTrTLtkLFRDaxmVfsN4KTZgn6yBRL2WInHgtpGoI3g2aOifnzB3PkyoEf
9SGV7WKXlVP/NQ3P3oXpXMPeIYvaGKe/bg5PtWrKDwGc39NJcv9zV+u3VtYp6f/j3CtZOed6v242
Ra3ZMuObOSYHkF330ilpLPQLE2KmFmmsqN7YeOxBSaUbnL/uUVU7hisLN4/5OdkJfLjDwxpjrrQ6
kJd5bfz1gijlOF1V/MmaDdhBPoWR0hWn8Iy0CnHTvPURJrjyNA27ZifxEzJqzgjkKioa58YkSyBh
A4EQBfmTLR4519Vx0hoI7VbOhxAS1HVdTD1r7yAGxBrALX6ZMuAjsfmdULxXOmo4IUbunV4i2YT3
ptIeSAxj3tlgiduAkKw+cdo3vFxtvTgIBZDPdxQJc2n3gbEjPo/AUyhUGEQIgoGR+HMy/LajrEvA
EcElG/l/S7tEN0a+rDTj6WYWQ8BQLhbpvHyzVMrgv3HvAzZ0v3enfza1Q8anWG+NPOP8FpT/tYGo
0FI2YBZl0yNAexYsULIkZm2OY5F5gwyNmqVCZHU1+ZJeGl7cPhplkPenY+MFa3aRX/8BMHeRDmkS
4mfKUW2wjWHJL3yZ/U2EOQ3AmZwKC/ax9uK5DrQ14/xnqBWA2iH4um4B9FLh/1CRgbrrsJtngMBa
IkWJBC/L5GSCQhDBlciPDVOXnZ6YRi90G59BoRIO3Y9jiMyWxt3tZ2rDwmpPRENhBq2POXXZv/so
yeMc4uxk9p09Kv/+dyzxZXJllo+VkztwYdj3clqiklm/EuuNLEsQfvFq7zMEPvQSrUvsfyFd5Dsk
++VX2zEfSq5vbKW19rqUAvxJa3NvYm8qbTI/aycWh909qIqtzrWsGjpdojLAU1Xp+NsJl5NlurCz
5MZE+nY/Lq+lbNm1cflEySkYvfPBfgYm4U5ZolDp4NFGiBre+WKn8xxqknOGf/YFM0337n9gamOI
+G+QyQNK22bRAqDMfoBBVOP0uqn5Lu7PZkIcuwL1y+8NtPD5HX6LmT7vcMulCzLGtShvRD9wYeyx
NgN9qAE/Mez1UlmGxDGbArcJTXgUDVCeaZxnxezXpntl2jzQxwuXK0si1mQ+G6wKqRbBJxX55A46
KdGlCVvuwPIH9t0kfDFrF0wlyKF5k9gaFljjLuIWk+F7d/nD/Ju/b8EA04yFOGvhka2zN9M7E0IB
ZxsXxc6NreW+7kVhsgpFyYZrctO+oWBi1/BOFHNO1v6CMGpPIlR1yrI163j16YcUwbYh8p2a4JMc
k0ffc3aRnv8bBFWsgEEa2rOifXI9w3PaeLspVPiBgCL60rwz4DkxlKZk8PxUumrkirpJey8Rk+TD
VsxKMIa6b33e0Iar8bUmMFJNnQ/bNR3AEK96NXX9fqwR0MO4E+iip8mhHWDem25Kp+Xf7Pjovtbx
NsGyG1FzCFHrAAF740iMZWpYP6HYiqxUFTRFyf1yvSJ60XJe8LOYL0XYzx2vZDplUbPXu8NM3cFG
iVP7EEoK8ySxfqUGyhF0E3oz+0WnsiYs0jLdJ1rJUVzUJBJEg4HmK77iFR2Sj54ncv0qFBGjy8tD
iPXUlFpsYPNFn3IyX/6NEvje/ltk7llvWcQ/ZLYh8HJ7F0KoYjvT/iRum1yQQlVzOt9hUF2ha4T8
VqoNXh5CBERS4OWtMdwXkMV+0HU4/q0M63OoUiF31fBgIy9MQQgOg3gWVGdWu15NNgbnRooVc7Rs
nfA7bSw3j3rLtcGtTr/qS5Q539Z4c3Ie25in3y7q/7P9Sb9N9PxlPnWRJKabWMxTr+Pu4bRdXf3k
ht9pUlR0PJ0+O0W7Zr4xUjYE1kzBep2dIHmNtklzkwsTc2gynIwwSuReP9kZKghOXbFSHP+t38KE
vUtSnJ1SKYJzwAh5ZPUt3fW/z4+Iqajo0tl0cXTJ7BBg1fdBFSFw81A7+gh1hLYB84k5XNaH6/OS
OywEWeEVcjj4smwbmXsev/I/oGixy2470LBROGWZrPTywBdJ45zbBP7OGr0X3cxVXp+1n3Zt4lp4
capGGB03XCzD57/HFAQ/yi6RlYafKvdJxrg+oklZNpCTKe1IiVRlD+RcgnVo1EB3MOnIikE5DofN
hLfslCSZNH1mD0czzljTzMd2xX/SCnChqphAmrEFr9I4BAYdeiamDKArjnwDDrl9eLQjlck4Mugi
gVdlLNeXlpESV7dnXspuYQK4Yvgg08/Ozosn4zJAc3ov4XEokZ1+pRUq4ZNP4+AiljqxVbsfAiQl
oK8w3wc2a8xK3cl/lUzFEXRav45XWgMQbnnAjcJeve21h3Uf+lFfReDNTMdW02/WsdHr53U7ROK3
1baiB/V2UxNzmEBNz6uIVzjMqOwwkPLHzeyyT8ZIBTSeS9/7VRxwOEraNhzmzGMVK3rxFNvaoaCq
tFnufVZETPPHcEEWJS/Vr+zjdCd/yAHg5oELgRngPhCl5BQ9TCWj2dV1KWzJFkNII76OthMyZJ7J
uL6UmEquM/PrgihPJzWXvos+Z04JY5FhPDTZhKBN97wQvnVuTeezFTbFTyWdy5DQW/Mmqhzc7exC
CXqrm5alXisCA7E8BBEQ1UaZH9PFKOcXurDFamsd7KcWtbtsg2FtsYE8D36nCjBar6rVdomrwfBZ
Nr8mtMH6rM90cdhN0k5nOdvIO95qApFOMmBrNIPBjdhTxVgmZp09YF3TIyIFU7wyNUWTgqZuFMC+
aYxyTH3Hj4Oa+n293DPyZM0jrx7bajT6b4GmMpWX2Rg+H2MbIXm4eXjGamjO6gr8pVwO7aSrZ1l3
j9O8HQ+0z1uvfobGgo81fiC/QMofUzJWZ0SrfwirSLIgsqZR20S3VdBjKTiX+2Ret0CbjCYQCP21
/gPm/Oc7OXcFiwr0F3uRAaCkTkVq5W4Lqhlf9SDmp80rTnHorw6/ctnExnUEbhNW1kp+qcCRYluH
WBHjwDL2ut0z2hMFIBl+wwGX9tdAnQ72ghnRyH/pCX9FT1ehMnJptF6v5aYTfAEro6ffXoAbUW2k
1KwU1fKD/E9NDABi9Z7vIMadK5NI/yNeza1LSJB7DGvACyL9ZQRL3kzKlVC1tAX6ANPfV/fIvxAk
mjVonr7zf97+0YaHGI8yFMf+a2riLPTRtwpAVrX08ZmrAboLdkhtTarwDitxfvuGmf3oF2/Kjjgh
u22sx0+YeZz8pNvsmSzVlz8i5gxh4yjDXzBopHuOV0CE2bwc2DJaVYQAOpJVJy+kZEeCog4Efa/b
cYwie/CPVAXvXSIaPHRK4ytBn4J0hXHCemYmk5uIHa7UmN1QEv7lXU2R2msGzlvxOdkfOlEQiZos
FicazbE76NooCjihJKFWYfPetBbh6oeUDelwe7jSl9vPgyrGnwNOgZehZQZlNybaAgpstcme9ltx
BPwSMl0n9zMGaQ3RFr0zPYGV+w7L4mthFfzV6WdJ4IrZAMcjyHmEJyvgUgoBj6NEDOBsgzOhruLB
fvuyiCl+FVObVH/P72O95Itrk2/lC3qyWGOu0Psra1/elyWU0DGyJmCMak/F632BOFU8JErsGKkt
at4pKoP9yyggqJRTyBofmQUiSLDHXQR8hIW3Tfa9P9ymG4wk/hyq4RJ1sCCCqKV5k8NU6NZ9WRMD
4ScfPxHCZ91JVLrGHY86dYf5WYjOhhpJ6Uocu5eBD2NNcMUoO/nwaybVhngrKiJxBNMy0xbGnkuM
dc8DcReiXriezQWuWPwmx8GSfaOxUW2k0i/CwFYwjOw8RvBMhowhYXpA32m3q9BoCvorz4mh8a/q
tbKUwMfCeadH7v5S1Eil7l4Efpv2bKn0ogKNqlMWV2dk/XlarC1bJqszEMYoyRXTvgC909X+8nKV
IPzsP3UZ4rj0hcFrgXfOKcight1OEaM0C0DcN+1Q4s20hgHWO9V07b2Lif1DJXFJ7BzKAnFyqWhE
DHiXgaTY/IPWlyeoWuI/dGKmdnNVsjyk6O5tMn8FlAS9OLj2xVo+ui5jrQLfV8NyY/UNbqnpdF/K
6j3fSdeNgTyiAExDCIcQ2VngSJ7gD7LHBGunttn874WQ66yJS9VxSiyxn1pgmCjCX/BnoTLoEt6P
QWbWdVevFa9OmpU/jVXFe9Qk6quzymsV9RbB5WZnIZjI8EyFNUBTMaaPyj/qt+gAoPhfdUyHCCdF
n0qM7GSwx85dvFVLOSKwbWYUvwRF2FYlJw0lhh+/UBxDrLcT0T/7J7f1bdpgfviYuujjqRoxGV7d
9jGhXb5Ii+VpZuTs3jsJQJM5B1A1Te68LRqMBHvtu7mDhl7FOCOwem31RdfWhOHQHrXghd4DfLbf
UFXicGdYD0GKRHb9X8cjpZLUZKxuN8W+g9hYyfJPgjn52pBT/4zPI6N8iOkYo4cGr4npTgNgPhuo
HlawwcW/8vJpFG7CTCYm2HHz3hk6Zc+9d2jmjZpFdNeZXY+s+F67p+ncQH7uYR1ipPrBCY+6ANuI
yDTG7H3WjKaqXWoDZehdowQwaaIOOIe8gaNUtlGXGukENBtbIgGMMH31R9TRPDxGvtZxhq2YCNSt
d1obS2xGo+jYPYiRklMCI5l7AUDHcMmfbrFIBfEyU4R4Kq1H6dqn5Ggbqj/+b0pIPzF7Ih47ExH8
QFNhHSbX4HDtPKlxSy26Ey6emHnfuj/xpWqGBiFc0EGRVUb+bvl1VnmXb9DUvM+q8lp487CfLKiJ
PpaH34B+L4MUQAD9NtbvfLxJvBDM7OCs2yaq06nf+PMOfqL8lPh72339LjRRLVbZVJLnMfOygxzh
NxJ5+45k6pPxye+N385PzmRp6AubuaXrTsRacvzRTbAw7s4uH8JXDHwZe2oHQ54gRm2iKce7Wfc8
vrh/s8/x8miS5Uigt2M/IHLEaAY1JNv1IPOvlg6Gy5QT4R742or0RO0heCe8RU8Uw64AMmXomhaC
7I308mbCDJSSTZTcsaIVwFj2HKUT2yfWX8MHMR1jtQ1b7PW3FrcbsH9ftw8MeWnmpVNTeIg+ET5D
AcRQkP+3op4IU8OhVbWsRNu8GF7CEc/UjBTEwtGxeQpqOfZ+8Z5T+4Llt2ywZTR+z13Jlx23555O
Z4QhkpoO+BeRRaOS0gWJYcrGgxNxJclS8H87Gg1BJtuJ0quWGx7RU3g1Clx4IDkxt7E/iHdDFvAM
lpuIg4g84enLt1O5zONusGUZx/qbm1wHLyjTs4pWxWXHhwkGhU0xCGP/QndQXIuNOnpxGQLMFOI1
mZQNNQgB/59XSLYCxczydoqWux7T57njeYZrGx0VkWxfm+NSI/o0OSBswPqkok9EMdZTXhA+0d7f
eeMKvE9jYhRge8h1lvbyRY4cv+5sVubGexWJACuGkTpd05MwL5YCHgP7e6doztT1T3M0j3jAzwYl
9ptsnAImkp6+npbnu+pCGnIn0cc8g6xCbkp5YfYFBUWauYO+caszy3thB292AvW2D9MiMTFtFuTb
Wo7lTWvG6Uh58mLYT6ukbmzgb3weC+MHmo+sL5XLg6+t9Y5RSwQwTAHltkjvpShNs8eSzut2mygQ
hG6zbldPQkEx8Ly+af9eOYj8I1ALQ5fYQEd74tKg79WoS49XksaulUqSZoBza8cV/Ct0kM4ojm7D
vKFnJZeu6IymeiN/9H/DhXjd+3RhKikjh9NG0uyQjDzcTDywLvHKw4VOBgRg8Tyh2GwJBQb3nCal
Inrh75LZrCtZAC+IV480yEVzJswEVV/z2Ur91YQZwF/dryE7cYnqXaJiGdw4APws2+8tUknd507+
Sy4WdywIiZuBNWN3W72yM0aw/3QZ1v+ymaOvGmoB1YTghxX5iQ7iYI1deXlr9P50quW1yZTZQFR3
UdbLvH43H5IjyXx+yncAPx8tF1z7TPJRcHWSAXn2qfDN31R14Sg7wqoNPK9guLm92j6umrfLbTBt
AxeaHBOCkJVW41FfvdIoRjuB+Kg2829sdUS59QyJRSO/eZNiNhUiJ/ZVkzDGsQg3kBbGyuK2FogY
Y1e3P8Y/p8Nu+vXBNBqSDJVSBEzQ3qQUKQk5ldV4GvIzQH8EIxsUa2EJv8Wi/N5MbGYqSy12KY+e
7TBjKX55uHpc/c1zPQ1HSM25dBcc1/NZ7BV7cTevImw/yy0it4I7jOHMQoztP38AChlPVR6pUS1/
DbU2emZfHIZleXm7nNxWg8chvYYr7Jj7XXshBKXs19oUko9lY0AQQn7klcF0io2OEmbr8rXS1X5n
hkErBHTaE5p6oM69rcQhRgF84/SMAePxb7CIjUV6hlwLcGBnIkiz/bGdrh9NszsXXSA3jCQkv8L3
m65cRqmv+VoMZi63P8up/FV1MCub/+QoZnQsu6WV0b1+zQmpwlOsKhf6kzw5Ndoii6D86cAAiZoz
TxcXqZ513CTFMBBsuIv2xOsUTfdk+DVEELGbXm6LHr8nyBrVFoPaQPRfHynrWcdzUuJbcAwaWi1S
O1VNIj7E3E/hORvoQqGAlYaKvWzY7McuLVgdKAfNU0vpjU0IUrf1QgEwMMvlKmHOW9fYwS+aoyrW
NaAoKsmLbL3htU6iT1NYffN75llcqDBBC8rXebvE1izzp0twmE86KL0B3WXHRIHzxFfvmYjayZ6K
HBohOoADY+omK4FP3nzIq4YEExOPPWHjv77MvIiftoRYANLUxgPDtxiPzoaX9IGbtVd2V+OMmW6N
kvS4C42RnBSnX7tH/JLEGEeVvn91iKaZx6+LlC+slgn6Byv97b87NUaNIF2POtEfmjIMTuLeM9ex
F066yvvUaM4T2J07e/+1IOF7CBHo9c4QvG5Tmxz1edo1ocV0Hrt7wSumb7LdLOAjNI5mQrU6tgmS
fqwOohu5ENc84r8nSpJNpJ/GXhz40Znzrx6O7fAYZNRiT7aEbNZLolUb2N8f9CDbfF5+lhpDFR07
oWd4JhSOkaZCWf1GdGk3YL8+2G+doUO34KB84kvD1rZzR+S3RGSVWnVpgnpG5sHkrxNyStvvPCw+
ky+ADwwsehXwsuzGiboXyYrc1OCQdosUieDi3X7FrWkTK31UqDPKxrZR5WMayCclZUJZ4913wPq8
jebxp4JhXvbgD/3+mzzzH0OryatXRyyOFSLQLQM39rXwXPrjoS6KKhUOPKqjtor1i3kQuEwMtXy4
G5WA/Z4I8vCR+2P18/vz8OwU/IxN06tpkSOfIIJSJIR34XBo2rCD9BLUwjsP3IX+qehOlD7ZeZLb
n7DEuhMFYvk1hDGwMopNkDcFlWFJxBj33tM3Hx0Z4bMe2XGgoCult6lOdvj42RKgBtPpT3YiCJu8
LO9U5sBftvahon0MWj7P/Vfa4i+xau35ABMoKnXbwlNvCUq95eCAQxHWVbReWWe2zgASobEVowsJ
eRO5/44Yl/Moq7oAvnA+dNHVOv9URM/1K38wjKGW+3xfTUhLnzzZ7cQ6az9b1yMEkiBe9uESNyjU
m48vdlU1xLt5DWm5QMwXYOo4yB1kGnenSV148VQ6nMHkVWtyiP2Eaq+23iVF0D+9G5N9rEv5WbRn
CfcLDnTBLOLR9cQAK1adaE2QiOheoCs7DgU8ylH7lpuvzHU7pHprU0cyg3LKkNq4GysXkSGWo8DD
/8YPXmDe7rBmwBZhysUxBh2NLer5Imd42v9pV9jTu714V6u7mpAPmz+R+IsNOsV9FuWc4AkuGB5y
djuAVrvbVK/y4BtxnPthzL9Aay9g+4BUltD4I+Zc4uemRauMccWAeCxkf2Ypc9F2PhmexvmRpWbI
fs0GkSvMFO18cXPMLR+RZB4g0uHU2pkDEldMz0YZWcXVEjxROmo0ImKbEg1eq9uFSHwh22+eS1nA
TzL774uI5Fv6ZDn+cMFv6Cg3p4XtlZiMlzeqd+xagdnIZph5bGXGGUZnuqFz4UaAneqc9yXfUtLr
HCS1swATxVMBFJ819XcZhw5QSL+h5a8s+Ry7AnYg9gFMjxlL5FbwrK8leuZdO+xGCXDt/UClGQuq
28yIET3NF0rO6lwlOKO0NZgWIApLdx0j4mTs2vAtbjD7jraLUse8AeS+60sT/PiYhkKeseI0Gpm1
IWNl2X9tabvq4MeEo52Qq26ndoXvjw59pnJEVIUYizw80O/Zt14aC+Sp2cgyG1V3IHfGzjSoTsya
Cb1ieJUMFuNP+p3FvqSivMowEKfBPCXeqX4w1+ghyP8IbfEhHQXqJMO4YIzOkF28EXUjUKUB9yg0
Ql0NI6N7UK8i7imgGo652/0cItEksXTbP85qAWtKd3EIbmDobm5un6ie6FwbrbaeK6L37VKat/dz
sB005Q2WDoMWqzJPLZvMbXaps+uf9IyI5EJFKbbuKBCWiIPgKQAe80lxk/zOvnSx/iLU8gf9MZXj
+OYetKcB/dUtsHeXtwSxqcKibGldG/a8KYsclGysbVzBGKvqXikDn6+y2UaB8MYJF1htgF6HxcCD
8URvh2tAK2484H5GxJuyCUkwtjZP8+jaZ4ro29jnBoniXTzMzCP/O0wI7C//N9qu6QvR7AuWlbOt
irU1ZpcLtafEJLfW2KOngl1SJ8bScpAdQ3ohwvm+6LtymrZtlYw8VB6SFPdyg1l9QGqV9u3T87xu
rgFf6uL231c9/Zo+xsBdh2vl/72z+2NGKfSzubA3E6F7zU8Mik8jhVyymubt4ooFgDZLSHnUKpLf
hhAT9ZoZ8fyOS/OBLjZZ1jhKdQCesWYRVX/voCk8DHKHC6MVgNMZdvrM/I61jcvwQiErQR6OtlB3
95JnDNWU+kxsLtt9wJi3TzSpuZXC+j/aUvBbyWZRgUrPeigGrJYSb/63GsXKNGUeK1Rcs9bQB5yE
+Cf9qB3146tZtykm89zehf0q0/+nxf2e7yFXDD9SoieqayPro/mHRBq8QGD6E6ueoW4MVjJdtcZp
MGGawBmBUfg4Mm+Em784i5Gm9rWWbFUL9MZpPeOD8ow3aMndKmKM/Orb6Oq6HbY9VPjuzrqo0IRC
d7t8+WwEgwC22S40RK4Lk6vOgllGRCw+eyneh01XBI6fTqdj7r6idX3b2OkXZRNYIUNqLafha907
+ZgrcGEHpHsXfnj2BsZjjz6vAFyg8v+p0qZhWQ1Nopm6/0WILx1Sswc+w9S4s33l8M1HR2N5NqPF
wMLiMYAzYsaDmrBSlBPtyC4R6f9WNeNxraTf5965WrwYcLJGYKuJB/1ExrJMg5tcy+Di72EHQgLX
Wsv44DsA7F93eQhCfl/TWyq4FfJvlhZVeq3M6FuRI3Rl+D9bL5uGEfrGgeIiCM6pn/IW4x0AcQr3
KoyZY8EknXGgCvqEhdbBKIj1npA5MSfaAtU/zsKRRelyIugevgwdHVR5YIrnebzPyupvz9AOeOpv
Ovtkfe7dZmVdQ92GCjZNPv+iQ+x4uSzvV1qva/9UV3s4VpTfH8Mkh1slOEIJxNnDa4bueQaFqaog
3YV3zU3OBenxQOyMtc2lkdjBOvtGboyBYfEwY74WQVfN1l6VT71CT0iacGmbs2f1HYVE4v+CB6ja
Tn94uCaH6msdMwxRVdvmeCKeyKFjCtQRKS4BlsJDFchnIiQkpu5hgxPUa/xIBHoZqaVyN0bKOKrn
7xnAvriU5LW4tav3G+smLl3j2LBybk+Qq1iz2jzrpqB7AAVIQOPCGBFAvNw8YcdP/8KLV2pMzSj9
FUTw/5qagtzFvdaaFNQRqJ6xPimh28ocIXNVndvGRQBaB2dCvG0G98RFUkzWJhozdhvIkq/atFXZ
RvKueYXiDJUMGfblHqldDiz7gsuJ3aG2apBtQLg2egQs1lcC7ttoNqpEv0swbFOCfrKVpmTnM8S/
0StluXCWZpXmI2Qyprs/QU9Y1J/2+It3PY0yh2xJ6USLvE1/PFfeumstneMiQR9cHGIoAm5obT0u
RdxjQTrghPf+W5OTZq0BEbe4jzRfxCZxOQbbNAev4mdyllT01lbRkw2lPwk0FmmbkhLG+AOA0M1w
m1TmR4lzkhsKGFmjMpFtIpvUPQGchrJeMX2ilHoJjMNufcoMX3oU0fH59OOAfO31j8HIbk1u6Zm/
m9BMTc+q/1GWZnwwmSRAXEJxJA6j9JSfQ1xBSeBMQsgeFwAocUQDe3AKrAvH5OxGzmuj3SLDRAtw
hf5TASLKsOwZbJ0N3wf2KHsq294aYdFXNMnqqW6UU29rF8dt81n/Ah6Ntig0ymI3G8aGZl/foytz
X+Lim3idRvrqQdqJO6/rtuu53gETmqoGAkWUGD+XGCItR1WPI+iywOUn5qZlqHBxmKa7oS2aC5DX
NTRy+hZOKCGx2Q9krD2ez+dOnXiGt2SAOWeOTrrBug3AiLrUojqZZSXcYP+RyM1QDysqHU2RW0GY
1qF87aCXjBuXLi7heGXd0adR4YBDdLuH0tzPmPXAh7YT1vH/tlzKIJMRSknKRZ8ZrFz6PKh1dQj7
JBrmZ84AUACIqFpmkCu0XTpOaGPaenPiWnskzDufAxGu+NxjFhNiBxxYTlhQbUVbPPVGVutiwuwN
67Vqm/e/ytCoptS11f06VEjFTbfol18J0oUof/CemHlM+1TmyojpdJYAGX0yVkSyCc8HmkJM0oiq
gpNnnwzmERn9+67KS9nKP2Ikot4TSQAq34ngdiAidyRya7x7zQ+CyTyHobg2sCsgNQ8a2IO3P0AK
QyNHBjdKQdSc13D0wLaeOa2OvRAtfqo6PZ6xXKgJ2p7mVKuFPU+UAHg+p1oyCks+p2/ZtyDohDIr
JbG1Qdqq0q4eo/7M01MKfDp+D1kAOCWmfibjX2E9HsffFk5QwMZasVSl3wHJ+hmPtUw1uI3TNfU5
O3t33LBmGmDR9K62hlReNd16VI4/Z6o4OcS45N+8romcNWDQsJ0ODUzKMZQMX6HHdbjj1LBcZEBI
DIvmhdASQys/1IrpRtim3LZT5oEFcxwn9GBcNxTj199td/ir8TEn66Dyr4EiKL4k1lObCZNia+6m
+V9VevT1NVlUvboaSJ7DdZekJFVwGIYuBK66N25kh9zOk2AzVcJUTJnhOgwI2Jt61wG/r7z4NOa6
dmZ5O/qDaD3TA6hsavEhVQ92ON6VLwnxJyCajNhzk7Ggcdkrk1rgAQ0X0XLVCNwZ1YcQIjG4f2ig
nhUMG06sn1ZOGlAvrt0ppv8G6RBA9okVC72Hf0VU4NAHbA1uirjhMd+T+KCNjEyX0FBrEuL/ty+K
ykM/eBLlRts6UsQBJ/KvPOJm2F+A2vCnpNbCq6zeQK2HBjJimJFEfIXdv7QgnzFNICUegzz7kD0x
/TlkTZGXbNSwz0ypenY7T7O2qb1gqLtvELR2GBG5taoyevoD+KttSZa3J1KCh4+OtnoCBCj7E8zz
ZrsHfAwV0/j13XCooEIRpJZ7Fq/9A6VLkaf/tZUPsDcy0f4e6QkwyxNDhqyvSVxj0V99RjhxWzn3
a3x4ZYkU+r0J4HRRrNnlzdjuAfHJLpQ0iQkf3WywNAdqvC4jutN+NTgjj4+JIN0DrzDNCGQBYpbf
u36cYxAlUsXNn9QU8y6a+iFFC4Of0+p73EqZ8vndOTiw2etKBzPUGD3bd4l2tBlTXO68OX7ECBgG
nZlzn1CC3Jpg+fwxvhWdQ140l1RS+6QZ1BIte+N8pEQRHRrGqjyJAdXudyKWx7tF5UlHCbSfrBgk
2QZq7wsOMF9pdPGryhKa8Uwml127j0IR13RcUJTrh6Ne46FH8UMbg2He8iHTTD5rpUWhdtzj7bry
R/R6LGdKzqcBlhC22YEK8mqh72OS4YIxjH5hratcxCHw0N9ElOf+qIv3YOQ6vpCiX9H5rJKTS8Qt
CQ2ixqQt2H83qjnYS7SG9iLgPEzeSvC3WM3+boF58pVL8EX/If4Olr1OOXJu0xLA8x5SfbRUFOJy
cXt2XsOuJZCxo+zMc5zXtAEsrq9pBuk6QSmAlQvjqDsbWooYczaAhcQ2A+23QxW7E/TEWCg2W7Fe
BOQk2Adk2SKCy2Jql9yVhutjK65V6ZkxjK5dVzhsoeMdLq3J1JqKjLk8ud3NNHgQ5rBb9DQZJ//Y
rNCJcT9KaIqZfqKCLa6BKQlY9XwiONYGBUuDykTYAPQ601xpPVTlz0k6BvvjdJ/Wsw/Zl1nNhZO+
MfH6BTlxpl9lNJbJNKuH45FIawCaM4im5DOT5OLmfb9cpjhzqejmlUkpbnfGJhAGLYh8hT3wdNst
GaM3AdpIWZZ01UHx6UNXsFzvHpkTFT8ZZRpNTusGuhreklMR1o1rdHiE0CjZmIs81VE7qO/Xupwv
JV7syidVpvX+QS06ZwEuOuC2oWBuQEiecKGvxqhOgVcjtgZ/OXQuK0BGxBAWD1QJyxtB2Jbcf6EP
h0cl8P73XUO/4dzvrQrfI/uF/aXB51WU1jHNTLgO2EWqfs2LyUYikLpzqK0M9bfZ5Is20TmigUrg
JMNktm7IorBFBb5ZSxlZHoe6fuAxZn9YGvngQlDRQtV0rQY7jjy3TJWNcrhjI4X+vemwucf9EZ13
ckSCox5wDGAq/6nP4sYskLYL1WGvShU/iiI9L2A+KRzji21pAGGX03Yz8kzEUWqN67DpzuHCAuJb
eAtstxGZ67GH1M+16N2YpVgxKzDOwxXuSKeTF10JQ7kntUHn3dIBunUF8Fw0P5YLUcwDuLl9ynBO
E1k3sMI+7N/bo1FaRIiSdZboB3utwJw4E8XxeSxWFY+1i28xEhQSb8rAKwGBrQj+sbvvin7yfibg
CO2xayRRbQU1Fpn9YVX8sxF9O56ZFBljx6CdBw/+P0PzLT9r0mYHZixpStHl6hghcmRKtHy2Tbu4
K1vbOC2JXNqgGAhYPHRAbSUNaGqKYQUH94i01VMcXqIUkm/aQXO0kcBpB9Fi7TQ6/k4s3JqVL6fs
o+4dnMQdiDbY9Mn3scv1+zRGKYyITvHnAmwQuFBQ8w2PuS+oPrTrI4Szw9fsEE+pjOUzrRVR3/jx
5/r13Uqs8uZ/MzDFroaIj9kl2/hFa0mghCBVp87s/JYzAeTOGCBlPS+uIQzC1nbUcHsxx+lFu6Cf
55cisW33npyMx1hiUxfIs5r3ARCVJThrdUTlx1yGOzDL7aEOu0ANw/fd6vQdlNuek8Dsim6dH+fQ
wFP6ILA2Xz3f3mwqayEv5cOCtSlhX5tgLfjDyXVD5YFOBBzsAPJ2tGNNFH3O3dFTv/CoO3ty6trm
hNZt9EDHGEmGgX+FZtfgC2npn6VVO5KkSD65pxS/835uHnjszeXVL3b1S6y3F4RgHE9BGkngiiCq
vq2siH72yPG60QlA6XUa5mv+RcV/lmZ0zpPBx+i79OYLDGC6BRCvvxdZUFvruhRdjnbzx+kj4q/r
YSj29UDTQBoS07hOq2JnRotf/tFvHCjmdxXbAhJ0+/DN7MWMyh3GACV7bYKiy2YuGoqofkt3tdlO
f8WVlm1ZuQv6uRoMcA4YiBohxZrhAtcUW22EV0zAc+SNrgP38VfEe+kzZSWsY+jGGi/buq45viLD
3ATlCZORUGj9BMIZLzEjq4FItqrdYrk/Y08GVPwtTTXaLZauenYFeZnceEMFYyTP2c9x6WFeXVOh
UyY8taSYr7odeeh6f2U+4Q4uh1HgK0MnWcikYvrsSlIqDKuUrkuInUy+8k4Eo9UFktUr6GxiRcwg
pLPJBZIrRDSR/IOcfLFjPUfDZE3D+j4/ijVWDXE4FUYNkUaA2WTli7vw5Nj16MW+HNNOhNT/iGE7
ye3R2SqWQt7GzSQWcXlW0tHARxzFAGazNyy/sTEr2VpTxUklsEWirgkB3jcV0x4/fJ556ukVJtHt
7yYgSEGORdg3qLhkhERYNeKPu9wthnJ1Bz+53thUQLiC5hMhsKa1DOD4w5kurO3mI4AXRO78GPvx
AN0d4HYDNY77uSJRYI/iIXlubG3hPTihuP3KNkwSPgbAahqgw8rSCI9Xx6N8Y2AH5XqjQECgsHkr
MsvlV9wFR/3coY6MAyHr/38Ih5Rdpda7LG4nMVu55mYKG//A069FNPGTB7Xrl4dk/g4G/yoHXdnb
KEYcU7LfJ5f+syITYioCvhgaCCxY4MnceLVV5UawIFwUhJ8BoxR0nRZ/OR4wTDVIDnAlNVxHH8Je
vrrHzVSwpHeAUWle8Z4EWThFIgDia99xR78zuBKASnYOnCgA4QhtJFGw0s8HxlKKIPuBnQiHsK2P
bLtwvvchzoOz2ZK/lrok8PMCtgXVWZHK0P0mCdPk/e7ZyKT5akaZwpR9bQxiGkFjEBewxhgze45K
EO/bZArd4Kp/uVr9hsQhvjxx86znbEYWoPl/GIveyfCTgtGcTxAQhBHOwexV3iG8XJdqZeIMfg5Y
4vNqOjHbVhhV4fAyDnunpu6nTn0LJ8DlZZKdiLzOCYLkqJB++Hi0o1rfTFwO/WlObRF6U3MNodTi
epjtcR9LMv5IFkY18TYPvVXCgPnp2J66XTFjxPR+hkiEB6MuHGiW2ifpXNXfsilkT+rNlch0zyE7
zzM5TW/7S+UYP5GjW1XdS7nBEJ/i4f+u2jPtXnqJ9wEYSdBRjZlswzHYRXXZOWCIxpDdH84OHZUO
8SO3rDlSI8aPR4QGZDY/kwGiPebgCIrznyQjqtzApZaiHYUUNqW8qS+nhCxrdpKBLn1d31J4s0/J
STzZdj2/ax/SIpa/7IxzRWka7vYU2Z4Hjv+bN37qhsIo6cjoNiHXW3TiSJEE3gsHbTL5DfN6531y
t5A4CVseytQiE3j07T+rdrfMcfFzPkBDM2ydqFY1TogY50ebcf4Nb7ZxsD7WH3SoBwdTN28PFM5A
3RcPrPGln5aXLMm6rBH5DKTTg3Zf2pRrsCPc2D9wLLu4mlHMwexgwLa1FKu/0ZNSvlR6G22J4ZHQ
XmiAA0fcKeV0ahexpCMIkKOqLFNn34svYHI4gL6i24OP3hD5Uen9Y9tr3fg9sPha3tb6tBJi2oCX
/1glR57x8t6zgBaRAxTpwYLUVvONqakHkDxQ/U94d8m8xHCG7L6eF4EzF5nG9UWOx5dLqLQuPDkx
vyC7bLcfZkpnyZ1oiNbnKG1QKn8rSqspCSg1Jae5lXqdL9YL+aPgGeezvTh+GZrVMKKttZ6bB1XJ
potVqQiIQc2MJRobvT7hJzRhzSas6H0fGwK8RTB8MtxmoYRp8vK7ZJuUOghVrrRZfLU15/C2Hx+h
jEN9nY5WBDm5a0JNkB1PsxUI0n6Lstxx6ihCOlPDxLRYnQTSSG83+tVDzJdtVnX0LebiBZKBPm8+
bC/jDHH89Nrdxs5RbMca8inFBxjEzniQeJp99LGITrKUopv0jO8VsCBfAKnxX/OXQA05ZYprN8E8
OqSkPFksdSDoydROPqNHifXVyWBkacGWaWzZIhhzZR6xohmtOLJ82TA7JHFBfik8OmTlSU6mEKCA
Tud6AG4lBVq6wbldRk1FtNO0DPtt6asebSPqJwqflXdyHo6GGbFCG11u0R5Qwin/5wRWsXy1WwSJ
lLNe1H3idBOUz6f3lblzxTWIDg5XEWLpf8jm7tK75M/om8wx9QDoEMNArtjpvs0emNfyhjJ8CaC8
YyJVyzCOWS0yaY9j1s1uYXrqIjF4vCTGvd0WnawXgmzp2/c6NHYnElQ9v71le/1YfQQ3vNMnkIMc
qlLGHqBZeOBzA0f54KKWIk+XqLL1sI3Ssw8BuRH6W4634Z4yzZt8oROO1IG9+9IAYn/rb5Z0tG8I
p6zjosAyRxeHC7DegJGBZq6fQ6l2zS7YUkz7DPk/vo9npWW9IwB5OJmyFBHW0aaclxkfpHIs6zd7
7GqllXOtJogMmX+u5OE8w/WoP4Lxwmr8jOTbK6yJj/GIQczoVpV10MgUOxFacBEB5IKeXsmRErOs
31Q/rHVCJPxt+j0mwjBqYto1HRKy+3wu368R06bFFkx1J3SmzVx7oxfDHvv1h1sXVuaKenOLFfOU
zd79BPUkxN0VDjNTTCiL4zsS4NhYLJLb3dQniDUIA4AzM7nhitc24PReeDlGucksNQjLRAFgQAj7
kf0rREj+xBFIaYpr5EYfgI6dcrpoXfjvgxesN/jdjJWCUAKqq1q4sR6nL67tHE5VgLQXEXds1nlh
akbLzMWEZYOKx0vnJbewRGnwpVqidUzKsy1Ioznx6hQwAEhao5+Rp5RrzLIOt3Qr5Vqml0DVL22Z
QzlYOPeHYY9aBeKqU5fCHm/9P2Tsk13NTYE6czsXPJUYcPdVE7va/A7KZTGyevDRQRTlJMUZnNCg
gjDmjYy8lbR1YWY0nYdBS4V17/xYNBesgxzv1QBsR9bIVwIlOOufs1e/dqWDtVCL+yNUTy0Fr0tV
hUOV/cHnB1I2KhBO2+B+vqL3KIfnmwfpAdarAKrd+ceP4tXLi6rAxoha+Gndsm0ekhR1TpVm5yM3
fd6dlgySJOlh1MaCdjfy7O9nnmMe9oywHdBMVao3makVsyU4B3PZc8OSVPMpxvEKnNvx9YxJGoSo
fF0JIowfP/DVWKGSj5Yp1MBiWJLgTn6ul9tIiu/MF4k90mlqGY1EoblBQXn9uMNf3XV7m5e77Tuh
/vj5rsh8edasGW2nm5qNKusk82P7Cm7B42lZC56h8CiabVI3Abfk9o2KmZFWYVhAIPxikBHNuVEx
DdbJFAqIgCqQxHKRpr7Swm7DK5VuOCK2SMlZd0tYBxKIaI1m6DN6ouq5te0avFNWO/T/7LMtbXaa
9rjWaHozgauVpCb3/4KmVGzT4rZnFry+8E7xXCaODXrlVLnp8aOw243tHayVl2Y2wHx1x/07lZgg
foEF58YbxPta6cAlG50WBrjGYGTxUD9FNf+tmXFR7ySQDGzgrVXIn/MOzK+VV5kTmGWGv8VQhLVd
5h0Zzq2Atjz0R+UDIywcSLtlbuxiMxRW2unkE87XQ9htRbUU0KqoZ3vaS0SnmdCIhIbdG52NuKiP
GytZe2ehcIL3YwNslv8lvC0umjIZ8Eugtm3AFUUxZeHuMQVVAzl3ilBA5gy6VhNtWstCtMvd1bds
NDwmkwyiNXKmF8K8L9GaMUb1pTLXArk1ObMSHnCljlTJ3vg/OhlfnHIVbkLhYbTtKlB1LiOynyOf
1+ObfzKdcvP3yvjQ12lPZgy6OAkc00Y8BGi6DglQPrZv9us0QliZabjic2wnb4Nj4KHPfMbQMkQ6
Hk8DmTwz8o12blXPsIyGKDfEmxovZV2432qeC3VlRApcw1XhdLWqU6gL2kDJGSj64h7C2QVJ532X
/ZK1ImggCQHDQMTVa+GBSjhNZIgucvXuObQpiV32exWTbOLp0bTjurdx/XB20MP93A1vEclJgeGE
aAUzooCOfyvvvU3/Sd0KPK2AyQHFwaVgmUVWBWclKohhqWIH1vLRHG2nbD7dB0yTmUbU/mbNy17n
QZ8ZjpsUwKP+jAFV0J3I/JeBZX9pcWafdgysWMP1tKJT9qGf6YA1FmXETKSdArE32QSfstnEbt4a
j4MuoZ9DYLLKQ7gck7jGmgpIVltc04OB7nVFGNYHERN2dZFm0K5XTdGp/JiB74GLcyWzpJgvoaau
WLGpagXwAxiuc/WTHqHpV4n5NxfN9tvg7BA/0B7A++Qu+Kn9/b9BiFUDZ/TOqTMqcpu5GuZyXqe3
2FpiUA27sdwSpjCMwM/Iv0K/TqovjjeXwUYH+3VzqUGzhX4p26sdZZzrXlWwD5CQmgCWVcetSVhS
T97z5ar9NT5PDe7SntewzA4vWgpL9gWcLUbndPizGcbdEg1oaXLVXfpdMy5RwvKl8cywsnxxYqqz
fYP8qX2Rtt+yDoWSU6gZVbPRIvYSzHSWnI6WcN4nidoMmUUVulOyeuxVfk1VBeM+fcvSuK337Oqs
T/r1N+4YKvkJ87nUy5qT3E5NSLoyDT1zrAcPf8AL1GbmMiQRgYMG2LwBlSQLqvpfSWY8wJkuha0A
ncnzUjXxroqlkdJSFFCLqR1B22weBUdYMXLrIublaWxz+k6rR5N4A8LwVJ2spdFaD5uFmVy0OW2D
ROZyxZNqwHZvueMLu5pGUdIEK89zZt1b8Lx2gelTrP9PZWFXYzVkCOWgLXm66OeM+5FXyqw07gaZ
Pp3nXaxkho2Hnl54sF7BO2WTY3KGrGmkCcCXj0lxA+DKdt7k5Vl0QB0OU/PzwL/5ZsvjBlIr6x7s
7TnnZhRhEJOSj186gPFLJA9vxSp8UyCRjxwiGBuqEDmbdfgjYw4VihoMcbeK+slPL+nGnv+EbHby
KjpNUrwQoMwzu2E1vzYS+e3cIMus+xfry6H6Cz8rQN3Sfp3yXaCW242h4I8z+63rEdpbzBhsGiij
1Ad1CPoLEH1MCZkZRJffI+z4m8FPu0oEZhqGi/V7VdUssGww1+HXxsXOj22ttylB88Qb9qUmoGhX
zGleaXgbZI27bZOCKl6Bt02FguXzRzPXdThOBIbQKXBUe1jCGLNndMbE5IMw5pBPeKiJo4XzRwFf
vy8vmzBR2Uv1/4MCD74LjHzXW3bToQLm58blEQp/oxrRAF0fQDPGHLIkGCJP/AEsuXf6jWnPX60r
YO6LJExAs0BEiWdgSwBVcAJeuXMVy1eer+YNxvarXkGbBb6NWCauZd1vu9BYUpZc2aafS1Fhl6Dg
w9EI8DNDtsG9AJ1MOyYarqYwZULv6QHwrR7QEj4NtWAsM7CbU4pw7CQ78RNBgosfq7fb9Py5FHPz
fMiyX8dXZRLfWS6vhIxa70UqJXn1/AQKq59bTMCRj28pM+9t0VBo2nxM8KByIlpwzvI+QIPEFYdc
AXdT2b4igWv2bGGkI5/TR6OCTZZolJrwaxZcaZDNtCCma3JmNbFW0yXJYCC/86+kxdzEdGdM7s7b
sK4ex8GMjpOnlzO+mib//O3MrLDTl7WRA/ctGcRpfR4I5KFhH8g5ZFNv+WaZq5ELPTPo72prJ8KT
Dk5urBzC0l9DgWm+ryk6zWwRQEuNjncd8Bd5dGJX25Y5VH6XeWGvv+O9Kd03/UVmNQxpkBWISWm5
wTnLzcNrQP1qkzHKncLyUZKPfUTAsX8HIXHSeakgIY9LPhOlIlXt/E1rSdWcfgcgqqTWaiwgoa/u
PSgBl3mPxY8Bu375cCrrRC0nyId0IrmFb6w36OaJwLOTlOCMw9a5Rqwcpm7Qaqg1BY3aDyxGSEq6
sDn1TR4YgpwLoFxwkoFB8pdtUz8zN3y7CV1VGenzh1R1vPxu44RfbRaqkkBGDCRJxMu/p6uTVQT0
Q9i9FnaTdRIQOwRPtEvuDsgRlm5tpK+fMbv1bkAojGmrgHcUIPVInwmoQsKZdtWvGEpri5x8BStk
oDaO5QErSO0zD6N9wydOanu1ilsJY+t8iTNJX+8T3X4KPjr4pvkKisb5cZszFQM2WRno+PUWa5tk
L/gKKojJvMeyMUaXy0Wbaz3Di0LVosSqdM0A/ii9rgpRnVdTpoUgISPJMXCjgHcyg/nH89f4ZVO2
kCQefogOfit74hYAa5qU7l7C7gCp725h06Kxtagr3K20R2nd06nDXhKwnIe/zyTMiJRrJmYvd9jT
rbgIhM4PSujjR2Vm9wqHBMbxb9knmGKqbXWvKKbMvI8eRq1r4mi9KYCp+9FN3rY7HRK1zXMqW1wz
VJpWZab13QroqhrfsbRSqRNjGIstQcxheJVuij6BAx5K9w1uRnBUDq2Q1y7qDN8d06SWq10pahP4
5rJsUSMFxi+zF5Jhb6jZU+SEZhx2YG5+FVoLJoTgwRhrVtjmo7tOKqSjGKy7zbW3ccIi2cGq43si
K0Rr0MH+mZITXcjqX/+Vab/tKPfblTZzSRmoJP2U1dyOPoetp0D+8YIfOSRRc9ohbZHyRY3OtxXU
V6U1tjYpmxlXPRdNLY7EyuhyohvNhC847zTp91hxmNz5OSIwZWmbQpJWjpQnkja6lWl7M+skuQ4i
3g5orZOTx/iYK+ZHPq+/wm/8txfuuf6zo9ytlj88MpzgVOkbmSW1F9yno1I96DP8HyqqtuaWVhwp
Gy+ekSanc8YegqImlImmdhksaGZiPNaIngG5r1h2Y4lT/2kAk/gOmkdy/9MwKwsKPkLh/lmnXWrf
RMUJJGY6wx1QzxbAj9ntNfyK0Ot70dOV654h/BFRKqO0Vub59M774ETLOqjSBl9MC7+UYovTWvQr
MKhOTT28C3/7haG0iftTTqjyzQZ1H/GsKwcEvoX0EDZWYHS8ZcEQr6Srtw7hVUj3BatzLtlT5CpL
zAdWE93BotxlSxmF5ADQkBEjT5oRNL0NyYbBzOyC8qtGGsN/86WOU5xqxYVoLlFXpFxhHwLA0dGU
QI7V+BxU7CaowvdfS+0bHNi3wCijMVbt4VE+J8Ss9bkxdqg/n4ps9xN0t52iGVjtZFYlzbJt6/nJ
cf9GVEa4l2BlMgS/T/tv5R24JEN7v0mLuVqeN8Z52aEUPvUp17sgN7nHXzeXYhY2/OIQhZuMPx2B
ydxTnnYgONxeasNHp6OnSiStjZb2+QEoKGwOX73krfw2vNhTj1z87QrP1YBNpJnZoLnOXtmoDD0z
A+WdvlmJHaZvu+BCt2Sm0xZUmdMVcv7jeY0hqKxS3KsIo89tV1O/cq4hTom4NsSaxPznV+cq1O0I
q1nxIicXcKNasHuv1LdihbJsEM5RkSwJTAfDOS7hSad0EUv7ZIK0e647evFln5h+7m7682T+qGia
XHhl0BnCZXusYNgiOs+lnZ0dR/OartQ/lKAFu0Cco1kEVcAxv8qRRt5tGoRZDR/Dlw1+adXCHbrb
BFS0aPqgK47Ccf4uTsw2u1pZd0+GJTYdB963f/X+lRmXiCvfpOZvWPtbjCjSMIf0O8j2vvfh15FW
b1f7yAwm0iErLFPgy0AiqSQjqj/ci+YdweyLqb2XC7Ll42qazBI9oZlvNGky1vhXRX1zG1tBt5U3
xzy47OIqWEwyNlIgVwztCk389SC2ApUIdwvpcZ4gz4l5IIQjB8L46P19n42uzrvTJgkbq0wlfL5x
Dq0sSLz1YAEVgc9OXzDvG/qcHCeJ15vZQXL9zDHEADD5fB5CpEcYzWbwsS7tl/PtN8YIXgDVFWOn
W4keCbDIFM5q/mEznvvJ5N56e1jzs7SIHp9huZTQo46Wiie2E7vHtVT2OCnHyMYWXIcB3efslyoW
Vj+7baEHcn9Rr63rSJ9dbnl3aVCib5nrcbozTNOCyS6biSZXTDpGwHLO1MeJLYjA5z1CEugx42/D
cAVhBPV7oDUIr2XFYf5IqqKe1szSXG+s9R7CqOYMYg8WTaOlBNG7MF29uqaRc1Dh6mRdlQCG6JcD
A05xeFyd9On/6ckqMnLw0N2PnEJ5XsdPjVWFdvWce38BX3haPhAWaYzLaZ9uPLxQn/ly76YOUEqx
Cuh8Z5DO+JdkkPToOZA01Q2IeZNsc4unQR0uVGRnaMpd22LCWuJZL/hkL4tKVXWGv/6u6MabxHja
YUhods24OwEptSKcBDHZX2nsiS6k7oCudcEC0D6NwKHB77z32E+M30u6P538fFTQ1eWV1RN+vkYQ
z8HMV4ZimUXpN4ZVNgES2pdLXTOXL4gGJT/bJyWieK6hkeT4oIBKozRR8vUghA6/54X59XXmhYSj
SfyQ6vZgQqxqAjjWiz7p7GffLtt38dp0wVzt9BeKvh8mfSruW8eWEQLmPdUdHSObLV+wWqcVRm+u
PMBJ8CnD/gbNPYu9e1NpuWSkFd9CN3mN9UmTGm+N/iwrPhsHzeCz3tcwzC26xqqgPgyKm++PBdZc
b80rQ17gVtQUUieMcY0jCDG+bKeCRrSmtsJVeBYZw1SxyOGOgKim9U2k2wyT9TAu62uQIPhXTRct
JmkbIC7PWdK/kQZGD9tqBrSFRkuUi8cI5V5VnQrtePIvSkN1eMVnHf01JXOvM3YIETkdQoKxlgwl
0Ai0Pd9GEiXAR46KC9vxy9j/Qfeo5PLTQ/X35RwpYFll8xijeMqddWqzY7DfYwlWD011RzBLsoxK
p0wnZZQK0cd/DKwqO/wdQkNo6Aq1n7dOQJYIGFAGFBsz9HfalUBMyZ90rqjia8NrOSrJ6u6dKdM+
me8MwezF4o5wS6yjZi90DrlAD7U9h1/HB7Hb+ME1sAms+eOimR3DL1kadIhddIenH5IcPcLQl/QV
FBMsvGeGWN8VTSGHjEpDmG1V66Smc5XCOypfrsm1JmMvi0MhfRG0tDnCrGeG7VM52DGzfQCow2+a
+1PyEVsNbL6Wm0LsTlgYDLSzlGzl5d76S1BK6JSgmVyM25CvKfGWfGm94q8MOW//PLnXK4iTDHog
w995JjLf34whJfQaROjn2aRZh3DZqFVdJcIo2byHeGj82933hhnYEJyQ8537E6YlAULs4A78yuxB
P04m6kuTp4ZA37DGFAo5NLyRFo1aYb6RpPT1NelMGNQRlKRf0MoEcIqiGAWrtQa3P1ojD9HVkuN5
Hz7NzfhpDvbk3HQaj0qcTuAOKfddCi5+9T0tRC3uqPPrAobecm009K0cJEhLiPa6B41SM/9BO0EQ
WIdbqW1hOq98o9VwFKsc9tPvkOOXkG3aniGUecSXaUUsE0Td99NJrnk71F1U5D+VdTetdn0Vj3Ti
jSd73OQrJdgopwep0ROyEPwu50ZJ6y9BHUqQ0PITdlnU+M8VOI0Ym5wSj/NrWBe1CdrZcmXrayHE
GuxrGjYcQU6ho7jCOx3kiutGTCACLFVGDN22N+XSInPYdhDw6eo0FTGJJXOAcmRejkYrG1r8t3/3
eVjwjYa39ik1V8pI7DfMw0+ooJe0clppialr3TvUgxrelTK1WYnQKH2M8OacFDTGQwpnXhWl8H3F
ChvlszADeFdLeUnaiH7VfVj02QrkdOp/DxiVZltABfxG5fQDMmyjtUYwDVWmVtsCkKDl6cCuCcWY
azmCfYiV7dLjtJI1GFohknwNR6b2CzKAL0qVY3BVYVZKycYNbpikfPpDEMbiJpZ0Ie3l5nd6RIR5
r4KuJJ/qEDkg4E2n7IyzQKbSF27Yd8wuj5SXhyGwIgtaVBwebsThxNwwFPqKLSrz6biXBbkN/4mD
OaF4eVWKFOEbsLHGN9IqkI2D8nzzs5q1KUivPpJJ2BSSpmHhmdR1hBaqFlQ6MCkchyzkjrGvb3nz
8Z1RBc02C0HMh2f4kE0XIUDGoW6EcRnkYyeCiQQplCqTfc0Jn0soyVmjuxQu4vekIPDSnw/MC4l8
/2GC0nOOcNt5N9jpG7OPPGAVGBurxZPGJNS5JRYVJQuw9n1jsXZ/2KrC0RG6E+bkMs/VUhrwtOFd
b8kvTipconCoGMf7d7D9nnx7L9iJKGhaLkDeNGyarNezAYqmNiN3lZlUEPf+S3tkpxboK4TTJJWR
PpC9eGXLCKmzAcINSyPHGSJVBDyso0PTmp7IBVlqna6DCK5JCVQDFeFf9ptnzISAdf01P8i+2TGT
LGAXJIjrMsHSIruEiOmOfVNaBgnbEyUO3miZY/7+zEZfB62e5ZRTKCcIignW0EkbuhlB+1KLe8By
YrwnkTFD5Pe+DMsEffJckFLNdHd397oluON2Q0k5+r+/1qBZH5hXOExdtuZFtE8qmurYiMiuShuy
3c/aVza/KqskD6S+Nf395SzdbP4+rfBt6lgfr6LXS0qQHmqwbx2MxMlvP6VZKp2DBfuv5c0S7wL7
HEYBfhVOFXuPK8GzTFBko5VdOj+aY0Az9pkm3KDmdkjVwqiddoo6P/eGmuI75+jphi7yLcHSf1hB
ltuc8psS5OIhrhrjdrRF14OTykye7tdXOJEMrFR4YfdTXWw0bxrsIbMTJ1vWmGH+5HTnUglrbDKq
MGcNX7mI5sJjET0p5JYYRhTxTsvFMeALZB0nwxxESW2CLdYYv5HdCeJx7uTfGZuAwFJo9pMAcpyi
go03lW3R6nkjb5PLMq3UuNN4YyiNR+ztN3QWPpHNVMx79GR0vnvsXLJPQPYvKIuBenL5t+XZjNXE
zlZgnulDpUmofWe1msEvVIdjyAdubZLTxFQIkqz0clPsYFn0sDMIMzOm3Dm340va3b89TlTYXq4U
rF4xbTrq1/kqxry7zvou0CsZN3TOGLCcrLFWSE4PLvls0yRMJTSDkpU18edLr0KpEVz2ZEZKK5gm
0Ijv+pKrb2FgmK3neTTpgcHVnR+pGJFR+RLmY2iSI9w7wUHnBVshvrRJNxrAyVKBTpck94bfgq0e
CY4JTboxJ5Oq7YSHmXKCDCcWtVVpUVbGDn5x2O1DhpyYZ6LIyrb9aR7DkAfTXwfbhqg3osDPTy7o
SxkTeDsMbfDtZjxABbcxKNv1qIbzzMjm2ak5H6aeS3LMmQHsjJ1p4T3BCNQPpzTEKzq1QV47Ikm6
TaGnYoQID9+OBixtRlZR9dSzHnvZDUWuWcms2ZOVLiKEoni0tNAt5M7aIWe3HrbAToN4GuXqN5s4
UJAIHGk+AYesbLI7Xzy3tecbXGBlxKpyUr6U23pYgADE85j8M/TC1KBjL8WDkhKR5FexZJwiob0q
ZCiWUWZZi8OuzA19Q9AhD1XWSwItWhoHuE9MpcgpnSd+IlWLw3fzNAmWk4ReMfBbvrBCGJLe6I7y
oTCEOTAo+iaA+VTrlrKG2+qE3bHPznilI33AZ31ogH1zRiyDKLe/ELjQxPG2TTgnO+KHP+FUmpLI
6noHpgfq/wGzLf8Am4ZTN9zsHQw8N+0d53w3zkK4cRFGwcJb0tQVmRt0IrnXg3yxF1fg9K5/dOdo
njqBeRepmrCZFmGCJCxl1gF9LEaAUsVYRxrGZzuSzCBzvfF5HzfJ0VchVnkCfEee5PG2DUNN1PtP
QxDa+jk7kRzQIQXB7cJqKs54sgZI0vKSYxdhSns8ihYbueN2SCZuuVsQNuuZ8TTyNgtJRlCSweJ6
lNk0/BHTFBeobSoQBVN2UM/8yEa9gcA8lEmypt8i/w4NCwo41h5URxFVStbD5vo5l7ht1XSk9/NQ
abFOBY0seT+SJw0AnqwmpSXdy10HfwL6h+zYGStPsx7z8JiulIPulSex6itDvzUD/n7bt2lvO0oN
IdY/92jk59eec3+Xd+2Y0fXoKjvg9reZw69XKPBAYWVALSDOaqKbGOkVrpDr+fxutZO6MpQ6g6vX
1c6/vreV1mmNU/5xrpSZyT9r10Wk96E2UGuAyAPvzatsHy7Dpty8cVQ1g7kuJkM4CWmrSIX05bVv
4r6MJO2Hd2pa3aYTx84xV1EhSVnZDim1Z5zG7Ooo2n2TfgXRhF/jHSPd/vmg8MUBPMMgKPe+Avyt
x61DoQ+nVMDidCRWSuA3iPBvFRlLku4Y5EV1QlmC1O3Fhtn/rAH0ggP9xRJmPGNtQ+J3Ta51GvyR
SkRQ3ecodpmteH1j1/ny/KZCk17QewcU0FOam/VtUKng4q2rGGm5ZwOiuir7ADWzsSUMsvkBXXGK
EDbkAyuXDFdxUljU+JvEiEDhG3HEf00aogRX7MYFs5MAMFY6eU/JzhhzDi3ftwp1lWmnQ1LwPl0m
QPQX2PRnms3jwnzIVzam1Tpz3VP/4WGYDGshledl51xDT3ijUd2vHa+QreEwFE6cOHNCjYwftemB
7mAko9kGPdXIrPpsD5f+UbkP6W1JjaBkHAfeWSLV+rTq/cVq7vT0tycULGVLbvTvCeW5Yk68Uxfl
n0rKt8cyRyrBI2pJfA58YAg4c1BAYa6ZpbNP1usysh1P5HNQW3+TJP5GcLONtNLlb8V051ZS6doV
zibd3TBjpevQXvbOvcKwAB7A3W04Qm8WupuAM5Xz8uTQv2J5Y5DutDkR2qN6nM1xldfIAXlN8/Rc
QV592U5rCDRR/PaPpKotfiyixhIl8bXwSuJhSGrwdz8jK2c1vhSZb6mF1S9A4id79er5BvQnmHfy
5Ger4i418HNTO3nRzf+prXicJT1O7h1awS9pWJzuOfBxmBb0jSqdzDNnGxr03N2rTf2O/AijI3WO
DtEskrJpAgW7RYTy8QPQMnc8B967k18U8q2KvLs7ehzNQFeTaH2ZeTP+gDls4J2XU3nuEsF4pBBC
DS8Qerp5UP1SNR8owqSYo5sNbdgGe/0WtW0jbK6nv74b2WmnW6j2C3c6Hdx1KFqrgayqhNIW0s1r
8JyvM48cB/2NAXijMNBDq7FdsG48ZGGjIBBuovIdm88cjQvNPKsC+ElxPhROroq36SKQqU84zHTG
8GviDwd1lJhFOmTJOG87c6VugFlHQEeYrnKLDjoMAjclJ9c3VsV2ALtT/Qy37oP0h/S1Vn/5ZaPN
5dHWvE/W0+S+lbDSLtk8gbbLQPIef+PEh7oIuTBH6enpr76ClGJhAzI71XATnjMUpYeRvTNfy51y
acC5jj+vmrDEVneCDA7cYltcyyZnCoOoLmS/5VZanVpGlNwBt9oMA9PbLm0Yxy0crjxC2RKzHnW4
sONlO+sCbKGPVNDC63fFLPlSUYpexcZWoLLhsyoQHod9pGldP/4SDoGGwcBrFMEzi4jrN5WO1wJi
RkSi0ZwOCm3ERwcdPnw6qRTq+SkyBcU8nGzYkL1w3pWZJw9z7qdjEW5VnQ2ilREV7FayHNPP1bc4
4Uwn/VBz3wzK6gITFNPyVzfS4kKUwjIPRhOzz24ILqCW4dUJDj6BeOIekHjnKcA+Fwm/x6St1OG5
XEJplkcJhYVNH7X4CpaNL4W9wbXeWlaEnxK9HeRbI5qRXsfJWppYstQ7GD1X26yCyK6EW7UJ+coN
EnIti9P7M2FKnpCQfqMn1pbX+ga2NVyIMKH9m0Z6qJlnIrsS/f/I9z03H9ZBnlajB3r3o48ZfmFQ
TaLmRn9REpVvjq3E2W+LPtoaB/5USM16KmSPukSTmgsZxl7fugsdLBW6zmopis3G1oZYK7jeP8iX
7ZgPxffZiH7vO2n/FYFfVdNTpYg4XiYXZtd6BfKw4UcdZJD9uuk6AuWN2a1P1FlVb3DOTvMGVlZ2
yg9xhnj3eBiyH1CALcKEpQGzElzIvFGlexllHcNNHB5v3bfcPjXmRNmRkFwF8m3aS42PV1m4zCpV
DRjYODUiRnBrTf8gE2L2VLhWYFl5gmcqYn7zpa5YfBroy3O+NEim5DCLc4FAEP1n3+bZfq9ZVu7i
Dc3aq4FWKl/DuZDH++GzYSxRWL2vJVJQp9zTfhQKRF9y/qcvfAF5017VXUstYENROoJ1xfk3UnbL
fAYdNjulQ9rysH59JHIkX0rbUizavCExSSMdCnpzlGw0JgyV/X8UnBhToX4jFdXG1Qd4F7f3M+ir
ZwXWdHRhbAjaeSIWzeCACOp2eC17Oz+Ky06bswy/Wkrd5jJW7ahSOHAHAiVjXFElEj8w+tGa6e/o
R9LgKB04jvw2uJ4sDvP7+hx1NcM8IFO6hT3T/RgHF7K2WSgRG3CpZ3i4on2pZ8WUzrf+NO6dgQ4H
S2kjlFyQtLaTH0NWlAymfPilYNsnegI3y7YqojG9wF/QDxiiftOOAQIr9P6gk7q2bHPovXkHQqKX
MrJB+Y1gh5B0h4b2kDOKrLnvuvNibtEzutjUMx3M6quE4q9mo4A9RDI35LjTeBEautZxRoF56hic
Vf88yrMiOU4B9yIZiulIMgTSXOXk+Onr1uJ47VaNZ3+2K1DknQPhkzL45Kpm5WsKwB9K4ZL0f7qy
nqehV7Le2QTtn1IgiyS/kS188wLxYfX50II14C2zTEC8X1nexSWqYkgot3j0ejB555QbrCMB1rP3
kEEn2gJjhHfR+cqRLsJeINhdjZGCToRl7medXiR0C3exVyKMKtahzEA1Xg5uubSimu2NjIJA7DUG
igmed1aLTPAjzE3AQEgt4kbVV6LIxiufgS+Pm9v0Z4p248sSRwnpppIOauTHbcaUj2KwHhT/Hf/R
R479+6eGCto6vDqlhEu1MD4/1k12zmfiULcWcv77Nm9i7z2HOmcgb930enILPA67/MsVM4Vgal8z
kK4D3qmsi+KpDZ5BrRPHIpQUwqywpYDEc80SNo9UOUOzJkyFDYm1+rq14f2zsAHW/WHUMJopFCg4
qGUTv+GRHtwhRrgByX8xLg5bNKY3txcXf//g1MCwSJpm65f11Rt8ayGQIOyG68SUPusrk2LtYACN
OMQ6TGGHwxABMXD75idWD9gqtecgHqBxw5RqndrDALgU0bFPVhx4EjtZzX/IyYPa/mmFdZTcRnYP
FxtjpwrlU+Ck5kBy0XPvqm/Cs/Vuq9zViOgWU0kPMsqCx/mDouHNxeSTChdxgbCtWQ3HJ6sMIk7B
K0ez+mPNoNUG0EWvhAOYCPpBXP/p+sgPSMR7WJ621vbl7gzW9H+WmlCA7RswfTBFolaFRKbSsfPn
B+VbZsMZ46yF5vBhzD8W5d2CEC+nd7lYqsaPvSB4JmslO9s3NC7YXxje3gtclQuBk6IzD1LAKbCn
YxPtBixB0wGMUgkPzyIDEkfAP4KhxxfkKCu/RBIxq7kgUQGN8bmoTMIaWqtVhl0PYFC5OSS97d+v
ipujqqh/bu8mGUGmsTkfc0rz0WdJvsOdJDczqlxBT8kz+K82c+tRMvG1NKx8sHFQVfUZATBObpBY
2kvwWmnlB1yGVqW1VueygbNOlW0DKMxJIi+ZOV3vq13NEHUYEv+bRZZ7n9pnGe+0ADAqETteJf0G
kRy/KDGTwFVhJRJiPznYQJ0486YzHr4JlBLaA2U8P3If0SlT2pJqr10MZaDfO6CH35u2UgYqyaYJ
gWWe2Z061eSLxAEaDu5/0AVWfRNtNyc6MR+uelmsxFTrtWBryqnSnXl3BfUmGlRx8DFrWSMZtvbi
a5FW78ptSkMG8LOMe6CPJTTChhtIx7L5T1VmKNaP08xfCmJ8Zz84yJB//HTTNOmjhQ+nOgupX8ga
HoDu+p9WojyKmrF8UGY12OSgE+2kq1cR9wXmbfJMyjdjSR7hHGCa/hmV/NWRcUvjbeS0BouLIkj4
dYaZrsf1ynqomU4Jhg8FY/XD+o+YJfiuKXcnb3ZmZbe8qv/ULR9J/6UqQePYWedqcXbs9fCbav9p
mgW//tazCQF270UtCmFLUvZQQfwJ3weRiA0mTsBHq3dkeUidS7OwkIdxLDnsBwXjQye3FpJ6oDD3
wAGT2DIjyFBGY69+Q73IExPmxT5Wqn8jCLaMVEaaUMqHrYLVzspAnhBaIb6bpwXkfkGI94X3lplD
Xv7Xzmff+ACOR2gYQK1Ryd4RDbEMlKAojpbk5I4KqVFPLIiawQ46c2EQh8sesEK7gaIspTLLd6Jx
9W+BLKI+I+Eu/5eCqKjTjm3W/iVRe01FKd1TG6qFcGApDKT/VdvIJElnwUhYc6OcsIDJx62Yth+V
z+G2cbTRvY9sO97/bXaC91LxQlhv0huXykEsF8YeG8/mgkD8uf2Ws4xZsMxHoZFb+t3tP6L34b6H
duuHZp9F/xG3/vtBbvLtufPrDtgRo8qIrIfHKbBizEYoqGOvfFhiz1EEaTfochm0vsHpQwcJ3PPy
UtDdpNYnZp6GzAS6DzJlZxYPJqjEjL0jTuXnyWF4oBsSkjvOpeXiJ2FtwRc5cD9xJ4hvzJNpJy3q
Tt8L5xBw5uEQfohKqCpU6P39rvRwrxJOtW63CPqSGYmXvvMvE9wKPuqBEY5RxFZuUAjSjfvzOs/t
l0ENbAN4zXLlUzTN+i0wsZLsJCx02sjxO/HaiNeFjdHDISQIm1aYsr62IijL/6YEmUB6IYOs2RgP
cy53I7ScgWV0PZxxVXpvd1ULqSfJiGOadszVh+QPLv40mzkdMSo5gXfVPB8zD2lttUxBZKFfC7Ug
f5eofkiIGTkequWrNA/tNp5wRy3WNXKlhzp6mANSO+OWUigA3FVdumBcXpCHX5h2VJbXC1ypbvJK
Wr7hLTjLmSKNcyOok/HLdhvWlyb5LTTOXWq/vKoagEdnmWwcJ9LXVIiheKZIoZHqgY/kTt6039s+
GLRQHV1mdDCJoPzeXF66ZjIYABP9z9XIEya69DnCet+LErbRk94B9gt8Q58gXSWG2KtXsnZ+Lsro
C1bbpm7rbmosfRe1ik3w9AAQFnGjIcA80E5VvqufTcNZjEGKtspFNJY1Mn4MELm0vT88uwqNvr82
nfYJN+y78VaWIaNK7qO06aT+MF5b5n16heiruXoODs+mvTJzgshMq7ektTVg35z5YG3xPCXOdUox
JCGSS2owKE7Oiw8HmepCpOYxeUC7TknR726HqjGajWG4fw3VLZayeo8iA3YYOeCFCFuW9ao7+zL1
jureFmXD7nBdtS8t3TUhunGDQp0c7zQ8IG9P9LANbPMtXiJVBHzBwm27KGPtkev7x+T9aO98xs50
oyfkAossUvp9GZnIqGZntNO2AByWILwKScSIlPmvr0W1xjx6JI2Ht3EQY6UqglAsOiknX40U02ZU
/+vUJdT13ldOK8DY6jsm3Y6h9jqBErGoFpBlM6SIJfoucIsNJDf/3WVD8QX+s0yt66IhZs8KBm6z
O6wJ/HxpFfJqkbCUj1xDcWnKPsOlXEguNAFa6zcctmNA1rV2J1FCZ9aZXrU1dyOVStCiGYzURq68
yuhZR4uIRWEp8vIfOKWIGU/7BMot6YV1aM/7+Qu0aQujcXOnqXJFx03lb1a2cC8qfLt0p0imotEa
ILtP9LxsTyt2etLxM5iTEXSLDiRxrK0d7o0TtM7T4zN7NPrubGTxNsNpDHGTr24Xk06Zw6D510wZ
OhvPNQim9fD1fEva7gdpbVnp6s2s1CaXMl6nXmOlG53O4Q/ahIWjN8wa5Tn5sEkndp30tvovssAK
I1BHOtDtUoQ/Eix2Tg/M4rkVoDCaVZHLODzP1WRbNNDbeyNL8IHxhflSlanxZf8kiOWlbAdnveST
nHcbwZ5dkww9S4jXAo7urY8nNKJJ1iUoj4NvZbIoo/Lgoh5DaO80ypeL0wDZA8BVGfNVeu5tU6vk
LYn5Mtr3KCJFMFE685AKEWuzMxdiqDJoSTilEKOf1j/H0MaOwYGHtzotN7g1S2Lg5W+AuE7DP3xu
yPhQtk1cJT2Y3FcU6TtHVz9cp6zqAJTic6pMq9QrI9JcQyqEZ57/1X36jcfmZSLTK1xp9s1oCX3L
XPirQSSREnAig34eEoYC96TIlAzwKAjHx0k0IlIDVoT0ZXPHi8jwj93VtSdf4KxnWTDsOz3SpVxu
wxhZsVfOUQNx7CIQuhRTTRQ8pDNt1svEJL9slKoHrzl57zkygAbVEaCU4ApwXXzsDttk2jpnCfgc
xtNX13apGQideVTf1CT9Wu+0o0CNJPDUdEOfqnWWlk4QfhMR2TbEJIDFwQgD1tmv2+vuvt6NKb82
HB8q52opzbyhpdqe7wDm8hxQGNlUfCX6LM7X7B/bJ93lflZbywaXzyHuCOdg8cosrqN5MGnb44Ea
Rjly/UFb/9bWgKTAwosID853uGYiYIH00ms3WwqH+tYnPRsRRkgR/G7nIIVTATwW1FDPdJ6JUSoU
/Ku/1K8YWzeNUHNmVy+Z/mUujOJ58L0/dOEgHr1t6kprBF60i8V6fu5hn1ump1EG1a7LI2Q4Ln3x
xQyNnWoicJzYHOeSyjc7pkm5xF3QOVr4UKZgHygEmkc7fySS+VvwA5p/2r5z2qvxi5uTBjDb8dSp
tGn0wtT3XKik1W0tDlBmmpWK3OyFqZsw4wAxsEL5bh+LdcFJzlH9+kRPgSaYd1ll3woRFlGhcixN
id+4SG19BjlsmMGMdsdAfhFWGeRCrNM6nLnLC8pdsboAEWCqn6/CRUYL2bZT300C/O5lDcevNo0K
LqGj5xt2VN7lpU5oAdLOJJod+846mkrsYaXp8Rq9gRrWptIVEVC/o7JzYc/H9BnuKp2iPHyGbg5G
wqN+hb5r732a1b85B3+m+Plrtp94jqEugjGbHMJVDnNUaQSU/b8bVmy5oAKZb/ZRbWAqQQyw8ggc
83iOByIg/y3/AncmeutCySEf+ZyDXjn5paGrj0VGhm6sRagaLQE+5gTI0jO9sfT2p8WVWj8DxZX+
pyWxxoXbJKNT3uUKaok03nnk2RtnO0FyvDFRRO40H/hjn/HiTtpBLFtV5wB//ZSdzja2NhE0EX/k
hVOvThULkkw4uBz6onVTQ9tj4hri23lvQ6pmn0kQkzifM0DaHBg2fVI9dNtTCgaPltIRQkMAh/DT
DKpppgxYeEBrmfd/PzYUOnnoEZP+1GK6kHReVD/oMS9hT1wEIgD87APqquVNzIRP66cBfOMbqmlj
DB3tyqil/Yqy0zVoJTddTyBiMX8/7Tvg3RcES8WRxA1CxIot53frQ4ZicnRTBkWVCMwf5zJz/gF3
8VY9tbTRdBYMuFTd+iFs1hdutPzuzDlAKhT3G05d18gqN4BDO1VtRGRLGcfTnE4JLS1Q7BZN/WfG
dP/HGdAVocDEzCJm0Qx0u96aCWnUOmYvHDmzUCisLLOPfO8gtrAE2M3Sq8DXeF5AClmsFTyznhlk
dLeQAw3aMyNLDx5mirxfxro/lgzihkadirD+onalYpH7DxunXODl6KaHv8F0n7v7EHD8cE9vsuYA
7Izr1qvfFE4cM2u6kyAUGUmlUbd2m4nK6YMtg+SuX0TY+cQCMdtjymfIPk4S0LNZltL+0BXHjReW
Uu7i/5Yn14qbYsZG/aXa9u83Z33UPcQJ2g0NSWWcGGSINfPiOztICo2EpmnwZx2b2rNPZwWx0dIg
LWuLB0TSHQEASVMnE6aPKrrmOuqmSn9hksgxTx9zIT/kgh4ZsKj2PvAM5BXDUuq/ZE3n7MM4UHvq
3Vqtj2itfhTzKCr3nR+GglWa8GHY0igwU6sI3WoEIGmjFWzRFIMrISorjGWLGLyTLQRb51X+JJgj
vGZkmb+XL8oBIenHS26W475sJ2RFoKuJWusVzYNHyZ5zZ3Ckji33lYKyKnx04/CiVeoNf036PP4Q
6uvD/g2ft+fANVaTmBQskrorCpPYImWDi8dW4tBct6IRGkE/lpTSb186FZzg6TcIibOzNOGkn5GZ
b/93TNK6ovrYnGO7DQd/6WKBSNiOmR9m+XgnBElBdXJe0l/dq8KgoYzpmUXq5e2fC0YsLs4BTM3W
JqiODtVs9IzZprwRHsGgiINc3SEIeXmdGRqilt6Ca0SP96oKly932xrmlHUZlp+2+tfAS5as+WTL
nR1+LIRV+S7GrDlaTml8JKBxmtYFyZCLtKJPr6GKY45SImuo1xeYeyk5W/9hS0O22ShFREKcY/I0
tvUNTDEZkufzgOCXcbuZZ9wGOoQgPMlqKJ4nQJeYZLTIqHgKqsU3yDmb7U6T9leAjVbGs1roKr+4
SelfzzJlda7z426CBeuAzGg39JZuvpTi5gIKld7/dC9c6TL1JM0K3jU+GorH9DGrjeHEYUL6XzI8
drAId/eaQoLVQT1PVJ2u+eCzXIv+Gs6JSIfQbaj+cmV8Mg+LSiM6ImD3/FtjQZLvUxM8u4jODeTr
F1pUWwsZfIy7JUIAIiqLOTKtWt3MhvTUylZUy+4q9cd+3u7f19bRX8+YMGwB2O4q5TkpzziNrZuJ
JQ0FKdgh4x5XcdJfaa4mvmELfzfjWUScG+w/WItNLlEthQJvCeKG5nas/4VNvrUVokEZXDghMHN/
9xep8z8jZTXHVb2QrkGIzdhOIx4pIBkiz8OOVe8/OzmNkREbjkw1clplRWaeqBo9gDZ/LK8wWAUJ
3YlZuTAJVXfhBXqpx0hvr2t2vowIVx9uJ2aX2gaWcgvcnq3eE2wl59dRl57SAAUDTDD3XJLKk+1e
G3CW6kLsbLtpyp0wOEYsJGQglzw1lXXkqYZxVab/hyB6EwgAwaYJalS8LgzAFjBhXpL8mBPKHe1+
Hbf8k3NnnqO9WTxV2z3mbekGw2sLsgYZQZc4EHQRL9rB2KcC6B9pB+PotJa0WdSG/dRbFJppkqPy
sBxS8e1uXrW5Kh4fLsDfZSsMKtwAbJN7k/lNcu2/IjdLGQTM0WtPutYdICKSXl+Iy4wxOXJgRU9B
XJx2aVVHodGqe2J1Cx5TXWGmM/HN3vG/gm4god2BYIIsBkYFkI5V7c6WCBAgctI1KOywQ+rK8bdA
rKKFRNNYeFfCK7EAiRTJhEmhr9ZAAceMboBFri6Uf3pK0yjj0exzX089dkU+fIz8SsyWUuif5EVr
h1gHuXHrnbZlPMue5j0PAlj8HN9wKykdnEb95PP8mM0cpb6yfXIb1tbPNK63jfZBh0/ykJ8Ia59E
NbwDhcGwQJ1yha/U5jrjElpBhkJFvbCL6Gd4h0I81bzirP/gu6Mc9MugD0RczGUPk/TbyU8RT4JQ
olYgS+a3iZIY93wMmByrh8LlAp7FUR1jvPMlSF8uGssrG7i/w8OYSZLBRhEPU32tMrhOncSQS/dr
kIoyBNNx/T1/wDm0CwnACNyy0/fT35THHlpAG+QfZyWgp/p/3EVVz+Mw6Kd8X/kGW5iYjwOEBlbP
so2wkVFpoen8AfpGmHn9znmflE9hbVD2vNctl1Cs4zJvfmRYrzgdQNcHHnO5pxpVJMMbSlkkFax7
7g4myBB94b6cp4u+p8lSBxhw8wr7AFvYijJJzI/tNFPh88WkSoS3eTaqJROE+ndOGy30JX63OeK8
6g4Ne9VJI1gKlAntdwGf9i5IS4vzZSHR3O8jPUO4Ntz41D+IAGdhwYeF3oOmzUA+qHv7xkW0bKMe
q/RQJA2kGBQtciIdd3nlaX7hW/FLPkrp635oCRFHblK0QItie56uW7IyIJvhb9bJeVZOG98+CukI
atbjHIEGmnW5lzMW7P6eIoC2Zr8UuWZaZwcb4pT0HtMyGDs07VgYCQZk3X4gWU3gg08KXC+VMOlr
NEnhy1R/1E4rC388m0Zt6dxEPkVRXyL05Dff7KDV4wm07Ma0AGYnCx0NB/NyaXRv7w2b0xgSP69z
Q4CmPexN3J18WSpuOg1OL2l44pHdPGeUuZKWlFlbFZp3h78WlDsTD85d9iy4lUsRghWYvkVmQsGR
/9z4oOoM2d0LYFdoosX8oOwDt3kPpCmVQEQ4njvf3+jE006/QVbgT0/PisjcXqq1wqeN+AIzBr2f
VxzfYwK8g7I560JxA4+0beMpk/5RM7RY8ZodXC//P+TsI5Upss+tNgowSOdf93M6czmErAYWHNrP
43ArKuqgtrHSrRzOfcflDgCWcaaHhkQWslO9C+cc6Ol95pqulHbsLz9E57XM5C0mGUySiCcBScNN
q5tvErw8G60nU5cL/bjF9QhULRPuQ+dGgEUKFS7ONgG6vW7Pa3mfqNEBEF4oBhRxwah7jlD7cHms
NRR8wP03y9Dj//+u8RaqEvCDIvo9e3xAb56TW/dvIRJOR0UTeLsMrkAy+MAIVe1vUxxsSq6ctDtt
8xBbCfqMWtc46RKZfHPD7baJZBzxmM6fUUPqmiSalexA2Iybzebohy+XZHTc4D0o1dPrf4IIWUfK
8tPKXSj8W0LRsZd1TRh0wigmVkviNYx7MXwoAyLr+m0H/4/2b++5TRma34UaCkKDSOhYoE87IAAA
0RUv+wqBlJts2OcvmSRKgdbwPpTX9dtxy06d6dIX2UV19otPPuNE5rTw/O9ViPgryZVxZ1gFMkjR
UCYv4SWj9X47JbBJrsuPl9ufI0tWSwNvgNB00hY4eIM8GVPGNDSwT5WFycIzzqlrjeEl1RaCawTG
RN4jLQzXTzNiaJYjSKklBO2hNbGQQbgJ3JKa1BXl4w0m2Izc39uJOnwmnA/iXTr/aO9a5NtWqYgG
OYTukrsdJHA91R7b9noeyqnFUiInz0ZhiJFgRZB35DXRJmw/xq1weE5zLtoIJUrZE8R+pZs1Ea9S
c+i5JIHLvVgQ4VXbCKM7b3mX88DN+uMXap1V4LtuecvUu4FYVdW2FVjAnkd7Cte+Jav0ShG6q31c
G1xRh2nBqGpUdbuYMPRm/PjQum/5TB3E6KM9fOlTScVtywZ2aYKVvPnZdUKquSMyNrGnJeE9YMg7
ChwJih2D4hbFkY6DpxNoFGhgcb5QO94WTVnuXiSQj04MeJRWemjGWUQ7BcWWu5OMy2nI2SepYtqP
rbDb/DkZDoLu0D7tgV9E+aOlGIwt0Tbhad+OY2eJpq9UmgRZiuxCHEC9Xw+pM9jbnVfTa8IcNTC1
Za+Qxf00xLGAVx3XuoG4vMRPAfcm0Tidu17/7Yr7m6PD6vUkcRtBCpnuMsjwAEk85y/66M1cvNG4
d3dcV9nGzJu5/z7X0/Oo658YzzRSWjl57x/4znycPqUQzcoQE8w66tQp7PIaTNRQCFq8YyDva5e+
xWLXN4ENqA3/0c615NdIRhfZRl79vjlesc1nzBc1X5pUDOewEOFNRae6MoPcU85LGwZoUkog+h6N
exurbb7U2QMY/1UzzYt9csYjlG5kE8VJwk/ywTNjig2wbU6Z+RHUK0IsDPzVT1ld8t+R5yVV3jXa
CbClovrqO2Z72mAfMGiwe+JXFoZJwejfIT5Fkpx99werHdkVK4tAcwtD8I098g5w8JyDBQeJda15
GCwcg9jbzqTlf8uBZtVMxlLy10bwlZnBywmQG7thJTT1HBtKSgWg+nJ4h2QUKI3m0lg63nlsRkOf
UHUmEinpdx/iTzoac7uYNS+h+zZKEQ9+bN8xHvcSNC9g+oGlpX34keZ30eYEynL5bbZ08Chf/VQ9
8oEU3RhwGQOtQBQ9Xkq/CVsbZsycgzKfI8QXsG4WfufOXRnlkmWffJKGi5xshMbunYF5Ec4MPCqK
wLnQbqrhAsaYCFgVcqUvVE9Se9NZnxurzteC7QvdaibD6dFHsO4ELAWw7434dDDepPVnmqWNkscv
yKv1vpbfYOBxGS6150Rb3e8Fy2RALzo5Kvu/nWlr+NkdxMrCUYNBIL6VsOsNu822hQnT5uKQeyEE
+xLAqII1f8xlf37HtCgkRC9XzWlEoHIflPi4J69YvtXTdH9n5Tfvwtd3zaRastrvAxnIq32UmJfn
1pI+sZ+k4vw0avIzSN/WgPwoEHg1RPJ7iGv2/XrC5mzHyr5f4lOLisdovU4eYntZU6l91xk12jG3
SrzeuOC7AglAC/bLaR2lUBY+nY3OqB+fuwYJnPyGhejm6CxEzX7sMOs4PbBB9VLxYQdbrVb53PrF
PmxASDhMmT2eJ2QBcaD2XuQ/3SErADfIYZ2carf8RFlOr8S/U9TJ+K1OKJNCd99/Cq//LZoKEb/I
zsyw3rdeykqEtFJHty32P6hZWtoN2Cggqm8APQTbJp4e9JZefkM/UI6am0+Cptr+b8u2f6ZLiX32
DZUciFVthxfmkyBK6cGaHBzaJtIU4xy/4+jxkzv6Dr6LYFJKBz9WCpvsholnudS97EPg0xJU0/Kb
KKf3hBXOhUdkhfKEp/9qP1e4r9sKW1nP5K933pQi77al8/KTIrC/aTmf5qRk44H8oeNn6tbERE+g
6uQwiW4DHiYERYul2eJeb33I0g64SeNzsOfMIgF8/g+MpYNJ31Z0fhTJ641nFw9UJvawJ+0TinRS
UADJTuGDhvm18gfJOEcPbjbQOd+aTqPPXJBrKb81ydidKzt4qZCa/4QDueg+IRzpYzk+A16gl8Q/
Wn4LUVqk03O7SJNf19CarxVKzILcxkO91rUwuN7u+U08VTp/oOPnD3AA5iBVlVDGW+Sh/6mdK7//
2vwHfv3nv2eja+HIB3towLaGIjEOfGanqy3v+svNTn9JT6A8VAxJJLkYNAZHGXpF1YG4FyUOkPcb
4T3WSvz3++1LmIw+MKm2/ZsAsSL/a+VPiTnUr/6awBLyIxG3f34c/lIEVb0vgNutEMUKRND9a1XT
bRAq3gtHRvRolnTzVBjisHEdC41bCZ3snYIBuNS2ImQ4mGjYOILwkN3jKmODkkohfxk+oWdZOZor
m4J+dbun78uEzr5PkMZxlKhFkLb0CbXl+TQTq6S0QMuScoZleaoRdCxzWDxL8yWSvTvX9SpquEFG
jyloG6rZ03dLhceQEl6xP3R5L0x/qGaTAuVAU4+oyefeQSwoYagm+7cck3zSRpbGkPzbGwVuy8o1
XqBpW+9JQKy4OStBf8pevu4cOUA3buexWcd+CvI6+FTf4dbH6BHt75rzEx/5iHcQfRnqxMIpcrt/
yVb/955GQ2xNhvDtIR0Ebx5Q1wYrrtykYBm4acV+RclpnyjPb2LGgUWg1rxJqfsQkFV/Tw0kZ2th
O0PnOB2mwU934Df+JF1ELABXlW05bcfPvpB5bZFfXFKI36YDOiGB6d3wErnncniFMQtxN5zcIR3j
rpowMGTWYHWwEcc9N/wbZ2Du7etSfk9BRQ1hj3K5K7Hn2jRuJqfWUYaVqwlNSX5yIBHJqiUsE/Wx
Y75x58ltQAU+jjWgyv0fSGNxAoCUSSmKw1BVAPjbWzxW6tegHCrIdQLpt1nBAQT/KQL+lQ/RYCG9
yo8ZEQ2ZZ3LyG8uHLyLda+bIE12hhT3HBPBuvgT1tlcocWtsNwQI/cV7uzlCVxXDo2MWb8gjcj6p
9RVGdNl1w3qbvkyBPa5fUDN7idWz7stmN36H9143RhQjrk4SMKPeDlyqoniIwRmv5iXkyVpmPkG3
dRQC+rnLIKzi8LDr3JxhJ/1tQdBDonZk+llbqpLlpT1oi5Y1841tOuuf2ZWLIk5Y4NVxToYsGhsx
BDOItALtyd9BFV9FSR/A6oE7C1e/n3N/TZ6TybKht5zIG4PeFdERPDOl7s+J1Upf2lJURRx33l+T
AsF1bXINLMdzJ1T+F0JG2Xn4wkD+bic6UkYGykQhwU2pfjNk/9wDdZK9IO/9Axl2qgauIlj6K4Xj
exEthnvEJfDdu1IWS+kja6PxL5sF3+NIz7tMYuNg3gBJ7FLWYhjoWbEhMigaY45Kn6FiWHxzFjDV
Nxscqb20kzvT6nkSTKbLJHrOwK3hcC72rQmZslaXNHhEDulfzl1ieg7dDf6YEtyWnw98f/1eYesk
wT7GmAq7iDClU9kngtNuxEo49l3VP1nCJlo0sIitpdrAJVzKvuJ9wARI8ZF5U2rD1SyaNtlNUi0Z
wf+US9GyFbaPS7WW8Rt4VOFhnxQdwpqpXOpIEU/+bOlbv1as5ANn0Q/NmJ5cbaIpwFJRjBbXo3Jr
eQ0tM7Uk3oYSedZWx3iFW6n4v9fi7uQT9c3PeEyLN23x/G26DVK5B0yEqUB+D/Ia6KXZcxG1MJO+
1HD3t/V5d3Ra0/L69mududf1TDAWPJJ4UqiJIo1rYk/sBApbhmSQZY7YA4WYeVRm2y86jLh6I/66
OejwoBtQmx/FyA+9hDsvpEaYUg8tsKUy75GW/HYhJdzjLmml9bFb9/0AM5eiYERP3NyxhGGBxuUM
QdA0oQUmGrc0ag3IyY687PEJal9P6b1uQAC5c3r2T9NcIyk2UGsKspKoNR+IEsC92Wrw2wPb6hrv
AfKbc9mVG47Z0r81YZN/tcW1YvbqPMlLtg1pzBzIBTTbswHr5yVD9zNbHBXgV8DTvC1hHB5KMw3M
ThO4QukGPpNHdQ0DUO89d5chAjlVj/ZY2xegVjelJaED2nSykg/dttrlYq2U+Rq0E9B4PuKuwf6P
7T6qNCsC+j7QwHSzmUxVdJRwSuACDEgqd6YtpDHsGks4unEU1cXD3cnZgT/TevZeB+vJyHYw3fiZ
iDOiuAgg+cVK7snHvkqd6LjJz1grevAP+4xxO7IQR2aqaCCTraeYRAQClvaqhxeBczhx/LuyaG9H
Av+CW0R4H/++6ssGP+f1/bkZmMFk05LROAcLTMvxDH74JzQ4q+ii2OgLaDaV1Lp4JexfyYh3O4am
LVaP0oDT073rfHbeJaLRc5BDxmt4jrLHkcVnCnWFVoWRQLB5QWPsk41v/uwj2JEPEUE9aVNrxSyD
+NkiRQEhpeTnlVHsrYrFZ2Ta3DkevqS7jzJX0dUn4EXWvmqk3rXOQV0x4OkIZj+9f7Q5if6mZPZn
UJvGFrKdwNykrNnill9KcCVEqQmvHZym2GuoiOyFIS01Z790WFUgBKbLK3ZgHN9GpddqFq3iL132
gdnJnAuJiEFT5EsSXacacrs+J8kZAqgKGxh2yVHQDvIfpN3A0A9yt2cF+58o+1HHiCA4vAiC47A/
NWdk9oFzmeHuh7rC5l+TwQsIdkHOSl6Tvi8KEjTvqDgY20Ga+W7f5cMuQZ0+o8OTODEJnM8v0+KT
5XufAAtxRci94iXB1YCDveUOUreDTSbxRuL656rQ8WWfBWO81CPV/4yS0mm4h+leyalQRadfYsOX
xHPOKpcTM5Q45DNRSKfQLkD9QclKaEOmfrhWQWamB3SJCBTA8AwzdLPMJYKoQ0lNlhpcTJyPIHpj
zpS8WdH/jJySAd4tumpPD2lFX1rGF04YqDL58+fuzkwu79ndS9nC8I2hzW4t6YVBHM6pvLpkGMHx
Qm7Xs7obcGDpz83jEU2X4yv7SYhaqMuQdR0xP0u8p3VUt/lCFci0i7UhcUT6lEhyFNAdM9cViNgJ
L5Yi0H7AZHYsyvOgMCJukFYFjKTkzCLNaNQoImUqNaCC9oYvtGgvmOk/4/3B5JBEjSDozYCz04FZ
x6WLE01pkxqbdwBAxATl9Xep0WqJmI0ajsn9hMAYzqrb2airZAenZE4h/nY+Xt3+GECfD5eaHPo/
FtvXSyvtNIMT1wVhK4m/5kSCMfVeioOqGuqoGljcFjgw79qHelfzBTUnKUeBtg+hUu5niUw/Wt+q
lLrg1DknfW38RfyGVLC3KKV3eg6YVGLA+0kx+a+fWVVADNFOD0crMfpfa8tJjHPuHQ7LURcOXGRV
7NCfqSaDpFgBwFH365KfyQGroqL8/+bvAzD2x5k3VRinPKbM0cQIr38YAaxdhI9a7bVOSGcUToQh
MbPljMKlLB1aH9A3ZKiQpLG1Gw1C5XHLQKWDi4+/TOkWQ6jU1i78QN5KQ1wGjvYxHFLxSj11VJYM
Q71rMlqGOifvF7saDakwo0jYogsNjgh+daBzl+shKzpXa4oWS2aKnOCoZoXgWE7wFyC/czsXzfTK
6Q5Q/1OHX1OunW/Yaud0F55ZwrQ8+6DcD33+TetmUGZbqOZS5p+ukbqX4mqVjmyeM8Vw9HM/j47y
F3wI9495udiVlQL7MEuyWTROVYz1Co80dx+WBV/bzLCH2c1SGbC9bVQB8s8q2iqlo5/dugv903pt
LjTifVDKFQJGRTlq+F21po1K+IoqOx+iIQowOaecPyTLEFHwDMU8fbMw2WOSnMXWaZkn9ghgmTnA
sUw4zK9UloIb1ZwPB5msZEscp6MW7DCI0AIZ8osNeaqD5lCq07ycRp6GRfY07hVlx82GgHrW3KD5
fxccU5KHekX6kaY9LXSdMrNOhCYpg/tHv5YH2YoaN43r4+iKqaoA5wlROFHopIg/ZIXlqzjEyX17
sVlnfvu6+dSF5tYUAZO3BteXGGUL3AM4rYzUhJt1RueOlZqb6R02g4xqzL0KQ0n7RyEtKJ1fIun3
x/SrtKROBWraJDiaG4wjUn4KKhbraElU7zBOCoJSyg6j0x26iF4JmCh8LbO/aKXYnfHQSqmqMqTs
5bWv5WYMuqdDphRjGQ0Tor/Gt/3CQ2hm6pfBMkmAvfYGOiFnb67UvYj2DbSqi/G7mqzSJ6SGSTK9
o56NBPvwScD743R+fpxdLjuCOymCqbqNeyHoGzg5EbgHgOLQN+9Y2YUr6r0lKOqAu1sfwVoTZlZ5
+5BbLw33nZ0mjiooVC/VKy19ACzpvM0d4Ev2WVaXNAHvj8+FNDZ6nyPaM/32rYC0j12ag2QQOX+M
KEUmZ7rR2iXRM/28HzJLG4ot0Fy8b+wH4Wwb/dN8ugHwwDeNce+qR5vgQmuzjoH8CTC4HkOkGIHT
9RypCCqzVt6Kbcptv+rJQ4g8EuIX/aLn5uABN3dzYgqZ751Ru9rzzGTxQRN9Kvj/zJLP7dBeVi8m
9/IZN3iVyTRhTJPcmU45+WaeUZhds9q2+ZeR+NJYJen4FtN5Kyg0MNSRRbmUBYUuyYfy9dk3XC43
dBLu6dU2jZFltfAjAgAF9dXWTkbEO1oMfgyNHHlYWiCkSgWCKEkjyLlwOghuG/8jV31WA2Dg8z8w
x0XKbtX+2jnUHlLSdHIl8o7gF9dGTdNvtRAqn3+OpKjldefH7O6+MO5GJ5mdmgPuTiVMMRnAZY1B
tM9CQMPC2ER2sgyv7PLWrP9TKJywK8Es5EnsMOIjniyaXcCG93hfcZj0IU2QzR/Ernu/O1iInFra
3h++b93m+WACkqEhr6Tlr2psIf0DgC6nKOyMVqtA0Dbxh1Cp/i6Qs+ixofKRLLMoyfBVh5jy5Zzw
+c0HglUBYkQQO7TKM1OQ9eTILQ0cFKH8DTtassY73q5SArSIgBMMaMpd/MvYegBgM8GyBpcQj98+
IwxM4U9DnJp3knueMsnENTk59s3utWV7GBvdFE9h5Hlz3ZZWIsvjFrvcu2p03a+uMseRDHgEYXyy
o4msMq58FdpikOkYie9gl/9j0eWGt38nvzfekY3XO04lgxLnpD3YMntLDXG2HKftaGRAOQvbJvDQ
3+r76b2xlgmtrMlbsROQoj7bUjpAQLr/LARQ3ohWSefZDiGkY4qDKGfAptkefpnK8/NLXa33gf3b
rSsv9iD4xxT5/e+swt5S9I2guKfjnh4j1VL2wsz1iGILIqr5ky2RVNjBMXjokT0etmxFwPVJDauZ
dNa0D1/Rl05L2C3NwtSddwuWyNHqPLjqg2zatc1m+IBNL0zWEnk26vlXKQ26k/Za6CL6qYKrDQHC
xrjXBLYRSU3GhN0pAjXj4NdOgTv0krIc7eBSWzua8Yy4rNvMcWPkivEcGZUSZ9Sgevpu7vKAOgx+
4oqwZRLXFPJOHULZmEopJgeoU6oir9iCvP7Ni1vkMP9IF4oy9ADhtmoDaDsYwRUfa3ANbbLOD03u
cb5/naYoO+zvG1+pwJEaM/ws/t9epZ6KQOFYtir6zvmTgJStJPEoYu+VwWeCLcUzLlaK4hZBczZY
KqJa3BoBpX+SbPlKhxBOpLusoY8Jh/oUETtyGSUBuCKL1x2lodPkB2FYI5YigVMMfoeDdgqQ3Jg6
E72ifLMKpVAVDvZNvuMUkH5xFEu5Zct4oQ1NszjCechtgstmwVFB/G2uZagkEEknTLEnzjqW3JrX
voA/WCjrxvG3InSWaZMztDPJ3lcH70NB1GZ8hlSiJHscJ0e5sOl5Uu9ilUKg9evXp1xoHRkOjXZV
+rGUz35vokx9HqGYSxFb5/0qynsZZip+r7mPp8DklBjVRYG+dAuSGOLtLDzaSsPnIJGsUZ8Djnyu
1ikMYQ4ivKDW69lyebJlEmg6jwpAhY3xv6p4oYni0qZMR6yp/2E1YlH6OUV4ttDkscDg2NOCqaY6
8HCy7iYKnUUxc24cQuX+aXEDDn83XTXEvpM3/h7+arraPqwphKIJ1RtF5xPsSTV4o8r3JhpyClDT
AiksxzMgR2ZLcLhhzOCKLVGg70IPoccb9jEKeXcsvhb4QWMsgCiIe6pyR0ssEJPmOD29AYtIpOG5
yUH0RLhmrDTCsje95t00QRqqjNGtJp5C+0jcw6qyt33Qr8OBMcAPRApmtdKswiMizxHUYXiR8VN2
wrobXV/3t6gCMfSJIOqPcddy+kH7foVUxZIFScwBneI9GpqOSTTqtJG/HDuFTJ/Rdt0fZQtSkGEQ
RWXY8/dHxgAff+b9o1MVfl25xjvXh/GNFvKaBvDQZT6Hd8KS0WIg9HZy/AJz1KKOAUNi0M8hlg2i
I639u5kMEN290dN7Xg+4bTleZoKYIOv+stSaoVtbqQjUeO+Mv6X5b4ERRupxBy0cL4LXcQ9U5RN+
Ol1ZOzRt+mB2Y8ImmfOOcWB6AOCc5LmSyUY/vlsTkE8s5z7u24tAD9pn5TCBaEXYNO9GJ4uKdcNp
i7CDJc+mezh6KGZSwniP1q5j6f2sW4N9IwESPrzYc45TUg0b0gqegfb8kRXaV3iqHS9tJWXu8KEh
DAoa7ZAWT7hsoZj7azxrWnhXPVpUq7RPNpgGRvmCFhqd1PKTfWKeiSzhJRO5Ob/bJfsc1HR8rxlm
toxzhJN49E/h0n7QRk+p2VWFzlhrF5tbSWL+Fva0kyzJ3VUtFMJB5LAoXbMs89jjKpNf8kvw+yuN
zPqz4xQwta4lAjWcrLkXiAg3KHmkCzXJc6gOmRle+AynhxNBL10ZhDdTMqBUedmarm+1iSv5zopV
UPgiCjNWsRiVizfPC1anvQyFG8rdvDtN61+2fOEoMyH3m26vDKg6wxxGNteh5AaIE45svxxGUCeQ
mIh/qNzUJWT4FRSV61ODiWkPLWQ3WehmBHalcePE+dMTnmUyZxlTXU3hdS17q7lEi42NlwIZXnhg
JzFBg0aWKoJhKzJUtcJh10ZbE7A2lJHXumy3k4D1N90JdDOWTHwU24JS9Ixlr+Sl0l2G/ZiBHE+X
cpsfZMPqhgpLbgEbqE7TJad2vx1ZbP2azC+nA0yhp3PkS1I9x0SPt46kmF67zRnKODPaQyzFeEvg
VOHeZhlsy8eo6OD7+xOtvFpVdESyV7ry3hMVn7D2+RNeHaKnvv6cF4S+Ggn75vS2ycUVBGePIcFU
lQplp8XpJ0eFK5QwTeu2LSrVH2pYxdYUUCrOXirGWdNNGAKASPGtXwK5Vme3JXJnnLEu4hp/J7WV
zQ92dXhPnGK51QdE6f54iErlaD2IX9Bv+HEe4Hda8DU8sqchgZuGfrkzkcD2Ob9VahBHwSFBLdNM
MMzr/haIk6F9P95vqp1bhY9+yJ9J4shgMOyz0apxxmNLkuqbWpe2qAlz/YXI1WaRcqjlcVDwrXYf
LYc/IbFmMmqGL7YD8ALWmi54qQnwF9abQkUoYPddCdySY2dMe+RyojeUEqgqKOEPWA1Vfu3DUfpu
g60lJXluJsy9htZsAEURCJ9GXLPR6q8G8Jt9ilNqPG9xts80sbFJREir3XoDe6S53dmMCCLjdxb5
bJW6gxLUIOsfOsMah64Nyhef3DYq8ov3AliKvdWvD2F/dKYTKZIonbhdbkybL50tmY4DwYnQEgus
3l5SGvOrFTuQeIIQQyqJotO0kXiI0zjPfWs2b99zWZuBYOATkfEQJ8U4l2d+l9WgbHRb/40glWmz
PvsnzrGKhCRbkyFt9tWs1CID8SUTjBqnahVcdxMACvgzTgiOePcmYC3JaXtZl2fksshT27UN1mm1
n90blruyB3mCmnSJQTO1zWnWTZaejX3vWA6SdR+KqUO8irCeVOr00KGhsfyf85rExBXnm5d4bijf
RK41GoFR4SmGPrXxif54pZxD7yXNCXOWVBj/K6XaXlCCaLxYfja4kheznrq+DjR95xmtcdHntLYi
eQzpVasL0j9PWOZ1Zeei9E9EdZNOdEnUww+6ZuZII+/pTxKpg3Mx5QcwH/gBahOtawR+WjPjXgeF
h5IHHHRrBCrmFtHdopngdJdwPladDTcAPpqejxXZo00QIAH8GphCMMbQ9UwvSwHL7bFUKi0kp+jo
gSuhPtVpq+tVQKuHm/MUtHxc6ilereyOX19xzlVD9w1aLNn6e3i8mMUjZszBPxg6lEapy20bdspH
fjHufkp1oKtqXV5m884Xkgb0EcaBPDRc2CxaCrce9aoYL0cUcs7wH+47SvhTMaY3JJoKzK2Rg0Bu
5YGvtulsS4OYu6kVSQQtK28AiOzOKZM2NHg3cXH4omR5qPQ/hTsoTnDlMg7FFQVEy8RBt6mAWFSM
/auASsauUrez0xGacUKQN8qNgoQFwVlZ+s0nht5Dj0MK3FyS+nIdkXjtYYPblnLEL5c6DORZIldq
pxjTlGCVqZ7d3Jvk0kR9ipqCmSApF044apgi3HpacVwJIMRjt6newryMxEzwV5Y/GC8fnpMQANXg
3n8jTb1bkJmcsFQqjwlKuWtegVKchIHWu6h/82eG0pZW7lWMEcAmwaaLl0XCApygwjtGnqiLXT/6
JQ3dc5xc64qPhdsCWA07wBb44s53YHdHqxYIpYBlSDteTZVky4kxrb675RlKcHPmw7GgigUR3RrV
4jzrJveahZ1UeXhB5O0LzQ5OViFCtgELw20/V5JnEosxHSoUR5fehTR/EwwH1t8+MTkolVUNW05g
Ti1D51qc8TL3htGI1WpdZ/+7eGgvd+CA60zfxswfBBCopcRdDjilIr9EbBAdYOetVyzgvI/tA+B9
nJ1UEp52gG+4w6TIW7M0pZeoA3Zrz/U9KM13qgrJ//d72P8AHnKPDEBqyyUnW7fMlO7DJ4q4oVhh
2ZHVFsOUTp81FuEOGMwfFNVEmLWO5894BvuV9EBtxWg4MCvAChiqVD3iwISdUlj4PQMzKQtEpjDb
M38Gdoht2XfpvP/f2QWdk1yiw4t4ne1a0b1B3lRB08eb8y668t6eipzXwCrMKs7D2VLTAt8fFZIJ
NQRXM3SrzJrel2qFFdR6DqF4lJegosmeB/rvYPxP4VmWYGe/2Ek025Ywm3o2J+uUCBo22NXQz+UA
S7NqqRXv2gMIUiQIMKhhpErjclkxGyxT0f4igDu0I0TIa1tYoet6GFMhKWdzi6OwJRxOkb1Qx/FK
Ph/orWeFJ+ZnX1r/Dx6xVJlRQ8SooMud6UaCNU/5/cW3Jzm8wX1fW9m9nVSyxccy8iU3NP8PFhNS
OJQ5w1JEID3F26iZhrUZNv7jlem4+hi+DC9w1aA8WqtC5Cz2dxtnVS6CK+x7q0I5GF+r5Tu4dTxq
jpQYAYywYYJzKXWoEYusHs7JJ6utpi6tQY3DVI6EeT1wg31YnXG1sAoe2E4dneSJM27R3PjEz9YP
Kvoz6Xb4SyZQMqbmgXrZSLuhOtNXKuIrJPGIXtDK1cP8LJVHYnDV44KeLL/Fko0F5i9Wial87VXy
2PRzIV7F66LSo86AG6WvJcQNaFKWD7OjoL4nVYN8lDe/jzNGncvDlpu287BcmTRLBjFZvUnJkrCJ
Z/NZu5YPZEXdxQWfcycpBSsXAGG2a9qDZLzbJv6SNyoZW6+bnNi4ymApGdVdgn8y+33q9+o/oCyz
4ksLdh9v5EGbjDF28tpHVUbwSiwIfxMepATLhKnLeaA2D+HUjCRhiXfjZQFhPbgf5NTscNWHCixV
CpZoNQxryanueFRJ0vv2uM/ZHAbVz7vFEZ1ivJ6Gd6HE0VicXoyZ52pSE0IcWFu0phl6C/XnhOuO
0YxU9utOWWwfoenHTDV66LFKBzo0AoihCeuMz4ImwrX/REZyyiKR6sHr/KoHsA7Z2ptrYDAHoMLo
k5ACw/CkvH/cHbTPWWWaAzQLKfD079q4o7c2M3ZjAisdlh1pxkdH+tWpnJx2vOUJEOql6WVmqcQ5
phzcA/CfWuBegjZApGBSbqvJqe+9SgL3W3vFmLdzY/l+sW+EggR379D0KSdrAZ4fKPQvn49m+bbD
CML8gprT5ihS6oTNGZBYovKGa6v3N64aCRG0+lZLEyWKGXGpIrz94JaZZSqtw5N9WvYPo7ZGgM9Q
ZKWBzyIJ0FFkUqRVmzZxFKuQWVh+ddXRs6KjPggosS5mVfT1SAC9oJPJcS02N2aaRAgnpkhFopLK
qE/G8tOwX1js+4Tw/K97gHd4BjQS0QweD83mM0zxvgxDm5T7w47NIm90cogadkSUqFQET7FMflD7
6v/KP8+tnQimUmNfSPw2LlE4pupJ9VCKO6k69nmmolVdKhXj3om9dRLl2jM5CjD65pI/SDdacfC2
e6jeGMjC4ReRgp123CNUUILobkGht82//ifRTpZVOhZQQDQmDDIrI+QmNV4403KgSNh4wmUfh4yj
7qWs5/IyQhfTDlrlFVlxtoGx6/atXM1VKqBu0IM7vzojVl2o3z20O23aVyPZaU8+VdziYzATp+Js
UFtPOLzOnahF8q56kYFLxFSVD6yL+dEsOENe+ObN4R/J0E6yuhYRMLxsSUczgZUnRfYM/6yK/Aot
+yw+/+3gYCci6NzOhLNAtDMUi1vDiCg9rAvuMZcXxNstvcF+gYQy+1sYItCFy4w3ufMzIEadtXc4
6ncQIghq04cQNoo2+m0vubbiT4rVX3Z4Ywh3hOvb7sc5V9RdLhlcUDLMCHmc399cT2wjH2P2lFjb
KGW8o1HYXZPJdgEt4jGbC6XeQ+CThMalmGQeX+Jo/+GmruNEgzOapKngzsXSl7dNcyJaMmtRcUcs
ObQV5QcrYKxQkDmdv7XG+UjK9Bzh5gkyP2FKbyGhoQdvYndhupkeFFAd9C3RZ0ppn4ILScJlchjF
PdNA03j91MGsqDxUw3b4G+Q+sITlhvH59Q0cVM/joa6WoUYuKYIpRs1cpxJXO5pLuVeWCqnAuWoU
ICljlCLrxoPS7tKXFkLPQJJTEkQYOjG0XbMRSSzOG6vHcTu8B0vQGzKl1sU6FM5+ClYMc696aoRs
d53L83SgurCO+dTJe6BTAYa8XlFV8hmunJJAEMp4eY1+8/CGlTarZMoBoY35CBiVoGtXocM08Ft9
2QiQZYOuw2rT70VuoE21LCDNt4RzDRrM7Gqv0kDYYPWoKi4LhCb18oM0gTo4a32RPXsGOKhSbpEv
Wu/zwMtQ6hQiuq+DB9Filgw5ttbige7cO76ISSYJrk8LNWpEcX/pZO0Jn5vi1AI2OWijNU02gpZu
OxudyUdLE9Lu70vuTadHIiefD18pN9h+s6BkRxAHukXBEJiWPd5M27MhsBPnnMT+zmQqentlXTum
edY+x3fAZ9Lu2Xz8IhzrMYp7HZEXAzafCTRoqNgkwWWi+oc44g3fvwQE1dO/SWxIPienBVqciWmL
k8c1QoBoTsETcZTKSD2sjG49NYVU7+DgoCF3BrFGioM/iDYJlE8K68GaJCI+EhL8C//EQg3trOEE
lelMq/bU18iv31x+N/QoeE/SuOC+lF+bZUOaYbGzKMDFnjsl7FvoWtRUV7S02GwB7sAs4eBXZ6Zs
QkGp1F0az/VH8gqXBWA6jgrbjR7Ugp35S409XlGW8lVvXa098pd02dB5O4h6dNlr7gI+K6R6gSvI
XLFJImRS6K8yHiS4+uMV/gWnWi/k2xnB0CdUkRbcOnsJI+XwdVzHjFJRpD7M/R5+w68R1rjHXqie
Hmu/pbhY9yqksND2sSgrSLGymwdabOUBjsRcCKk+/MhUW212aS6/raN8MztjbJ1a6374pBcrFz2H
bI0OmJtOczlHdotZeC/ZHkRJZJxo2GzOxzJMeAfOFTynb8rg/uBf15Utwe5dOpVsdHoH8jtXJydk
w1HUeZS9s3XgHLziPpkhe3dL6174y3bJ8c+1cU/Bl5sM15uaAEkJ5A48bLgluK01vAyrv24KDNOl
8aSrNgF8drdSa51HE20MvgP3Hp8VNJWqRLM6WTaEDC1lK58GVnqe92AlJcrkhvw8yWc+bBjTvr1K
FTkqxbyPRcn4zh6y3OB3IDgEP/3XdxGNf0fWsN5WZ/jrBYIQTCwF7Ns18+JNVRgYkAwodXx8xOsS
TMNan0z/r/T4IGaglmG6wAZ6PNeNfQrsbZ3cIKQla+hBARuzTtscDQBavQ0VNKscAOhri8c/L6Fb
jPwgQSYuMr9mMxArnWT9s9yRZPRaDzqC4FnTzQfjhFnCH39upILmlfGZoEoAbft2WTECc/xAlVdj
+VFIhm/ud7vZ9j9zLllszYRG3nT/kcWOxjEpbjE3yIPP5urt7OkneMakw58iAl0EyQkxeNMJtwIU
bHQYFrc5V4EWKMfbnT7roocPqumvFeb/TdunWaHbPhLIgAQHIgIekme3e3nPm0UKsPEOye/c6HyL
+8FQaoKv5NNviJq/ptPNrrKf9YD/oXHWPq4yT6HV6Fr5RyldgjnlbFnTccLu0QcyPxaX2iOKsjd5
gknRuAG0BYI8gvXE5oV8gygxIXef8riYD5kHClFa1E78XIkxdxh6zsEjUtZUi3vK4v1ECAqNn0SD
OT5zdyZex5E9LUIEupFg985CO/TYupztluM0XS7bp/t4otb6PVZaxcb0dCzpLpr1DD8+l/nt14Ew
NKIgwRF/pIu9WT8fpBLN4x5eq2h03xbb35HE+9jJqS3GyjcMeCn2QVBV2tvFv94nZkZv7mFpzQaS
zS+5QJqOfVbkSvFRKMbAnmzP9ggeghGIwJg+4WBxi25gvaEthLjprd876ORZZp0Ta1uh2R1IzQ3o
cdneBAL26wqaZ0/MAtsUpI0cxplI81N5HPYycPZg2xAG0dqHrbChkycTEZGjksr/mv1Bs/6hzgxj
Rk6XdgWxJCK7rvoTTUe5ZdLxpR00/2Ire5QCeF7zwp18aJXiDEZurQCRacXA7ROs2zLmxCE6zpOH
wziMuasa5Y0shAVHaKmdK5g8IfHd+dbYNmNjsFrragcWY/41sTGcbvojZk5wkEnPhZLOmMAVKNV5
Ucfp/CcKDFqHQUjgtPzgFJyDBMsl0T2Hk67Hd+bcdu9IMvR7aJ2/94FCC0v6+waAls7VFGUWOzqH
CNEwj99idhL+gcLsjMg2kGApCS2kjs3pKzSIjlTMHYqxom64Q0ymXdhAwMBs+aUXCj0CleeerpOf
eQGMoUzLayJL2tPlersxc6JpIGvpc2OxNWW5AOoPkaxWc+c6W5mRA8DMIdLVLC6kcCEekYeDgpjj
EOueFPtVlcwoirSqMaFFFQgMpD+dYucW2ktIDiAp4iAs0gI/i2qDnVeer0O+a43ED5pjOU5z3js+
FX9bfj5GB3RodkozXH5/QEu98/YAym3KsMCkgTCTpT4s16bkVmi6TUtq5VHU9AVZiQj6R98hYxHC
JmW74R/a8rZ2a9EOokbdyk6+s3CjDIqlq0zKZnVj0n7pbGYWW2/eLw1eYmU+6WU1pIHjN2oQ9hIr
NrZFf+dLg3S28FXlYpN17t3pZti6UZ0T1e8T8plNzefoLOT2WH5V53LUeTyuszqd4xMZH1dmAAdZ
dXnENzmzGOIlGAxXNetmITs/eGnJDYfO0P7U1ykgT/rCaz4SIrWnRV9M4rRUa2QJksNNagSUaQNB
//QoqhyWnYpO4ocOLcDqUnpAzo8IR57ulXM7xc6FsXA47ZP/wMwMayf2xI+RocM55l2h6EWC2SLi
+lz7K5smRFmtXL1cP1XW+d68mKWXjQvOX4sWtFV3hlzs2PPfiheCU4eMFJgjpyo84zPM9se614Lz
zeH+p69NVGd3TrgFwupQresNGO0YMjsNaFRA9Q5hdSxQCrxOS5k9bNCJOBKFoW98ImqEzP32BFaM
8zey21ojx2OpjWGqPeOmkZaX+cEtniROvd6o3yhQzZSDXNy1GtVQX/N4M0fvgRKKDSPED5WUcFkZ
jMhHRu/gEUO9yeE322UpCvbR3Bn6B3AjwmJ5mPVBvUvNJWesiSl9XIFWj6iFwANmJ/ADZZUYQBM/
OXP+eWLE3Ew3XMxj2TQfuBQsE3QESkO1a1im4NVLn1g50931/1NUA/WozOC6E9dL1vdjKZ3idIws
W1X115abxyJ2UegPWiNvMCq/HhIs8BBK6H4Dqx8ld9Azlw22iVRCJAdEZEaw9CeMmCrUseM+iylo
Pe8FWh3l9PjAZf/66A7KyXFGa6H17HTebBYeha17FJw9yzBT9bbCSzi2IEAwWuBiqLwqpyHVO+LH
8AvChIr/2w2mix2YFppPvTLe8HHbNJapKTaImEtykEDefT89Sn0+0PjQOeVmTqwfmWcC6roWFQPX
q12WtKVJN0p2yehNRY3OG9UVFFKlGfuYl6uSw4kTGqGE630CKa/PYVEmnyIF9HeEEF5/8YXTyNWY
14eOr2L2vweDx2FjtMC5T06mXE/VvTttA21REWlxz9Zbi5pIBaRmCp84QJN24VsPB7jezENXTsCi
3oOqv/Jir4duEVF+lPWEJJdyK57JpIswMg7Lz4mSP2aYWxFiXbano8qNpqrYJyeNxhWJstUgppEC
XVmRfXTSXIuQvW1plYkxCEuOAhaQR+BpcEe0sGrxAs7zLs/XlxRiH+5S5Y0q69rJb0ut7RIFsqGl
DozExY2Ara+MIFflT8bvfkj/i8GOn16i3lGlTwQ3Ek+tNwa4KSQeRlQ0QALD10smSa4tqMo86I/+
mFx23Ok43gVriwrG7RomKzs8mORANHIiYG+QtiXMt5o4ZH7vLe8xb1AdkS+rswuFTkjPeNotqz8q
00K3EFLRNXYh2M3L7vouBQ+hKZJk/bUzHAtVr2DEWnwepIThfTTsAGfYvHJojb73CAwEWatp0Y+y
zPnoexFrPzzzMbljBbmXMdaZkejyLyKpVs+BQrKwZhNxnd4/7B9sGKb35w/RBUzCrsH07RED1VjC
2a5ku+1b8xvTlQ5eWfrRHwDLK6R/68nxvGJEWTvbJp2/D9WPcxmvOcozgew2WoL2kc7xx+zO6CRB
PwlcGlRoGUyTDUdpMIMHu1wvCtWmNAT8tL3JyoMDFghbkSHsK07d48Zml8p+K/xXNExwfBRT5kGZ
q4i85ms0QJqWygYziESQtYTEPjUyTBMreahBY55QfPVrmK5xomMknLOYQXKphdLeGPH6pN+fTQnd
HFkWlGaX++H6pgeNyk8HtgugeQbnJSfDitK4yEYdBLLo7b3UDjN3P/K9T6KraR6nt3EBarUorhDc
0dzTvSv03JJ58nczwdsghTsHbEljBPqYIBkbEtoKNH2iqQmfdT0gWgErkKFnIBaVCAeBj+hy09Kp
O3m7N7Y/gwM3Qjna+ylktZtGE/7dGHsGfp7yX8w1AtVZ/DObANutm75HxhzDMHWd/fjn7U2LuUSv
VZ1nojjteCOnyzsgfkugWLlqzwznXXBxoGIDIFxszgQsVeuYShOA7FVvjWzJDcXK950xCjRMPYH3
L8kuQ5M5nmMDjdF/n+qTUz61XXdUB5Yc/tAvVF2nJ4SR0DNbITb2exmnbrk1I1ZM+hy808mbM8EZ
tstUKVJqUCr1AzINvotGynB/0uzVXOD4SlBi3T/tri2WjZNtB9ekl0l/YY3Km5mxyb7I+cXCr1lV
t+Zd455dei2HEGMhvPFRhlBiwbzDZov1qkW//hWQo4VeC/Z6B7eFarm7IYmvl0Gy5hvqu6Q1zL9S
AIUAgx0ink2Ivq76VAjGApqkS6NgIo08qL3gzBmURNYl44hmhmOVW0dBfkccVfu4t9mivmqoOl8u
fbYAkY/C73grOlOkT0X4V0xKeVRB8zY1SXVgPBZIsL/Whny1ev9zbqXG12dNoxkbl5hltDP1YBj0
/Ed66KVVaFmulwGEacLrQIPDrCDDpisB1jLJn6A8HAJAfAYRz/wjbB3HiSDKZZz/VHUIA+SZtXw2
UpGPAOS4L+23cjaTgdgs2lLF3T+R4DPM3QQBCWAbBmn5ZJnRjjZNW7PbwA3ZVnq4/QgBjasYAis4
tIgL0Xhre4nrpU1Wl/+L60gjA2yyLyddD4HuqhXwz4U+W0c5xXXDFEXuJ0f4+4A4M2s8v1uGa3Fb
Wt+5id1euA4hziD3lwRA7YqGL/ok3hMjX8Tb6ABbjwq/PsNKgYNoZh0NUwYza5CYJAXZXHuqBCuz
BeD9kKRNfQSSc1u5hmwHuk/d8rI8XAb8Nmhq66+YYxzvzsnXVN4SvJcozjeSUlsjatgVpfjiv0my
HiopqJC3Bk5e9BexFaR1D8H9I+oA70qA1upeQhkWvMBxB/ppsuebIelUa9mLy0vni7dQy0CDWTxf
XgjssjzLE79RcKzBpzM7p1XiPqeCK0VDOCC9Kk9NDb//YuK+Nn2OqP61FnXV+h1E9NqxG1MtdUXZ
1f7gv7XPBTLaPOLHRKAiW8DDJGE7jpCUQWOyPNkEmtYrYKhItU+geQxIp+RfzNrZj7TIl9R2PqEN
s5HzmotJcbDDFmO37pb4AENlJPY8pFh+xt75v9HmzecZIqchZUmnLqIZTeOghUcMw0naJ77Upv0t
lg5gQ2shmzutK13yBcKw8yj9RiSnpFqLBF/AQf34OUBbWLTtXMhDzlp/TfZSZ+5Pa5d1zMPzJH7/
ykRk5EQjnJxMfWDdBLnOpTDz04M/NNBDEtbO+DFx/fKno94c4pyT301MRsxbMbSch+Wcix9G+dwa
qLraOVorlRc1yaCVnKW2yTnpTkDnXwkWjeohL5LYX183OOCraJ8ySl9aLEL4imgWP0Bs95kz8NQU
PZOjsI0ryEvaTeSUGkcMr+HxqvhmO84v1SbHi49XUz5QY9LLTfRTJVWwpXNa8b7G41kYxUUw8L2Q
yeAde7GqG2JDEHRWX/MHkIepCnjM3yZDeNJ57PcikCk0zVS52Pr5wK7wpycumayzpt2/Jx51n4er
QD2rM5ZPJM9grlh+yELadoPTr9nHbLsQFm7xsf19CeOwBEEAqDyjRf9NvQkzla4JvRZKWLVbmVp5
ht6ckJRw9SetBuna+u4sfoioUos9ZYeXekGv/SKgsbkeOraRUlItzWNFfURIIRfAmNpafBRkbg1b
i4wdcv/L2/v5Kv5lMtTj1ykqWqO4QIGIJoAphvMHgG7jn/0FtBdhkPGZuSA/cYb4S+lGgKm4y5LJ
XJE+RrRvLWzLAI+iJRL9BxTvdGoUZ8wlRg7V5ZX3G5RVGw2erCbqOaXPw3rnxcQm41UtjkM6AYAP
5aUIeKN9eOpRLDx5WgzaAnH1tIzvjcbgPydotsoWPtFpNLby9qaCFZFmL40G/5IjHJivZrtjoU9h
ed+lxjOhTKsFi118o3nB6gOmBwWzEcKbuUpFEEw8LSD9mLfi9qWsKdU8JL0FNd6OsJOYNBlfd2zP
rApI7iu/Hchl+yupYiNpyzLoJ+REcylwx2CeM0HFNI6S7Tmixj4K9zPgaOuq94iHl8PAaEd/++T8
zi/X2HYDLx3KnCsnExgMJG1tcY01PsZIFNYaWFg/DJUN2oOkDm24wTcKLVk6GMAr4DZnBZ3mOCI9
VT0xARO03wY6kjjhhz/TkioOLw04+Mq7FMH3LH5KZuMU0Lg1LootDpQCfnYjk5BZAqJ2Y7W0pvx8
XZe/rMiaNBdmvNcAo8BBsML3IHpHX3PIPL0R3YdTrrn3rDt6HOXgp/Y2fbpWATbUhsLdao229h32
G26lVVywy5DWUiXwKAGVX2MI/Sk3pqv2HxjAdsmzxrXzeYLjcUTlIK31bMdFUUw2tXM1IrqXzW2g
4vircYp+tXiFKPIlc6wdE9TKPO7xvM2/7Ti2MAZAKG9KzrxdIJe2EC9IqrKkp+FzNpvmFGe6XLqh
u277gISRxxvsuPp+h/RNZPAcmI2vAF9ckKFGdJUeKseGrDbxEO2yp23oiuDW9w/d3RW//mnL7z+Y
o4o0+e3XAGrmjwTm81Oz0AIupJjnCtp+MycmkTaB/gifZMumgoyilvjUHzj2q3zpeothI5+qdF8p
VJ9P4ON+EfrqN9cK9ra2lLSCLTQTaqoK1Due3PRihLwzNVc1HFjt6OCv019RQpXSIW0KAJIdrnYa
R6QlPMWersQk5hFuWJ76hA/UcPeQiooouexLErK7EnE/ICJXIjQhoXLVdK5jqb3Fa/xEweYxAPTo
iiZhSIsrbwK0xX/GChbTTNqGieDtk5GAv4R0oN/NA9E3KdQu8yG1ouPPz3LbbwHQDbbYSyFMmXz5
IRY6QRTMcKqr76pxguKZ/7zFnmCeJSABy0cUnTyZC9s3CdTyF2/sq6R0A4QgcoHpSi1kHk91wupt
VS021wvJjpuvLRrLrb76Rh+i3D/Jx/5AcarPGkpH+4xOpp2pE7L+8rF/XUTmXolKCN33kXqBiQFZ
502VdUEhCwnLnITWTY6ioY3AnPySAP8MOkiFbQb3G1cosHvnBDkie5N0QT1IrGyA9Yi6tIrbL8ut
zr2msOhURjyEvrtDBBfppLYmx3vVrCw7g/GXyaJ4PH8VoOdm4pwvW63zZqypNPXklmOGT5PkqU69
ksFRQIr8NrlekOQuIIUDheWZ1ujnUoaamVkGuqTfwvEwbGRm0d9/khWE+8FJQNEG93b8RceVU79P
0wxUQKKPWvmPx8fOFr7tvpks3ZOENASdtu4yVzwZU2Q9CrDn1jg6kKXknTGvZQQ/UMSeUCppfoyF
g9yxt8JiE7ZbTSZfyjHr8EYG82cXTck300UZ8J3cnv5RfvRmg199LhEmHxNoOvXZPdycl3PzBKdn
KuDci1kIdCn6u3PXyzOi3MzWM654/OnmIH031diQX72HovB2yMQzk+dEhXoXEEMbh4lGRGCieX/j
OdJlgBHl/GqliJ1X7TG8hORMIbn6Et29y7djQ0o36y09sE9KSqbs8MDoObtvPqgZBQBIL5XdJQ/N
LR9q1Ld2Zmmi+sBukNWWqozMDPLur1ZwDyyYRZrZgGYNSrhObLfbNb1uh8IJqv4+ps/rJVbEMxAe
Btw2CW+HKa9BVkmjz0WSPeajfJuaNKDeAoalp54kFLLigIs3FE9HB1FDe8jbqZ3wsLdDMzrU+Ecc
73mxlGkVBt0BF0RlOyRE3Q64cDPDohgev49se+cNbmanb7utWuJaQYEuL377rToBC+jbVQ70xYcs
5hgegvyRQAMu7ER4JQFIAiBuGTVhEvwLh0styP0yEBaWPcrV6d7bh9J7vsvtjWG7bBO+8h0lYH6M
wRgHdlDRO31nYn8sD0dyYCQH7LBUreyx5M8HbWwmaniiEVXDuIp1HMA/SkpPRVy0vKn3NPEcMwW5
qYyUxnbWR2DAus5+zw6BhO8H3samm85Irnr1Svk01qoT+htxwUPqHnIZYT8Sc+/0mMoRn3FBbbr3
Gydz6TMMW5/Qx0feDPs1QLY7kxTIFVY+fGyTSVKSWtmwjc5BD6BUHq+PiBF4BO7Mg07+XfyiZENL
R7HpCkeS+8GvImXEH0aTSvoAuISwEppQn1AKBnkj6DHw2FfFjHMmOkcIEhRRz6xvpBGvILDkrNuw
ubzJ9TSmoWyN5u+W/729MF7Gx/XFKOUA4+y5J8l5fe+UnQbeMAT3G9HHmSlINmBniYJQCH+6lrt9
E5lNAfgRw0NziKGhSmGClvZEw8utUTC0zQimEsq3/suw2kMsse1XeqGMPfTpNERRPaTAa6VLBWD+
6nwPCokivTJaRCad/YnOL4bz6nM0ToaubY0F3Dj3OoZ6UxH2HpT30pKKWPq2k8HBhKWCNKpPDgj4
7X9is5f7j/YWmWPfXt/U8csRyhTOm7rkTGwtZYjLV3oxOA8oSBBbbJOw2Jk4Eqs2KqrVWQkltixr
6e7UhgJD8RHgH9Ql+mHY7FO2xJ0bRs2/Z1ICGWQJVlW77ONV0I0qR8vviA6EB8Et+8KPl+YrS0kL
GKNvs4j8X+BEPQZDpPnBohvRWlSqq8NcUyQJDCoOfBVfciSFdEPu4X+w1XFfkXMZyp4stYChzAUK
FgVTWW74+09v1fJ9EItdClBTbdZaO/wmJ4t8stKUlDe2E1FVQ9EbHOraj0hZpETa3PTrZ/v6g0o5
aQmn9DdEAkAUhuP1nzl2zo6z5Tc7iYLalS1eP1YRK1lmNKj/5kEUQV6JhbuTXZ7TkDd77Q429Mxv
mz1EmqxwH593hiqqAl/VG/n7kkG/074YwW0aO2ZBfOD6c/XgLR8XELHZI1KCiJhcjJVPOFH6RqFB
KuVImuEc24oDfrO9zB2HxedRW7pAj0UZZx3or8V4KEU+6aqb8fQFO9vIYWWiejJgLuZ2ddAgKKEo
Gmi3cmGuEItzjtmylGgm01UvP2F5ZS15AZW3K7AHsE7ytSVNA1b+q/QJ9vT0cPcx4DVAjMBptmxh
psFBh/Ecddsn6Y2NcQP93Bc16smslB+ycUI3PGf77nVvqrV2x/PzqqbSn2Wmrv7AsqttX0KCFXac
DWMiq/iXriI/1WouUkxeqjcUX/ZSh5buSFDMzXK7ij2kj2b0UHGrxy3+bl8TkVTp8RXatVaVSNr0
2LEkCET5zyoFnayX4len1D9SH9pDHLv7bVa73atx7LE4suPfGXWuPc9esGwyfcqY/vLxXECDf2qA
+IwWgvFq3FxL0WQMHuUUlj4kRHGuYu1yF4xqrUcCekFA2og3/MUCzfPUC54uPrchwnwrIOtUFVMx
QeKARMiD9vHUMiRsNR/vbAVZQBsAU/doyTwDtWMLPzqc44o7A2wzV76n2ALCsUmRihJQZx86zTD6
QLeVePK3Y/quwZrUMII8SlXz2y8kxlasx1d9zh2nSByLIzmHcobgDJMMOWUn5WgNWO3TfbWv2/K6
WEHWMaClRwBLA0JBUgAJqTbsPK/SjoBnEv9rYBm8j7a92sye82ktvfGQ2xg6YtsAd8/sDy5lYC5w
32Z6XfilhVSGmflnqoLonhz5RN2O+8q/BwbxG1owbEqB0PnJH6S2K/4mJ4Lt8Aeq4FmT6iHB2O5A
PvFo9+5t55kJEqFgy5T3yaAHRTv7SKpEdnxpgzZcXCQvDFsZaEF78bJkXzevgPiVn1FQHaL3FWFR
Ohtt0IHd0dfQdLGnwXSnVnmnNOy+7b+p67/CEhK/l784q5bbIBwLQNlJMIrTuC6x/pClohfA1diW
ELUsxdzSMsNch7XS7EK6qWXJofdY4yYt+yfniyFC1igRT5bqlqTjAvesGp0VoTSmhXPa03SfCRVt
DvS1AFJvQ0nmHFh797fvOkpuY8O7K04gr0kX0rMQ3MZT1kY+Zd5HEfgaLgq7/XRuGiV/rksAamqV
aboawA6MMOIkRJaAgCjHc9401JJlYdefL/TDe2pAa0cZg3aPiqkw+SWVlrqGjuuJpK93Ocv2yEUt
iXFxlYBuGmfFn3REsyA/zXF6VrMddFkA+qvZ/rX3VNe0gjmPN5xgoGhn2kmC5lVAPCh4qejobcP+
9nzlrijdAN1YSX9rsvN8/CLh4U5gG1E9syfBAF0948PSBaixUo5rhwZswcgu4vYree4SDK+6BqTs
89n57F55V5Yx0P7V12imfPHu9Ro83imvsablD494aQMFWvJxV0Qb+Ha8W4QzK4qq6eux8uAmkXO6
Zxgz9rN4Rz1qDir3DHXtld5KrXlkc3WfyKbOT9K5D4K5y4XrVG8yabMtRlmzuq56BIF2TVBD3PSU
4Ng3ma922VsIVabagoyJ9CF/cDxzjy4e7B134/apsegngi4sGY7EaiOlHZ9cXeJEcU0CBAjBpNil
33wrq6TH47Q1p//mgvEidkPHpeDq3HhQA7qTzA70G8kRo5T1GWiEZVEASiADhO9cPJ8fBcS0/3rh
CUy6m+/LO+DqwdBQ8ZMpHFPOKR4RVsPb6VsrtPbIugv9CW1oPYi+wyFbYOz2EaAbQV2W9bOxcetA
tpxz+9uU2aSjBdty+vkAGIdkNviLYOqz02msf6GgiP/ha5ujzuSc60fZ4EIFAOTTQxlrhxNAgqNh
4RGVvACRDij8fHkXX2+TVbSilWY54SGOh42LB039D0s9fXw+06ueS1rJa2lO7z6aU+aLhbCu7LG3
HeFFzFuII1202p23gB20ZL6ujjKMOwVwO/P61lQQ7ox23+17liO7CKKC2pOvCx3h6i+js154TTgq
50IFlCbNsMHzaIfkEz/rzkuBHereevtsutROpk8VelTkdbJCCXWQj4Jwp5P0e76rKos3+xMbYabT
4zefRfYSdEByP4tFazpwzddLUJzlzB6EaC32hboeOaywi7btebfAkunvuOF7kuibpo4nf+V4VZYb
4XUmLHb9qeDsqmECbXzQQpUmo+icwPIMA84Cnx0gzXUs0XN6gBUyMbQPX0LowkzC4hkSMuWOthhn
ZYjJlASS0rWuHdujyqZSzSHgXrTheKPdZ2IgIrcjpZBbiJY/CAJ5I1O+3QI18GBew2DrbcuekkIP
RjpDFxJIMqMeE5mXtm1gji0pX1qfIXRwoRn5oeIGse89SMrYnBVXnO+ckGn3xnJQN+1Q82DclW7D
gTsMFQPM5k09g0nfpwIyhgtqX0LXausouZ63GZ86VjXKKXN3OIV17pbiaDuAzzBhkJz5b9xKseq2
hj+t/UiTdfPwoBmZ0yNvMITt7egWip/49By49xAD0fu8cxmKAbFG27gMsJAZjgD/so6+XjSmIlXV
bVmMQO64kNtwFbd2R6PAOQ4xAZZ9JsAb6DIkbAUvIsTtkx2FWDNQo7ZShkufCKvQ1a+qltJq82z3
cHj1RybDzbroVV7pmljH0x9r8seF45Qw/XdVFzSskaP/5YK7LxDNBQoaMWVvXV9057n+UT0X58GI
tjom737bA+ZJEoKfvOZwggkyHzfAvywzPdvolrL/1aLpS2y68DlmZSQtZ26PbsEgoGFwBNmmBfEt
DAqS7CrqIygRy20/4+v9V1nMxjZJGpvPkFVK68OuGpuirYMdPFqaZ7nH4IXzd2KLEQ798wqig/NR
Iausd0TAbSbql74mNoa9DNm0srL0SMqp8bj1KZuYB/8HyOKJ5MPLFqBBKrojWP/uzTHB/8Fl+pIB
N6Ktk0bD2eXaA4K7hLZI8gLKO0dHQRz1jd1IPw2WZ7NMml4YEakSshZAjqL6BqUkmJZ0BXYyD7yC
Se9J6K2nJgkbuaGQYHNqO1Xas+0lwbPxAVMlfl5it9jn7lphXLbzPDF8vRo63PntM/cJd1RqkQoz
H5jLyfV334uK8srhi3OGnn4YLHOMZGyG9smcJPfmv4R1oYG7iaT2MB245Sv0rCk8wPxDrKDvbCVG
RO8/v2GMYBcIbI2k5Dr0kyf/sGNW1Wg6SNubZ8v3fREApLnidW1FRwDdCU/39hqfotlQtKb/cHwV
F3H7QExEsujDZpJmKD+2O67bFoUR4s7zmlTN7zIvsR+OObjOve/DPB8iFcJXtNS0C8IrBQjCJlvU
zZ8tHGw5vblsfKsD16y7RtXo2agXgh0dXlxaHCjvXmwECNHx4oucEyACSaRJnfFu1V7BBTNg4Aoy
EOZxlejdZtCt9BrboscWa0xzJMOaBOWzI7Uk9kZnylWzqAybEI1S2G+eh29Ggt4DKiujK/RzaMJQ
sN7EvImbibafM8/xfu/GuQ+JY5hxzAd1vYlq7DHXYRiaVyj1kQbmM87ujPkK5aaCqBoEUq8oPdwn
HJOHiLln+J3oesowLiSroclgU8Rzx+p94tKdP+LMl/ECu9+EcNTpm4wD8v37TsPni8bWI72nM8CS
Q5Xx3Brzn75Zfk2UGkJRRqiII1Xfe0emXb+K7nx5aH91jcNC5TMPH/5yuwb8+QtR/SdEIeI2VUlt
NRGo6pBHMyBCDftdIrD6ml6Qby42Vm15slkERzWW+uyy9gazYMtkW0undzcX7qKcLUNmG42JVxPK
TDFtS1kms9YKCkPh+ljo79yVDvZPnN7ubjQZelGhuzO7UEAXKtdPzj+Og86m1iKjaUnjx/T9Wfx5
9bJzbhZnSwd2QYuEQjDFH0E4iKlLGS2L9p9UGe93muItVO+ZV5b7pTBaMRyEL2Z/77KujhRSn8MD
uzZ4f78jlmDelG4rm7KH/m0BIf/PFtJ5CK37IWwjMTvqCuhWU1P31KDN8dLQzIagyiCh1vA+A2ne
FJu0Dv8H80sQzNuWGOEyNAjsOT4Z2+3VG7w9FOhOeGnzuZ8gXkUar+gLzWRDY4E1X5TtcwYPwQS9
+Oc5hugDLY8ZsllnPPvUQQuagkpX6cxb/Zn1jaMOhfl0aw5Xo/+bVxSud7MZWgo7Dsu1gN3AQM4b
aznZJeDeowVAvqOdQ42GMOBDwhbY6I/IISWp6oyk1I3/WxZVIzi3+7OkZXdCiQonafyg+PRqWDAd
yU5baY0+YVug7jN90gydZn5Nnx/YrmOPwNJLVp2Fv86tGXBcOejH8D8IqfPxno1POICauHs0ZRGG
ZMEGk2Ti595vHW6bVn3lwYI2yYtNvy3dNBpTRsu3ZsgNeayOLCjicPqvRGWG1w8sEBPmTBz0OyTQ
TB/SqktPo95X+J3Mbe4B1S5v0cYY2myEhNm7SzWozNQMfUkF0aOjUD74pVwZb2F/ltirk8TS4Nys
JigtL+0AckrXWAaCIu9RsYCnnUFkGKArlzlz40vsFKf+hWF982Uv3Z00jpn+/jLv4Jp4CDs0D4TT
O8WjMqLzwbYSoPJyPsBagmRwCPsFSy59tNzbEmNU2ZR10l3EeM1IwH+RoBJQEMsU69b7SPXAZYMe
QgbS3II6VRrXjvTfuVF9K9e2U7+06o13hMYt8wvEe9R2VqyEkGS4U2VeH/w2K8GUgktS4QG9Nh0B
/V1sw34fvE4yIrgKrLssxJAxVpj7dCpVi8H8Zr8uZsVwvcsFMRGgBxaoTM3dJqf484p7h96g3Ycc
RLl/+RKJHrnA+sxUmHxQnZ5y0yLoRcYvr0c/OruBQwLD57my7r5KEaoNsczVnPa4EWnXrVj3aR2y
do2zDN1YzTjOTARa2aagIAIZGqGSLgE2qRqk74kSZbgbJkgeJJ87TocrQTyfMvWYgFZMifrv0k14
ruM6qDIiV8NeDmkoqsXv4RT0h9x0Sed8sA7N3gbzNR4tuk0zUjMLjBQwLMnBZfRweepGDjIZ+qlJ
iHWypM1DykvnnbEQ+FqRFs8rr5qncTY2AuCX/diSTpsM1oBOtl0vHwvjoiEPfYDwxdZPwYslN+1d
iZdN0hxgRg3JB3rQNunzjDWN73MUvoCVKsS5Oo7eKcz4V0rd0F8plzT37Dgl8kIZ3PGM8pXLIU3/
bVUvGoMiKxU9xiJUFad7li8H3kKKedsKFvJJOC8cq8jO4Y0DWelnvz2+M4p3PFE1I4sUUFJyfT6d
k2MIP38oVfGTKhzaa+IvEMnWW7LYPxXB8Py6whBgy7433ofh2KhYe4xUJp5b2zdAPPG2hqOfD6pw
ZvLeRxaJkwFHrwZA9zPgJDqUZuHxkUDyhnCEixoxezgcG79v5jaqE3gweddjrCtZuCKxh4SoDNv+
3ysDcSl6f1z4Rsd2C4lcUPC2vrGpZSqlw6LWjcjjNDEKEWE/6MsoA1cu5Y8Ul6lzU6Zp2MEBYh0w
Ig7hZtSrHPyG3ZPTlPrPppQ3hBtmJ5wzYuNWeOxZvxr0SaSMdybsY+8in98iet7kzJsWKkrruMzP
pj0SqwKaA1ytykvZCBdDxOrN6bPiM/lfDxGqGKEkYB/G9jukJYUuqR/CPx58+iMU1zUiB9qycLZt
UkGux3hLhEMXSHBmMDXVeA7eD0d+u78+eVuGfw7swHCvm0xbGTNCZcwtEYmYxhNRrlfQkJJOFNpn
uwTtzz0viF1hRGMCEuYWdgwXlsTASwb5N6p5C41pXke0FVJT2ZbyBNAf2cdcamacbzTr3a0HRJa7
c2+Sk5UL3apxMZSSM+V188sUBfe/7pGfEK/0MSC3JYIn1b8mME1MqnGLW/yrqcg/iyo7tg5EK5hv
Q4pzsnBFrMoIgMqqxUebPf73t3j1mfDo+ilevmlrFQAo9dROAM4Xk6Y02XOqWcClIe7vPhzLZqd+
VEXD6wlZQW2TafYWqDkZRH8j/7A6XHR55vcpV7wRuFufHo8O/Gbpyc9dyV7EmFb4JishiSJSxpb/
kcyGfVapICbr9tyiN/bty5wlPIpeffL24u2Tkz8uWG7N2hVFg8oyBsuYAXFPveLqhmM/uhIBbni5
kfme27rRHzwRsiN7eY6L4ozqrKVsyjO4caGm8Pmtdr7X9gc6p6dDZ5gY+KyKkjSdPrUJbPPnokEj
wVmeEQSRreb3KpWpcfuHn2NXFt6yEpQDpZZdP8E5y3By91byR0sArlg1gFkdhXVdhAVsdhhPqJmR
8HXZh9nG6Vq4SDCe0byhzwII6xORSuFtldAVLN1J9b0lO1/qJoO4Nb/cb20kWdNiossqi6ZHmgym
/juhDX0oY5q5fjO9Gi9HyLZs5CZNamzMZlP4g+myhQivTCuU4sXzemtL2u/JPYj6Js8xPX7iCmkX
cA8O3J+2iO4SyPe8JgcbIl64b5OeDpoSpnnW3pX/RSAI3b05BwID01lbUdFTFpg8ezEpnbrKM48t
Xm6wnuPn/CYs+FoDaZOmgRVYwi3XUPWSEVqD4kBDRMiuRr/tztHegTDpTbZR38c+aKEyg+/I/VGf
jWGsqNViPAS/9Gasuz1W7Np00LAPyi8Aw9f4oBb2f+DCrkiD/zzFOpLy5Vwy5mP4ode/m/6lbsA+
OmhTCBRiYYPquqiO6nYJUW42hyn/kKoxXgI1kJpuh9G1IR/NmxzReLmqP5jLbzyQk2LpXzdIS1dB
8IgJACJFM/ZM5P8yTR+PRblXwUgvJxxBG45nYDh9IQlkhYFDR6pc/v4EWFv104tPOlWot6HlHvrI
+BRfyOv+GdefsZk6rsyhaOHAI1yfPZmRL5TwqWdeomiYf1ytRPEyrzHI9PyUuWWY5qPD5kVfmSz8
3mZbsa+nxLD5NrReyCVEpEY1zAr0jcoaW3cE+4XXlIRjBDcSGfivl+bETFp47NTxu8rCqnvDNHgG
4fJ1zCJyDgwq7s5izR6WNikq1seo8OcWyYVyEAfcS5J3T/epfhBd1YrxcFqZZbItzYxAFFtev1ri
4fSW23s1+z5G2Nz4EAf/W7maw+HjHxJdXbNTqYfJ0HyKSHqhbb3JBhktPPPl3QcETfOfOGgei85C
X0exeV5ElH75oVWBDSLRj/3Y4M6M3hcIP5EnZ34noyA/0XGaWcqdS8FZ21pDPhYtxb6+APfwMuVy
FGGe1HKtMC617agWsKnsBNQW32tcDOkzi1cPbuFRbdtb4UpJc6itf+gugGYPRr3dJiAXqEIU5PqF
qf9NM/RdLIwFalWNreY7vs5nyzESQ651cLXqwLqN6T9XyDLnaRc8mNI15buRm1gpxXA8lcUD/HAl
qVZXw2fMSXlkdXlcrSjXo6nhnfFvVcZPgOKDHMPJgR3Bzs4khuFUgjyhEUNrtl+dIhZbl1TMcGmE
6XJ6dCI4ps0wT/WnooKDIXyvNRItuFn0fnQtQLRDgfAwDFMbHuLihCv0cDsWk6Rh5KvlkizIgJ6U
txktFYhXMaqnAp1FzHi2e36WVGrAp+C0LMV762xAEKPob6hx5h3HHB7YU7YsJGHptDey8YwYFwzC
LbPNdKKc4ldZkOW2vZ/3Co8NyoSSXzSVjvCOV//bFeELjg+TlAoVH9p//0WiJuieNX4MBjE42WQ2
NyCoq4XhxLWe04YOlId2f8/WzPRNg6d62Qc9FJJ2SWSHloIPc4j4giLySioVTiIvZtv1UU5lsTmT
U0ZXVTOmDqAmaZLGX0pxAv5VhDKoNQNJ0FVkOLtSAWQcX2kbHKrlf/jh3C5WlcItJkbjE9b6aGBv
qLsxAKisthbtAmz354Bmdk/wdE7JnBRTgMKHxy0gkdzMBZzHLp14OiRZG4i9xUBF2TlZbQknrGqT
KDtvfzbpgN6PdiufvWcC41WV8bb+Ucz20/PD5yQfUh0Bc8eqwtlkHIBT7kfmDOg12cSGnM+dpr0m
YxYOEddmWHcgiwM8BW2A/G+ORgLi5xGhfmCmzHS1Io8zvc6RLgOxd7pfmFe+wC0NMHWWakyy1rof
zjsMMD8wdQDdwh6a/e9hPNeBFyz3p0NPB6zmC6qoNjTyMViK+bHaYHHGiMTuP4UK6wuJG6nVi0bF
3l0kBKPr53BVNe9pgcKwOveiymg9OjNfMTxUEtAXyqutw1NN8oDxVzNzNTb4qumzgAPLVpejtf6V
ndQyi9m94TNo0WJzylfQxChQpmosP3C3TpIgjAqt8niGlyKo6mKYTe10ZZ0haid/TBxDR+3treMI
rVKMxDtUHhq2lh+mIMxoDMTAC0z/qxwY0t3jE82wJUmxkS2YA8KtPnUnnfkds1Ld1OoxLe54wV3l
I+Y+zYCW0+4HS9yKM7qaKFQHcjEXR/WUg1uIzHbRy/g1cLL0XwsZUtnyQGgIsNOnkZry3mtFXvdm
a5pqQA8I8JiFRWf77NZTt9/4UA/mhWqxGZWZBidPPQDPydWYscnDz+VfQLEofViaFcTnxtyadNvc
ZcXclsCefefoLy+ZFCPstvGbmnCCxoC/ToBZfefHSMWBGsss82/xSoo+xdjEskoZ487tkZZ88HGt
GT+wVt3W3mwnTAnvJZYTdLRH4G4r7Z5tD+Auekz/cif0PXIO4SWkjVVNzaR9pcMhsq2TTZHBM9p+
uh7HqZFLXHmbQIa8k28l2l21DJV2pPTnFMiuM0vBQhuIRQ1FA5l2H7vpJygYnBo+6/SJ7QJXeW7z
6mdHRHXJESxwoP+Vl1T5YX3C+D7oEsH8dXXmB5nCZ2O9o2MTktk6j5nJouXl92BQasYZjYwNBilM
+KQ0qL+Cm58J2bDDUckyEnEEs/pXHMzxjk+lkNdOrzdgKEuvFurKPO1UJpfnIcDxerx/2ZgHmZDb
wfdhRr7UqglR/rKy+T0g1MFHZDBIJSExTacXo46xijVwosvwVcnN2xafgn/Q92Ip3ID78Xyt7ZoT
k0wKOnIf8EGCisySSpurKLrz3dF+2/Q8hjRgGsEhTBl4fLR9hRlmU7wcFiaBaGrjoZ2fG2aXkerB
JwhuNJi/qErYEdxP2mfWBQ/gbYbNaFcVDcWJDXjjvOdCHZApZm4K8nwuE/guTc5Gdgcs1ncjTiDm
ms19H6MBN/x7OiHsckhqOJW2farIcKjsF2f4eAyI0Crxy9VZa8yQ3dkGFcEsgiHBDYIwKYzmr6T3
hPBVviII5n0EFM6nJePyXrPS31K21ozyMAM65VuMCIeuwJD8xX6rcH7/cvscROoD6QqnMXv707XM
fynYeex5kUJHF0nSDQPa7COnzNyhNRS76lyL8cxgoreREe+kySM0Qe4EoM1L+Ic+f9e0u8LHPp1I
+d+17X24XxBh7pCiOXv0OgpaPXaRPVuZQlJpzItr6mqo3r/yzAqQ8iQOlektQinArzPkivGEXlMX
j9RX1zD13qNBvE53gjyyfnVUNtxkNtXjP3mdl4bhqD4NletwY50JjB1bb5Mhq4oKcFF0Q2aPluFg
4pGqcbDLq+YT66UjtyET+fo736d1WMTa3ekR9K0/JQkX6wNxMXu1UkYI3m+1TGBJsrTZ4TqoPTjd
pORwYm7wqYffMTF5WDuODSyBGfDX0YsnxYaZ727BYp6t1I3/5gO7LZkfI7qPiDDMwWiLYGhrDKtA
RMji9owOj6QPk5R0fqSQ+7c1ZBkIYU2vDskfSHmGSOY48QWq8a3lfldCe1nKrdw3iQ/xLfC47oNR
jnWyVJiTHkxkx4Il7StNtZmL3sHkxYJS421tFNt8BkxJwXd1rNAW/0UpHW17Ua79MqK9W60FJ8VP
czgxLjzL7kh8fLe2rF+hJ3faiCrnA9pJUkSeN6qLnZogaMwpMTZWx07wu+Nf5eNsRGJTQ6iz+m8F
A0RtS68ZBpw2TYcugLPWXJkyJupj1XICZASdPxlFEMMKN55aDackKOC2qHxUAxn7/tHjqSKeCIkK
5xpuiByL4evC86F3GB5FJphprmmGxH4fX9y/n7N3dvvFjzvcyKk9fHDJXUawt+XDh5s57hjuhfVT
hCsig8/ska/ZgIsUnt+kp7xj8hKnQe9EP8uQoKdhyXMd9PbsAFTWUMUGQTB+4DX4Y5iC02pFMW0B
vNsKrz8LyLv2nH2ZU5rgpB3v6sKcjpPnoRjw1VDofZ0D7eqwl1lK9O06IcNKQ2moTYB9rkqLzjbt
n1QZLFJYfTfp0Qr5Flg+AWCovc68URICPaUU4nXvk8oicahiNABs6dMGFGabszTjmA3gouCLbZJW
Ma/cGpwJQVFbCbh+4gjkp0kNLtRKdYmiGZNjoUROwdeYdOdk82gPJRaJ0RZMQzIwVhwAnqofQIBQ
UmBT9/DEnG+X2Pn5Rdkv8j+/PUxGTSibDLlwpVzJMTXhd94eFCP4O6X3VET8m5ykomysoNNAbK2E
ruXEmHnSTEG1vOKUEC84Q/xZz+iQBHrNAkYGBZ8yyTB92ybtIIaNPiQgNbIs86haRxBvGt/nfupN
sozf9HuJUEht5YY45ooTLIJC3DyQfGwL9dXlxNaBAfoteYyyivD03JP4ICm6uAByhj3hOME8IDFT
O/x6L9g5kVgLiIHlJclXy8915vKyeKxK+yk3Fr5jJ6in5YLFyVKP4dWmwiuZnYcitLFsE+/0yNTQ
zoVnEPLZUGLlK/XyvVcGTXOM1ZrGtUV8oubIl3G0GcdxApPN+DbQ7iMpyT2k8tYb6W/QH/KDm7re
Q0tfn7iiOn/2aQ6ku/DHHK6SnvIYBu/oCywyGZf184Vwuas/i9Id23AclOxdwuAxFNhktS/stdo+
p6SQZwQTMu+/SrIogxseoxrbxFEaPXf2wdwIywmdxY0CVJ9BWcQTKQ2nYy4fftDGHoKaPEfsn05f
j7CmpfvWR9idfL/XcZevXWsNy9AlY/ylE1xm3JHqX4r10w51KatjmYiuuU9miywuVpJyH2uRFuf4
MeeLA185JrSZit+d2VXpf1lCWOUn+t2ir8L6cci14PZInw/dHG7T1PBcUEU0KSUCmw4CZLGypw+c
pDBx6IMiGpIwMyLg9NtkpiTdqvv//oDmux3sX1wA5XrhoCi4bqlTFErMydKxVTA1fjd30RzO0EIn
8rNSvUyszvWPqbUeekiArPGxJqAU6ZCZYocPnMmN5CN0uDLXPPWfqXSAYkLr1KefGKSR61FO+3Vr
Dnz5ZNvIPgvD7e/2wjoLnadyw3zbxEVoo4tZJnn3jDGr4a6pwQWLfrEFSgJWui2cpEHRSH+9Siqq
6ZvMjlqTWKTmjOIS7ZUiaptD2qTVXaO+9E+03AkLy24bNdpvoM3LxnHbLspsCqzCjiK5fRcVD1an
VKuNc4qQVJlTxk4dLuN4HhlIAzT/3zxZ+YyAQSMIBZ1a2bgh/ZEjD46BjHWeHC3C42jAY6+cXiUS
ZcSg61AeDkh29i3/NbRz00IVA1YDLZ/foOUqvFbFxicB9QRhYat0XkLMYCnocgFsZzDFxqbS6hUC
XXGdhsHGHviKUxFOFiA02xrKSfWRxOOgXsxGQFb31aBQ+6zS+QC6kCiLB0seE/FnnbKPUwTVasEQ
xkxzFoq0GENmjhy9BGSCY3WILrKalAFTjt3WeBsCyNHhUVMgVkxotiR+FR4rH9pYYko3E/v300lc
d120u/hok3TjT2CdWVJk/p+Esp1qNxMpPiJbNCrqi+WyeJfctW2/UA4wN77aRmVBYY22D6+vn6mj
9fmDG6dLk9v/by+5lIaYiS8Fw424q4R6ZA8mNHIJH1N7iQCKHS4wlf4XvwX5kEWsOjGYQkV6Wdam
rj95CuxjUBGY4oPRCBihh/DQvZr1TPbxituy/rohLVTPkfR6KIgFs3w2JFY7k3jfAAXoRwjHttKz
axagP48iJPhWy+X+dPFI60+A3Lvx0w/p04SoaNHsZ9hlNUZW64qfRr76w+wBfyqUy97MsKDz93cT
pG0I1C4CJxocdwSp0MzGtiAYKx+uBGTjPe76172ZHE3JOpWVJENW+uGM3I8cOfq/ohiqwZVISNkc
USe0pnhJEAD55LZ5fhbxAIyMXpvA5V1cmkQaJxBi/4rnlBPIfQoM4++4KiyUyXZiLlpk6CQo53Id
gcyzH3BgqSYPO3cQiKEzRRNKAYLtexYc2CCILB3Qgh7fUI3kXhcf7m3bV2JPfq9gbYO6qfS0jCkh
f1rHaAmvL1RNE9TqiAMGRVNsWWPc4vGuc2utWgRtw+4oSwcK+GFITK7iYtoQfBXP2ZcYeTeytG3P
V+kLHoq1izrvbLPqJU3gHWNafUvCllGFZX49sSJA99ObH/NQgWZQlx2eUIMUHT7ZpBWVVJT0wrNn
g/6WDwLiBKlAXQB1llWWzze4ahQoVG76CB43uw+onKW7CpF72yn8OnJVKFhGbPnDmTjIOCdxwNG3
cfhKCZRXwsbI11Kg4EH2YY0oPQs/WeH/GuedagZpBYABSZewOfE2iK38WyFAHEkh7sUorRFtxQWC
vTVE1EKypDW5eG4HWGn6tblvLPsW5/ZWoJVL/aY1w2ei+G+MRRHsF3kLqoxBYadTg1KYQ+8exQq1
FLMbK05PAOQID82hUpdlv3eYZHUf7jcO3rLfiAzQ3khBwwjXh0rwx4jogUsP4zDujYpQQneelNUV
KV4uweY1ndU1lBw/u/Dj4VJHqv8Dh73UZ5oNwgoc3NI7q/FccAk93psafA78PO8mRW0p2x19xcs/
iK25is5oz5wteziMffqj0KcKbS3oC5xK4baCAVrSMM2YRrbKgDltL8oQaJfIpYuJsQldv01yrdW1
6/XBe3muegChrqkFpQFhhFaOp4DA3M95TXlD2nXtodMZEw9IZXMx5Yi+4TOJk911IkgMTvLlmaT0
zCsJptCXfX7LHGR9n8r8VxnqSgEoryWW9U0AT1WyQjea+T7IKA4QPHX+ss/fI//jzO9X0BJYW6fU
5CN0o3GTAcAS2mppTn2P3EPu3xMgGa+3wFpm4wa02q6g4xmTpbEqxvCV2lO5Px1Ow4xBrBo+K2dG
E4rJoi+gS7R97uCmvd6b52H4tJHh2fKSitSy/PpHAxp3Dy2TMtXpyJpRaZ6x5nNS+jTh4AjnR8/E
VgWGeRonDAb/gdWgGD3wN2udbOEGg+M41fbFqQHaRn9JX8ZJAqkthv5Q5oyYIkMm5Hbx0Ji6LAh0
HdhZewMIY+WJTVLwTOsVjNYU1Dr+4sXw4vSmdp51oISZ9mi3BLgUYjCst3LPgcBdbGoobpuvV1cf
d5IMfL6g93srgOOmLmVPNe6EymRy3N9eoOYvWYnF0N3PvAwYW56puz40c+UA0MjeDe/3J9q6LxPR
pQK0i37RTgFg602e2sfzYGNcRsR4Cd/2CBM2Lxw3kuCprNyRndRVjr/92Z784IJ1KDMsP9tViS9y
cGoHg42/u6TtDRRPIjSVX7QBwRta9+rQdUQxv2Eu1WAU3StDt7Yt6ENIABwQyTKYBy8e91w8utc2
+Utq2a11AXB4ttL4T7FN72wYL7RGjdvadNLiNfJup8kMeEVEvV1bPOPC/TCAPniEqQ2onQfI0Cxe
GCmVBmpkWTlMLeOT/oI+ekgz0uMTDEUMkKVsuGtvu/LNJKfU6+jk/mQJaxSDoY28TaD8RK0Z8sj9
fIs9IaviCVTMmXuFGZu3CAFQGbFV5DxNlBDlIixyVN4uPmKUrIc2q2fNQIMrAGRsRhGqm1wpeVBl
JH277sb/FKNDXPNndOong+nXVlrLQZ6CsIVCf1UoWJEJm6k6W/N7Np849lG04EOev6X82pMZuieT
zb6+bVVBT9WyIghOK6vVEmQR8/2R375wCG3EOW1Bz6TpxvS79a6LayDNFLvO+f/q6iZHEATAHmGf
KwNudLeYPa4AdraLYyy+JESeUngr3SYh+hz9OysfSetlMPMiTdOtBgAYn/fFoNl7okHWcqwNC7Jr
J+SoU7o3MCDlXkJMm+hFTYrIzRxIrD5N1HN8fPnqO7gmBVAQWNiwbia9+I8iIDcLMFMNrlutN3OS
ve/Lcg5uti+jvv+QgPZPO7oEO3c2/m3xTNJf6t1jWQEhNlKLLThX3XcmKNL5jWcRuPhQNEi/wdfe
+3Oe8Qb3D3T2R49bkGkXvkkJ88F72gAtJHvD20yCQ3fISfvdj07p3DLi6Af2eyRq3/r0Hu+hPVNm
zhU3lfPEKINTxShM3ciCyiU57xCb21KcKt+SfB/CkgzZnhaniKbGluKY2H5M1G5CY3RuR3rr6Jxu
A+d6Uu7ee9YqytDjw/APkR0GyKijFowZSHuIdFHsU8zE8+hpEcizKXAslZwEYwnbWqyzrHCqe5Aq
iILswVeWBat0C4FU0YiBqzhWHQ46qbCHr75jiAINQAW3IeYDnQHB0ZFRLZEGg5rOy9q4Ar2OGusr
OFmRX7jpAo6bdCAPTmklBvwdBoHlM9ucH0Q5XNMw7aeslRLc1penAsadiHuFdaAvTwNpJ2/9anxo
dQhAmxoGfPO65KVTInHBhRbLIod3ilWeUPbx14t0tdWlllVtUUtxXCfX4ygpYRURQ/3RuetUqc1z
X1NCWA8TVY2xJkQjNK45qSNHKluNAOl50RLOsx4ixJ7lG2/zjqBRtkS06ymmSZ3sYaqeLz5sUwQe
IjPV+NDJXmjBy/b3S1isH/1QiVyG9S+fgcXOPFA44prPi4/bjBi/jLQNT+o1TW32WW2nuGu924dq
UkVHuKuVMr9QkunfWXoRVfL1cvjSPr7ijhhYLtRGLIt2Y+HSaO37Vx69zI0Sx+0d2N26cyO6D03O
h8p0he/qQTWwC9BIai0CT0MIDb+mfkd7Q0bJiDTnuUJ9O2YuSVJoEVQFjMVW+GpDdsCcyo5fv6JK
zDO5cO+/WVISD+X1pFydK26xGbBvle8Xx9zv4yHe2zjJO7d/5IN8nRX5us6cJUoDDheRYvYw6UEJ
ebk9dvvPySNWKYSziwwAN0Wtr0kqLNa7C9f6mleFfMZxvEDSykb3fr4KCGAhd7eVEs2SQMLlibwE
v4pMQBd/Hxx85OGBUwNExJnjJw5k+rlLPSLwdAlbOojbWEAGptXwn7a3e12jlumnEFQdc/On315o
xlOHNa9AsYgiYEFzm/kRJyJEZOfo4JPGF4rbUEgi64NjRxy8wDZZFyJo9I0YsqqZ7JFYaqnkieSa
hTp7+hfj5yIUtoSiHB97GhjXQskj8zNgieAwx3TfAF691fQlkbHgdgWHFBw8fd9zpK5fQvQr1/aC
yx2REI6NQA3bcIwfjlTMhuA+x0fx56v93XDT0LkF1PnaSaIz6z3/oqdKj0euwQf/WDCkCkO5KomR
a0OQZkzsa1dyHyraQu8CznQsFU327eo4rVaEaMiHmUwA2QVitGDbb2XGyOCi9wonwzKGvXfi/RjV
/tICweKBOPGx7RtzviOntBvlO5+gnA40YfHiCCsDmJ9q/nHVnr/9gHX0IdprqtgQ7okvtEyRSB5d
G0acY+y9S/3ySko9NXignMAtdD8lSB952kVuLV0Ej5FVsqT0XDMbHKEHvvSzY7pQ66Rq6uaMc7bn
uXZ0ZdVDUduKb+qq29fj0vzSuMNk3EoXl6B0cPBuJYSvnp/CR6J32EimPArGgvEYqBTz7FmLxchB
V5Te1NFLBW/zXXkhtVnAgghNXLVF3YG/xqKNWwACBfPysdTOLGqzPmgVw2meKNLPIC7oFGQn/QXN
VZ7bPJvLbDAp+5R/Go/4pVPEVPM+rXhqu+bQgg1NV3XkigmqQeGrYP0qFB/htKmYwg/C2JAhzD+T
9qgEiE0/rLuDJBrOZ3euUXCJVSVugYc03sDEsGGz3jVQ0F8by/KqDsl4+ZHFldibTm9Wc7Os8JhU
5q57IiJfzTynPRiHcAkBrY5pCk/2gKHLQXAzf+aI54IvXE+C3gysJT5FHDNjAdOoqNVgCb9Q7sZA
O1N7IjkEtpTFbFb1y4lMkjbDKIeDwO/aPgejJFPgTTZoS1jPIhqmnCGTUY6vq/6Sji+5L6CvTbKe
vKHGmKRpR+kNK1aYUm7HDdesGn6hbYJGORvG1DKQPAoWLY7dhjFLY3irg+6AlEXityxVMwWIwf+X
Vhm3WEDb1wMZtuR8Dpv1vFOU+B727Ts9wpZISbijjHPZnFeMgiYoVA1oMoPovwBv4pWHnCQj9QtF
BFg83vCblXPjOFAr67Jhl43SAwuPxt+Rd60RueIpVEEVoMd4xc5tm+fMg+yhYPmwN+Q+NwxiZ8ql
A5yFd+4aWoqGh86gOQIG1q0KiH/hmeFSKf78yoA8F8HwgjH3U+1/m2shAdeP2ci8xKoP6jO1HJPA
Qqs2jmyPWJhmAji/JTqZiquB7a/thaV9oBKKD9KozdAmLF8umM4v2OnCQMOqbXbD0ztrV79BWFf4
I6o8DfLWrq9AlILYo+OfBRzAyafPypva/gwyUtNU0MQJHnhSm1y54aoAFvayoC9f34iwI2gtVENV
Zp7Mk0fw3Pz95kCVo6/EiKKAA22MzWL1yUhy0stHF+y7i3xZwEYlQHhxFKkY+4wQD7OPBF3TRE8x
T5VRSbdhbXUaQblc7DQg6UYjKRuWSnAXLCylNUaObWmQlZi+G/pFUga7PPPWlBf4LyVbOa+lK214
P0yjA9B0CH6x7IUu7UNx0+iqqbVWE+RP/cscrqZt71k0y0lJ5VA3XHc1sXXUEcQ1i/EMbiDu/Its
qQ0GCwCncMHj2rriKtoMkOAjS2MI+BMaZbIGh8yUXv5gUftevT4gMVp9Svmd/2GDxYg6DzbuKFA0
OPGzMlUxiXEHzBzXuYxCFwbkUqgBX/rOXPz1843XdJUhRaieYwbCON2Ld87/6EiW5BWfkkrjIjK3
xc1ErtbhEL4sB7QV4egVAcZm2rqeMGB5fmiLTfjuR8S201CvMmccmD6ny3SMaPzRveOqkrnvGvpV
nH6dtiquhZfUhrg+ryyI3J00jQ0J78Xfv4g1v50c2nsePeMfRmgJdRkpNJUc9vxJxaSDDYgzDnab
0g552RsgU8HSngo6kfxelI5EPu9gqIlJ69mCdfuVOdgc/wwyG87u+CDaJWQrtu9VfhizShz6Zp11
wXrwX51gzeQfXx1ug30UwE12+0zwDaBobefr2wSCDPzj+5pz80JDZwWy+YTZpS9HMNIiDyIx0Yla
nbjJ9DF7cZ0OYXKlg2CRK7mcFZl2Nxhc4rYRp3Gd5Zz0p6kERPWSjXO1++8CGcAkLzjy9MeGaHdE
easLq+fXAPzDI5V/CjBObUix8n95wxIHLCNX4rxDOkWuY8e0hs0uDYcxjANxkr/yHPNLM+N51Axu
/SmiHUMitOquFUGvYnr0n5E5KGUKKHwu+set7g9f/IEFqKmZJcPlLFhgfBLgkbmPIU4aKZF2FLDS
YVkjWfK8xMqx4ETr3TKqQ6AGscmOIEJjbLC+s+1sCoiOV+Obp/KZRPh+H1UF8eXdnoJuj+5aZ1C7
C771Nib9jAUeO9IAUYqGs0IEiyqFBkNSytuq7VglrQVu2rdvqYKwuwLNWBbefj7zBj5+x/FGMVJY
EoxrABkoc6BgRMuRxlZ2i1qD4N1MeyZZ3GdEjvlYHqMom9Vb26sMRKgVOESh9P0vcs2FyGNcZ3Nf
GAAzurG/TTihEaV4Eb/Ycdu6QMU1UayWnhFmQKhrn1yV9LtsQTXA0FbtZEICKBuMyDCrqCvj3Lcy
34nXFf/sFR69kUEjOYxNuieQZ40huV9D0oOHa8Dn/PPmqImLqlPaznBHf70y9k0XL3+jWuP9J052
nbL2q3iItpdvZGiMK6lByQekly3DKJzCJCizTRCaV9ziYFag6DJweaoJxRcHKxOdh5/o3wLtrq0g
tWNxuMXCfKMUNqe3GGuMPdg18mjjhjdy2y9AmnpE70ozPC23Q7T9cFGLnuKMNymUI7cwkIvRMFly
GECU/xmdG9pLdCPl044UE9MH6pxt53frT8Ad6lBMGYA2spQV6EQiT8faZGusT3KPoGC62X1sQ6qW
43L+vPXHA6CDvjmkhftsk0rNCzgevY1C7+vjBPIOLZeV0AIqDzG22JCueyz5K0zFiUWbNw1y6NGr
zNYhZF9cOOrnr1roZS7TuMmGHvdR6J+pwvWHWDqJyq7IG+YjBbTAY9or96GUC5V6Y0dp1mLyc4gt
Qs96Lzb3ZMW2H+T+WTDM7KCF8lsTSIfQCttLlse0ilQF4LUy893JIsmorGlp0Uaa+gt8Gxyr/qT5
8+oLVuSIn/pCnMkTObqA66QIZs66GRWKvQ3TBjy8iwLODxvOT7jDQq1rUknVBQ3b20z7dADbE5ez
MXeUU0oDO3ynfteYQsowDwi60qfocwVsYD9Yz1nxrdhNLJXNq1GmEPTehZqFAf9RfE2GVP62RzIc
DMXkJvk2v/XYZSQevxmhjkdC0o8VsIJjgeFUlZ3r8SSyc0vh8iI7Xf70hjZ7+KYANMtN+z6mX4wZ
Yq/MGnRGv2dzs+flqLAZI3ZD8VJaAh9mvtWrBgpQZghr2IxppDh4aSrhru0QvWzgLrOfURa6y8Dh
1TE0+PPS99Z/Zb4YNlOxMIKpdj7SPJhs5AYrTNHUcYnuRVYkgTYWFEttn7X6phn/WD1asacG79gL
yhhU645dR+pYOPtc06M5ACsa1edkkuhpmlIL0l5O1aZgaOat7rakgDUFIAbTbUrhGLHGuP2Fj7wY
mDa8zjc5+B9uHY0AFdr4l2ZDZnqguH7AJ+9gY2as/g+dyaDfwbxLWgCR59KgU+cZkKhLc06WFYed
3Iv3VuDwDdRxvHs+0zprQdR61XwlZFG9xrHwH9nVHh047X78SQ1F7UdIW0xZf2IU5rfssrAxE+9n
XVYEQipkDbcXp1Np/ZZh/4ast9dGPX/jAXHtVSRsk2QoruPW6K5VuD79tFsDGlqXaeUHAa2SDPDH
CY+QVKYEGs9IHz15UevPjj/J94II8dD4szyymnNW/tWE2aNs7Qj3r2+usJ01TCG1BEnZzYUn/eDZ
f0XBeT8D8+ANFcuPRwmj60WGBioJVroRrOOfYl8EhmR/zHssWu0IBNG7cLYOMgKnPztfM9ywqQhu
d3+QL0FH+Cl3AmsM69rjRbP7IELRpmXim0zJZeIp9vbywPj6qcOj2gS+qowJU1hgpiopCa4bkaWC
Xyr++DY6Uj5yazaJWDf2VT73iAY9Wciyud60VNxX5pjS7LD9e1FYkML4kCo/h+okVDrcB6muMSLy
0w/ZpTc/NIK8iWyMw2QH7hxR/vkxBpl12D5W3ZCPHasLSw9wDVtKVp0lRO1QnBWUmLDH+UkXVkTo
aMqd5LEROepbM8QD7PraRDcLJ2acEMXLhCGHpH0tVGuoz1aiyXvY8uaVDxxIqadsnnvbmyRpQd8Z
3idNArVivQzJLaCGWQfZ0QJR2HE2qzcg1oPSYG+dS2Axd2xR5a+GF5QQWzoMy4Y0Hm6QmNR+D4Z5
sWCDyP/HcmNekh89NG2lbun52J/LrRdqYKep0twFdneQoqHaIc10roNcZwtcaog7OaPlleYQKS01
yNNwYujFgHHHjcO6ZT3jIJH6iDF+W0v522oCM7KqD5jR5IK6eh8rFL2gN1GqrPvECc8hDXEFp7MI
zoGRrHUQqg96pl4knYrkKf6Xk7FuTRLpVj8E9J7fZL9yzBK4jlC6HHQ/sn5dFy+hyBgyxm4WIMQp
y9ymUtSEgGG4b8vKzvtrsg/d7qJz7D5CID+oMHOhE+ISAAI+qgIG0h32bh4FklMNGFKUIQDR7kHz
j8gE1S8cNAYledT7n39Bb8uXX2RGWh4jmBbJtpbCvVELb1/xnliK/NDF58ES1OCbuuJfqqEmf3qM
DdNRGFHk2aBgo68eJFvROTcYmAkl6BWIDzxd4HlxNL2pLf5+ONF3m1tr2uY+b+rP3EnBGmTo9kSh
nFkNkks/jPFgtQmdl1aWb0NMwMbz/elb1mnAunaMhFIwt4PUcSSooKlczciA5vfZ3jovBB5sSdiO
IC3T7POPGL3JrGvuPn5IQ+tKNffGK9sYfjbu7RZ2/3W7P6UXtU3Dzg1zTCfUNKEv/wKbCoOnVrm1
3daaZurjowFZgur+s1qdFOF7F5tK/eSgYPk2bIq0DHjMVZRBeEcoPVyZdAJGsV7RPr906gdBy2lK
t8NSnw4PyJsPDsNds1JisYgzmZ98nmOy51TN4orwujXoTPjpev/IFLDd8d2sk5KNpAiN8rz/CniR
DGFhV9Bqt3cn4VKQl2s3FVFnp4rmjEkCIvozbAknf4+s59VUScjIEjbwNxdEiDFd58zXCPb5xk8w
mIIQbCUmRtBVYMMZcpwjx8HP6NUL5I1lssag1IbcdTfKkfhnjZsNYsSNNyVhGgIrCSEuiauSNX/P
pPfh5Jw1deFPZLPZcMIMI5csiytInorzDRg+HQdNbCWH5DoGs9+NnoUqlvBz0dFr36nj9zCjAiT5
IT+FBB2874edIKhE/MmQ/rxItum58AdUy59nWbQhGkY2TS0TgD5eSp9/0ovrQKgi6DcRlqEBhHIR
qD60udkZwpDknkMYXDWJz+ajAbGeYfY9eynO+f3tg0zAAOsQGkma1OBGWxKeF4XwQux0TwCcXGIA
voL+QKRH7uyRegmyAqJ5hXQrvEN7/bwBgqwmXQAQEJJz80maVFzVPPOeDHGdJYdN/+xWPSupcGVr
J0vXEiZDN8LqqUdBzejELns9yXftx1jvgjAQA4vq60SpHJsc+Ns1plCEcKfkZQuATWIACsLtwCq8
cQARxnPYb0iXYfwzslrJdySda/FttwKhhF4Tls+SlCt1LYqxGmjLj+4NQdXImi+JK6jAWg4O12vL
la9Xy39rUvZWItUmwMTQ3+mE6iSe/vjyxec3yscJ75452qVinGh4cCBwn1kHkQ5BykcMxaezHXT9
KdrMg6wZkFzPOi8i9zdiJ0cxgQ6WXD84ICXMfESucpJsEa37eVnBo7C0GjuVMl+FnPYei6xk11tL
7sJ4OyNhmo3ic7/s88hX6Rl8BwN7NvoOaSfGphX1jjm4rR04F4Rm2QelXm3cCAVMNZNaBH31vFJd
NGy61/a7aIUX1Ju1Eied1RaOeI9StBDOb0kOxhH/98fC3QVA78wZS+my1FeQLLnXkuJrs/Lmpp31
7qgCGSkUyFuLCf8LnK1hEw45OAkXiLGDtWCbildyKQ5CVo9ryPNTiOpBl90hrE3ydEH3qaFD12TG
v/CgcQrp5zPA/RhWtwhI62q2uza27+BNKStBFSN6hsYoXnGM9ACqVIECh16Dsz/cXn8uBZA82YQj
za1MiMdlB9xVc9Z0ovkSWFvxvWeZyaDJSQo+ziOzeQ/uqRyHPc5Sedu5rthdL9pvWXZ+4t77tJhL
H0+Ou+GtY3XZM3JttN0MBmYHDknL/aOCzo/Ubf9TEQBZ1dHyL9lLvgAuLa2PoVMGMZDIV8GAKvs1
NMQlR9yaBmuwLSnTAdKrROHw90KyQjefClnMQTSz53xRpqXKmPmxDrxdtwNIrUDKNCX3H7dnnb4i
tq2iHYq16inxngN+0C66SINxMspdc644N0CXeLVMsX1zkgO4XaKNcogHix21tPrZxddSCxYIIdwL
v6Cg5x/bbx45WibkZxKjJrPMlS+TILLpDvYWVH1OzXCnfGPCf3Af+nBUXFB9Q6UZXsvQWJ/IpfM1
W4g2WXUiE1ojdSyZBC4X4jKl4lNJs7v9rP2dGiO7WnPs22fgcm8IwCRIOcvCliWiVm8gw8pD3tq9
MwlKGOHRtaZuot4NRNFF2hs8mTPSeszAADSiSbweRQHr1rNdrcGJgoldo5nIntnZKfza3WSckHL6
tIaPo9VuXaANIIZFM7akMk5ipyzTb0ySVHlvN1eEUMWN1cCrexB4tesNV6idHyckD9aQz2zXuFvy
TP2O1vDUudoiWB7eic4wJ11svCImYnHSiphpUFIKN3VssV40Xp7hNeUDnymBuHeFdDossJiT6KYu
rIQnz+HY6PinlhpFwg6/fZRF08B+5OXwmPyYMTuQS1zO6KI06es0uub/ITGwjbAMVAORLPIm8jvv
NQovr4tz7lgGZg7m7TBOT/4IatPGgRG7L4oo7HplN0GABuRVQoOCzWVXkiQ+L4sglX0PcEHx0FJS
YuRZYZuV8OqJsyC1SzpVtl82VfzLA8xguEM6KA9q+fqEHphRB5nfHqRrvNcooXJfutbBhtqUEuCN
fvsEBSYX0oy1qxfkQwvK4DHBIxFmrm/PKlKZbsPIgUHpenPopNWo95tgNhnbOgNq27htP+OPJV4n
WPQi+cs0FYCVa4GO7thtCkYFwqIt5zJou/GowuUshKHV3xXR4eyJTVdEgqK4ISO3Lb1VC5tC6+g5
XEW30lZBpAcxs6pizM8PlVOYc01eFBXmgYWdHfXhBQdvGlAqHOE3+LPdjBQMd46gxerSnd41GZ4n
mDt1U0UFzX7syli7+DT9erAXtGasCrgsWYoJzEdUtnGqF3/KtzdLm+EIVAIXX/P4I8cBz3s/h87c
lp1OfFlnGwXyccfEr6IgQvXw6hEOXxH4xlpAm0rTQ+TEGvrppzOIHEUIity+Su5h2fkebHT1SHQk
qaDjASngCgEbte2cbrZ+Ge7j6HfxM9xzufems3DOyHK0Jnc5aNZvLq5v1LlXhJYRmqiZH97Ln6ws
BZOVaGQDnDvXPTKoVh3VEHCjd9MemC+c1zeoSV7YG1qgus39379GWUUOt8g3s8XhD2sEAxSjTCTv
bNM35IHOGSrvwDiogSmPdydytmroEIJKkXcCjmS1YjCZ2WFKYB091nOCGhWz8WWaI6IqWqXA7PEg
A1p9O1nhB4Frlr+2bYuKSoKX/6BLzffLX1iZMucSQiYyEctGYQTXZqU/ae81hyaWjdBxDax/DQmC
XqolNSpb9EIoX++fN1jpDmj/f2Q8ECJITHfIoiI+ltw/u3C+nTpU43a21cE+/rV3bViRywcFPZCi
IL2q1XSYzgRNwVEqbZDNiayala8N9USE/ZPr8GjQmrK3vFYQbWU/PzZUHyAehFi29KD50KQxm7Lg
HgCogtFjsdp72e835HL2yOhFxPQlDtQhzW/6hzVGUaec/S7FsE6w6eg3+1qbBNCUAx+XWi6BglmR
hORmYoiSllUm5lSIVBfwswkSzg4PdrV39Ds1n6ikjJEXVybm7ZiEgExLW8TbUymz7c6A9FiQGasA
Cn5CwzDzzLdUGWq3tiZQ5qMPqTd1c4l8DPMZafPOZfEHMukhov/qEz3fjRQwYMhdolpAZiM6fWTN
X/ymrng1x9aYEBlr4PGZMeulQ5pxMB2oc8yaXOMKldFFI5YJUYJKCAdDhsYcww7Tn30lU/S3qNu7
VIUfXuX9Jk8JZ6rYVaj6QZBrJ7kS33wUb3yik4JIh87LvZ2Q4wGM17zbsBO8Mp4KI+Vl42Wu7LQg
VKxCiXVaGvvZiVgYdn3gPN1xeYyzTrQGqu6NnSUdAW/8vt5hUY78/fcCtKSz7KNHg2Y2KiJXWBTx
QQl2PuNtyt7uUsBxWnbcTJkDUzQy+t+d452l9sZZy9QM0GykdxvPN751qmxI0WXsOIr4+O5/dCuY
B7tZgeYy2a4zd88kQAI3xZZ6DmMovVMXtPiEXOrAfoYXuz3btqnwA7cSm9tiuDBJIzoG/dAUW+cz
n+eTCqDD5Bb5Y7wDUrv2X61foXS9XEGheR/waLBmx/5p+R0ayYopS6LIerPgkvrSTHETEI2k5k85
gzWLb2f91Yjc8E7/1PTfOMb4+GWM15ymQPLtOASv1x0Io561ER7EmTTJSAChsllc7kvChNswY9EO
AwDQpPx1d2YCrZsVZFsGjEY4Iixx0x12VvGjupuNL61yeTUvu5pmzYmMbk+fe87lHVIYuxi+ePHH
+dGU20yTAB0HQU5P6zQUo+BXliVvRFISmWH3KKDMcC5utc1IzC06Wfse6/2wEg76AIO7SPBPkkct
n2l7owzIv2Ag0smEtzx7I5Oj/jSWrUQ3+YoPQUSXqa+kH+wzgFw2nE6Sr0wc8eJ4Z91puAxUnjI2
IqWvHnPBibDelhGCapvbKwkydDc3YKA8c9OJiM/CvEdm1YrHf6jSXGyabE60u25mcCHd/UZUd394
0eHo1aham3KvZNPyvvDlJylaWgkb8IMPS3tt3gtnSRFRe7In6d4GkyScTQt4Zpzcr1b4OhpreaGo
Yeaah7wA3+yIG/XQXB+KTKoCwg1XtAiqh7cR6WieSspV6osgSYnMEJ/SlEASqQT9K3FtFIqKunD0
RU+zy8q3T3ZOIcKHSajZTfCkw1Jh1xPU15NSJpxMFva1WJlAhrh7/o40VTKBBG+UGAQ8av2JWLhH
uKZiO+AEDH9pCv7CcDEmDGk3D2MHivvQYXbJX3zxRRdBjVGJ5ThJPjp7mcFZQQugM9TYC3PfmRMr
U0pz4IvUFmLvmVSqs+p0tcK87E/Bl+AoyT1cgUH0mPavZlbQelZi/lnbN6ZRUAN8CepsMXlt2NN9
GQmXnWJXodLxd91JvRwBC+nDHdjWHk1IFo0iUCmtjHjCIjo3vasWuQXjpLMX5KmIyHwfgP+8e1l7
0mM4pCTtDg1JCvej556vNztPogbGq6RClO4S+tsWtDyfA9/epfliHcfNAdpo5rla+/OjhUWp7CQC
bBz0XKr6VkVafiL9/oceRchCXOgjpGB8YYLi5HVqln4ALtjXyK7+ZP88enYgugFM3h0Fc7XRFJdb
lHMtoqI7wi3rqk75qyCmZh9DSwB8MtDO1JaYb8E33xQZyWsIkvsqJNH1IFixwRKZg9XJVx9mUayx
4fo+DC4JfgEklthqkDgsfZXrqFThOl7vYJcNnriEvIyIywgnrSbFAKE3X0gyy+unUM9V06W9iEOe
jLKkurfv59vbtBVCOIn3MQp6rVdjoy7caBX4zVLwOlNVnAgNLZaxmpLG1F6MdoPEw4fMJPQIS6DV
0CLfYqdXIzTCnEPsWW/Tn996xfmQz+kWxRp++S6LMkR2nzbXdbJcqobEUUNqh9x/aPrc2yUCSMrt
4q9dO499Tf+UA1o2VhghA7U3jX67eiymYFa8NS+T9N2xMutsWsd7dIjlne4kuBEkOOryu/AbOXho
QHbJ6G4rV5G6gPS3nmYe2GWSi99gsYDJ/Q0pBjSFDJqV1o3J8yppjmNgqjVvjoCGlk04ND+Q9+Yg
v/bnNoTH0VPd7tBrbnSLioCwoW61//aox4x8S9O3gFJqzr87+Ky90dakFgmFX4ISZPyVqtqR+o1G
1HKBRaT9aZx3hp3wcPfo7iRcaTMOkbXTMWYXLKk5WxR6rj9Sd6UTAAgfJYG5SOyVoUX5yW8pINK5
0EkLms6t08pjV58hQcq34yysSDLReVEvZTOmUSkOjgQBJ4P28RKHYEcSlB1Ds+qrgP1YoA2/r/vU
sGUu2DhpX5BVBq6yzDVQ+Ds/UxQYOKYkgR4xS1HKTJrPtn7uOcYmtJqtLsmJhmH9joI0DE+jOdGN
7OuS7iayq5YLBleeN9BIgFACSpySSuV8D0e5Yc0b1XNno7NmfcXP/Io07l7sc2SeQgaVydKfLi5K
Sdz0d99P62LPDnpn0FRrWsJiVbFu7O+Z5WrAvAo1M+eZmlUEGgSfnihfniW70QwelVaMgnBGpIFC
KWHoVBNzN1SfSkIJon5OQEtx8qOkQu1i6nGY1gX89EZENQNIb8Jbqmw8MMO3MLNW3H7cLuATwuqB
n/Qu6jNU3vQY2fB8YcG1wzrmTBBTgdVO/i33qc99ROYzCayqIuKXKhu9B7J7zw3BBaf6oCbztSZH
CNuZC71OYEBS++uzOCe8cfNHOkDqgwtvXGwJdPQpt+sksgV9lQ863TIX55/aeUjQeM1iDJMCjS0i
clzUIlIBAsNFXwfxM7OoGy0fjh0X2M6qFKB/uxzKwA2WTZ/lX6j+g/+kAVzjvkX3M+zztMOov42j
4tYzTw1u944Uil9+/y3qkHg/3NTtQd7JD+e04SBzMCY45TnpN8xcy9+9iDMSpYgkcE5x0JLPqT+3
UCqR2mJwmMOQT2dEfEl8D6hfJWILAFXyuf9ZdIAdLlU/sJbwahm1rxcaHoo19/qrOipbrIbTGDG5
3PxfLgS+310rzIKvpCLThVrtWgCKaTvJHT6gBa2YZ7BVSxKFMwpkRwkZ4urqQvwx6i9JVscB6CBT
lJ9JEhC0lUzrzTrdBU+zQX+ISr2Ychlw5tfmYrORkB13ajFoXdxyaDRtqlNJmaPH3V7k564vPbtF
Lg22Ob2vSSGalQQhbgOWb0u+4SPpGl40PuNNO4gYkrucuKxm1SBN0WAJF2Em+wctsGfHRX1FzW/O
WnbMMuwIC3KvaqjdnxpmEopEgc9rD56FIqodBzu8HjgfEkc/bbxScjbwxow8TXcjtV89Mj0V1TG0
O49akQUL6rUPS6GocrJNCog+YWKuzAnA5HOi5Hyw4iyQdly+T33W1mw7qNbeVrzj26TJ1BdO4IeD
ObF6Hu4w25+c36qrvU5G6SwMD94bPsP55O4OVeOaqkEHS1ABPe8HJT3cMUv7s90DKDh93nNzxpnM
eQfXu1h5Z6xZWShQX1dPcIPrHto6ZCEAmyc8nyoT077b7NFNcABCmGbJR0dJ8331eejg2ikcbPs5
8PZjR4C4cpSY2oJ2uaMqQmyJas0/yYnFJgwpR+uigKDKyYMr443FBSmZPbttzu6/MkNUixSI/uad
7QDGPXX9TyZaqBOXuRhxMsEflexeyCqzZF5f3TAMu3kFKF2Xi1fm45Afz3v+q48WhfkAAI4yddQt
2G9FdXKs9M4DwBXS6PrD7a9m4aPS1qZ4Ajvyn0V/nOYrxy4hMdqW36bcREhZzqVGZjfS/MtvZvxn
zHkoG3tVYVVVWUrd9PlyFEIecCvVMWnw81zKWwjD4QYaOldfcbH+J2HQZCATHLLWCSIBVgPUiB3r
EZ0r1WsZFHvK0Fzxi5xWQwsvdbLpJYlZVGp4HD3bvXa40xC3Fd85Uu7It3vIJUOXNX1ur+i1R4l1
8mCY+z5R6O8hrB09VrAe0lPRPjBO/jMDALN6Wyh8JGUNBLQdcVOreSd8zXFL9ucV3/0of89F3XKa
AjDpVPTNj9r333SYpVUqYQaAcurvKcgf6q9MZKwCLU5do2El+ap4VvwXG911j7uub/onahQ76Jl8
aFYPgDf1Xqr/xlKah/bEIlh9PfwoohTSELb8vkLGUoDypxbry8wEDPmqBLHDbmE5Nj2VNbUzscAr
I7OfDxHmDbPKt3qwc5v2lOclEkaBgvLSXtx4ncLAd1iU65/eTvQOHlDa/+Jdio/YtGrqRuK3PeKh
y98iG6VGwy1cygjgWXGagCBFOfts7K3IqUOyz/y16pxlP5ZB7W1iJAaC/jv4XkWqUGGbAWjYruTD
5/Yb1YWIT5fdD1eswrIQpwRxrBRRjKmahqaTMzPikI4lPHY8atxItEpm81jAAqGu8T1P3uekQjVM
MllK+14gwJJZnbnkGRFmmgo1rbHG9+gNgbWJnuZ5YJbdebkqCv4xJ6yxC2yES5FWjZVs7g9YZu9b
encJ7oXOZ5QmYuE2iXXef7B9jb4oSPLpST4lTwlWG4gkX73ShYdiHcu3IJa88ZEgsS3HJKT63KV+
ceQbcEFlC56/U6C33ZWzaah+LoVMvu8JhObIKZNYF2I5FB2xlsw7HXHoDw7RjpnLxULYsy310tUr
9OWKOOxbL04kpY3epLmbqiOs229LKTUSfHgXVdnXdyK+brlgnbOpR5SSVG2+29Ilnh0cf0F0luDR
Aaj/eTWSDKV7ox4IzxFgsGKS6k8khsq18y0V3b7D0PNUSL5wkU6LDHhFtgd+YTSuBnyPKbw0O36f
UPEdBVW6Dzk7/jIOrdtnhgu0jYtpgV1mW6VPOUL5sKtY3wl/iXATDjZiFnUv5Zi0kaTgC4GEr7+M
FUfPSTL+vq/7IK3cRzgvFp7tEMdGARIFnP7BI0CEYEv24ZD6GlKcOeowLYW1UHOI/urwWy6SRXoI
9nqnMkfGjzjce8GBkJPcCXy80CWLMywme0y2UJ3AtNeg8fJYdtfkFLDckSLJYvAf1YYJH36psQPn
D/bF6cUZy0FlKpymouBU6CZM5x5bQHCh9BU/ua4e3xbEBrwJ2hi9MCFritTd/SB8NTi1ghdU3xRI
SUkBhI74pO/yMSGmsKJWCs3GvYgnivT++CxpJyOzdq0VBK/uLbgPRPH2R4xGkBm1jI4t2TKhsM6P
c+AUy77IwDVrHD9MzBtVKEjg4mn1PeE/SCXbIRiG2Jg0kslqXnOyDXQ/qniO7EPmgNQ1kQQT5MYm
3TiAWgPhlhggs9DeZqjnzqBxe+Xp+bdbNPwVjKIZmwhraIuCObhXZDg8utJH73sQuXE2LYmLrs1v
gbxS/lzHcH0me/7lGbXkK5GDYvNB6P7xJFy7ODPretItdGzO3DB96Cjq4di/kPcDgOqCOUn14r5A
rKEhri7WUTXcgciqysvQK7JY5uBjpPJgz+MsGRSZxP93mJgcplAxm5BuSiUie94bg77r6t2VbiOP
jpZIg33A6NAr48NTTB5DvkXwbRZZw3ftqFjPBTcCrSaR95P2VBgY9Z6j2UdrPskG/ES57zH7EftC
dI9gvngVppuv8R8AY+K0dVWuxEv5eLR1y/h6b17ebQk7LLa49kx6kK6mCpwuaxvQu4y42mMwTovq
BAhTRZ9+c7rM7s3Um7Vnah5HAPZ3azGMgIQSujKcef8MLxVGfnsqg8dEI8woP/JETs4NJB4AGn56
nfRQeWCX8t0o1GhZg7Ve+f0Ha9qzSirjZfSKAmSVghaZOXlw+5i8OQxywdLHm/8KIpT43/9y5vX1
SZqUAZkaA9ZD+G8H84q/XuxzDkSota/WMgpAkWWF3h/HBoBARSuFG0Ro3W/F8oQrstpmk09Y77wR
dwp09fZcZIgBd0daL9DzK7szLtEpX48l5p/Z71yOqnY6Hkdnl2WbPHGjsH80QGW5K9zTOv/9SBV6
oQEPwVGU7fsic/MNw3ml642NJfxUHhfjbY9xkvByhYt2kXYzdEFcWGUNL7lI6eockK5W7pZ0+DSF
7GL1JH+KVpU2NoqXqFM4s8JiiI5PezRpjGybYpiK6JF3r+MZ3FNHoM4Vfqi6zCfT+NMpnu7L3IhE
rDMPQJQhCVuIlgvly81asUX/19hpHfjSjFsANqxwyZRDZtiZpNHEvwaTIgkSbbMiiMWj6D+KA5RL
8+Ac7OvofeSDt7Od+uFInHXSGgtF7GSqw1JKrMjRgnTc+kvA0tZ9cebmCfAseIe870D7NO8C9G9F
w9hGnp9z5zvXgrwprXEHx1whCEPtSlMFpO2syTPkSZ8rwbX4c6g2XmF2M4XeazhJKUm/OQq/dioU
Q/7bCw4mZ0ZquolU8p/t/5vco2YTbDKzRzCytOtj8OiGKCgMnvtOYusQ1k9UhEQUPP8wwEg/yBSw
WBNm6F1P3gzfF3fQL6PRONjE8tVjXPvYZBXaeBz2kMoN45LfFIm6mSDJmHVOJGmbEz8OYcY9ROFz
OQhsUpnxLJD/yfR5cR0yp0CHa43q/y/tR2e9s/w92RaQSuXhBACqOTiD4YIg/6lJa9++I7KAZjS3
l4kdceN4x1ZzEpDHbGkcYZ9rS9XViio39NHCXaXuYrGaYLTXYiM6bIU+C7k/bsKuWrc6hzPz0hf0
ndcLG1ps4AF0ob5AcJ2sLxXn8Dj+eNxMSn7TxeHRM/KGVxXsa7KeipCR5SdvbDPchRG2qLgboJ3j
4/yBdmiaMMH3UE/ZaTdne37ib2Pro8ScLG4cCIIjSmuUTZQs6Cr9gCwEjQ/JCKN3LBTSP+tVk0Ij
Zqic6FJt7gIJO9hMu9pwXHRt2xbl7WSEfPKD4MZidfnK7s6N+fKESrCNZUlAEZ/rgEhMWWigs9k6
hRelcp7G+Sl701rqe1E1qDeu9T5t4UTdGFCBIFGk8RjEqVaQUOTnjaeH1e5JtXGaS4XkAtywNHmk
X5f+IMspJwCDO/wlt14Qezi05Cc99C7e8ySwMNRCb4Mi0heVnw5ele95DvkAqOeI1u/B2z9Troob
bsvr/cE7ZURuVW7nPpMPV9s2KI2l9bhP2tUJGSSUYQNQ7Vl33QEl3UFvrNZAdoYteu+PN+cgs37G
nywW12pdRqerCjj3z3wxzXhlRDmtR3QoqU3T8Ral1wp/DXvrhnZFSxiLanIEMpFbw7Pbq3T1QVo3
XK40CfQjDPhKvcaxmqDJdrOoav2PlcO7JKZZcgo6rtlF3/JsXKZdTbc8JV8z2dzTtzuQhiuqhGca
eIONlbDnMekiDt0czm+kdBbD9XEmtdfGCV9Ip6IWDi1Qo/gMEUQ1VCyCZKNlr1ffun61/pwVxwrj
pkZG5DuW9uSuZp8U31MYrYyuH2sp33WdPNspI0tWeYG5v3Grh4SF60Jj1nWZIbW4MD7g2tMwEiHz
YwkNLjZbo2/wn7HodG0lqrGKp/Ur34VUZ6yzrvBovuwSmAEFOzPUY89nr39YFL7eVwbEUlJLbEkC
npBuIMFB15YojgxeJWs2NzwTot8GTHnjgp9auy+811OlUz7Be7t956BfKkHgjGB50LZXYBNtsWMn
GMKHhi7LMwCr+bds3S5OnhRSiY1bkzaEekUXUXUfJnu1if2TobeDbNOTLW7K/bJXtHboTeocY9rX
XSiEs+DnRqHOX+e6oYodrfncfZ0rCrsm3hT+YjaMXrp3/0GpHp9clRCMfuHCMz5+n8O2ySDWxM04
sV/ytnw+pR3A9raXXRi/9bDgv9qSE2r3UlpOvHrQ3hXylCqG3RwEtmFEBz1pB9T3VS3RGu6MyJe1
OgFv1tBKxfebAbvg99IXBHx/AdIHJvBZW5Ki6dAxfcqtqBgfh37u8z4ZCQbV5TWVY5lbN8AVsGyR
0qsAypjCMiDDibnoknl17CQxaaz+hLRnzer9OzhM3PDRoVXHG5WEC4HZE5X5QJYpWTpyGpEe+D4G
PowvzlUlYXb3USFQaBzGY0yoripKsNuPklaupqIg0qvn9ZMD/EQOiuZuSBEi3SIdvbvgKannVWnS
rsSMVYKgY/RWm6BMYuXnT5I7JUJ7RgdbMIxdsH3B47DDJpjYasl8akgnze09T82UQFJoipTIeA4r
PIf+Shbi0lRE4ydf0G3QUP7fo+ZHmZMgEH8SfnQ+pEk9o+d9IhwZZflbZ/jC+q9NftFYZ9UK6UDR
JtfX7SEwQIl5pAdMEOteWefUNIf63Ovi3SW3xr3JiZ6KgkGDmNyxJDdrJl6EwcFsRVCz60evqvkx
VhVJcwkZYpvnTRRaekO41D45V3Lrxlb0ZkACZ+tNV3oaH2ub+uIc+r8eHrMyTGnKmarCZ4XB65KP
bFSEJxU3a9k8aCwZNvk9B/+KsLJz5Uqat2+mIzdCE/wzHDvTazV9iVf7dIgeAd2SYavn5Bao4MqQ
AIRnHSIz2jbfaqRxuzq3N7lDJ3/huFZ8MtvWduymrLpxDlhNglVmzGaxeb9Ap/vEeQ0rpfv+lJGL
Z1fXE/upKPJaAROb+xnFoPXWp+sbCLqO9Wg75N4NkWWOtAOEw/xr36PLVDuGp7zvKy5wDIeh2vKZ
mhGEHRQeOdEj+pIjGOEHRomDtuI/eT/3Vdz5OUs8E8UNBSn4ieWi4Nv1CbP4XY6EH499AwRBPpLP
cWgNBHmu2occcwnOA4T3/BxUPCEd6nzBLhmPEImFyqhslw5lUyvxyW0CFzQSk/XI3yV8hGHX2D4V
TQ1CZuUIbwWmVRAhOJnvsDiIhAGp+7z1SHWzVvwXtU891OxitmIDHy2Eka4kd8V5hvUQQswd6q/W
Y8cvEre27fAdDmdQLzH3fbhwWnDDBNNuHWe34so6RKZug2gBBtiLvCVuCB1gGi/dHRZGM0zkfxV1
7sClg10tfORRm1Mc3S2qy4dI6ARAdO+cK/XUMXDuqNFyOnLhi8AqHsNldWxpJd5XnvIPp4oG/Kit
CK4DKd2Ic1CcPUxf+2W6kM9iTLPwx7ihJfLo1lde3jveo8oeSSZ3SJ+jz9uRALZy0un3dcqIfJOh
drVRYcocZxFjPeC7vudbuBdWX4THz1nUTuojXaoPeuI3sQkHttaGxjGMmmZyk4XyzcEYqwc2rxiZ
eRob5XsnhEmlTYqao3aKVRnWD0Ids2EqOy5SgK2m82bwBQvQUqqwg6h0eQRmTztkUWmpN+NJgQMU
j6LUqE789NnViWRRBTzveJRBDWKwIQ+LFSXf75W5tUL/licqnFEOBIHLQDxcJZ6SLX1lt0m1uG4D
p3KMQhqPhPwSothsmW5/siE8YrL2bQurXMRrf9NOe2VMo13GbZR86witQ+5GxJEbBN64+LkefLP5
7YfKVl4e9+kcVMPqhZRlpEcyxZtA6X4xb4Yn6N2WlQvPWehL/JC+Vbdk6hByIIj4PAsivrIcrEdp
V5GhwlE081alhvRxFnJtPMS5mU0bWzaSpXGTXybFs9WJpZ9FdomAmeZiKYum6V+d4VxQU//k3652
cM0GjPVFZJ1MPkyXnunThx32VJJzZxFNpkVFMPW/ics+1yq0xytFfZn4ucCvNKda95qzSOsrXHUh
1lxn0XebtE6zfzfB0oF7di2RD9w10XL2kUcAYDqvYeKzTa9+9Qc+bGPEzQ14l1+KkoJTQdgD3N/1
a7zj+POm2SXHTuLHaEchil6XnIMudoT08efeorrBKZLBfiULiMSA5HK2DMLauEe4JeiEUGZ/6zHz
Nmxd4IdPhxHgP0/vqZmiDvkaiyN9TsjHNx2SJP8u8x7e2BRGcuo2LFgghYuH2VKSCLUs0fQEZGny
WkdZUDIRSy/NguXqtKI1Ygg0IQ4nybk2wljtNeSUdkhJS1tNPOmaa/sLsGFtL3jQDIeq2Q8sw5PF
tEUskZekeQAUe1fBIrcvzJ4wO6ff/PavobGfDcl+7sE8wFy1oxXzwDesQpUZZfzctC2A9qs3ilz/
c1aj6yTzwDEgcjQmdFVayxEU2iU7zYeBBd/LlDvVgu8Li1e6cVsY5ihkZnfyk0Jt287QcQQJcapn
J+GXFhtwuXQVLOuyhBjENpc44jiXuZ5J/u3zNBUy4bn8M9ZXd6T1aJ7cxhpKCHEiL3sh0RlcZh0H
sdjpeVd9js/UhKiaQaActzspr/x25393LDmm6oHviDEdNK/twpnKtEn1OP7TXx5EXyPWvPQR3VOk
zFv0ynvQFXGqhHVvDj0ssAFLdDl/8WS0lG13xh70LWHTszCP6atZDkjSC4cU5RzhT9DbB+vXEPmM
IczHNio+zuqKuTHJtGjX2xHaoropM18zQT6LqdfvPfRyMKmrYC/aayiYKU+XBf7VpD4ayY6o3wj4
oV7fW1X+7HFgFCNom7cdFeoiZ+qWYSCRkYOTPSNLfbCOSPVoSBVAzgpmpPpP9JnVc6wK8f57OzI/
3MtZf4VD24BKS14X/ygJ3r+fX1BpJfadOD8kqjD56ApTp2sg9iKt01d4K5mqrEDIr6y/AfhAVEDJ
nGZkhy9aQ2nR8NgcidTkomW3bAAVSiIFMfplq9EAYQamdIkBXlenFeDMMy/H/dVs+mM96mwds5Fc
hoAqxvMKFkTDRZglLTyWBq9dbc+6/uLZQEJ4/9t95lraeRi+xqAAKnx8u9Pk9XfVSwFrh2UL2jKk
jRPbauNAR6naHhyfgztEJzji7QG4Ly94q9yq03JLwxITasweMD3skama3CKH5VDRAibLRXrMtD6L
FAv2LKy2aMnUV+OfOAKHggugXkhMKeRFjdT0uVyegXo6A3kwavgRF3pRBxIvg7o1deNUC0iAVVLu
vinfek27Cy9JL6Wrw2CNq+vHvew96rGtY2kMrBPRoJ8ZIbfJhqIRtsbBYSdZiQANvf97hth680Pm
cb9EoZbyOYcRKC8IN7zso5wXuFiqZEIwUqJ7PAcTCnXMOEACdt5KOOcMb7yQDOP4lRpGEqByjMrw
unpWShbka4xH37WDI4H3RPL31C5Jsmar8+VupAM6pb7cPgK2y/PoQ6LCb5cNFcE227LLDE8i44L1
yPiuhQw/Ee9VK7zzguYf5+CqnEd11D3AzvxJFaPqmbcP1xxxAMdYLESYerWFaw7bp+jHh+UbMuUp
1RJ6D8w908HV6Ui96CvzXKsBF8NRBQ1dxmHiQPRfcLARDYOENFmErMW2+fzwlwvpOsR5nHqdtsej
C3Uygu8dwQeJrZfUZZ6tnOTohm4OC9Me4H/oi2lRtb9sTtMBE4vYev0FUbkpu0+63wNwWpjfojhZ
h+lAN3G92/9hVHjXTFxwB0ZWMKYTtmrXepTp3sy5y1TNbaXYPc7YQ3zfhf8auH2FC1mA5AXg/vIN
+3lJ0YKj5GE0v8RvWctp6zauN401CvWkZZRw0DIWqHnM/zu5SYLO/xEkyYLm2/ZGVokbAPYTQvQh
VbU83w/93B/2fZ20bRP7yaC4WZmjF4pACb8YQdxKAzjxeN/HvE4MOuLHZU7lqWZOwgJ0J5Zp+JdE
pT1tlAo007aBLb7B7V81+pIe2C1Oi6JJEspengYXrziRy0DBpRPJrl+ZxOc/jUU6EXcEwmWHz4ik
a3UhBNEeWOHyw75lN+z6kus1w7pOW8zscWm0tmwAJWT5uI2Aqbkf+0LilFGSD2NtChx1zynzZIgz
QvEcYB/Zo1JSQdZnuf5HDc6OswwvTenvj7nPPN/eu9O1YFWlolNPZQzHQ70hz2NV40/S+SuLk7BM
t5auSAkaotve0ci/9A6C/6zi13pClk0lwJm55lPvFgNJp6EgcFH0SBTl4tadH/GRGoPQQcXodTTw
ghkHZGVBVmSCBxA6+e2FfnWw239MYYPW1zuszJxmrrBO1oaccUWigzewOnDxGGTGwwraDlZCWcue
laKYX+iwUC+WPUpIyLvNC6YeVnHLjlbFUUsoAEJle4II/WgmAj5mMssegDxnrOGUGtu9tB6a87Rn
93k+ODD3iFZ149g4rw4YjUhkAOmiZAWWsFWbf9qdjDMcu460IsIa+NwrkKgVTKBWetcvm7ra0RsW
sYiyE0wIjjCZFhpxp0okLwxaxZaBZx6fo6bAaoUjDeztQSvMw5p29megzn2E9CiQZOfxT7S7x1KF
CzYsAg4mu5GMYLakgLAorlX9m+hPcRqrEbK/ggkGaovtmbRsWbB9kvYRvseQ9Zj6AZbaKBsayu67
/opr8aNo9iTpihfuyTsqq1+l8xWbrKG43pNw94E/DVmCUB3K1ii17S8rQnenfDv+u6aFPOkZK89P
f8QQ/LaAaOfxqRv1KkE/4rMlQPuNvCo3s7LO0l97+dWF33ErKd5X3N6wOwWSp8OmnrkmwSnYRPhw
DJyu8+Rwaq7B1JcDdXEFx1Kdgvy0iS+N6LugD1NS0Sl8zAX7/PYRjpxGTnzY6ykqH3ykaWQl2YdE
iT0uKi81T4HGHQI9NXisAaPVfJH7MINhoEYaWcZbSxZmzBk76045tThzeyfd0wQwCvMOcn2z1/ED
G5anSNz6fSNZrROVd99UNGTRYO7WSC3kHKuGnBU8PGosv9opbyau/ZSe32aYWDpecqvxH85kXaCR
Xqchx07B/XEbr9ZsX6J21WBLxRjETLkM8zHD372Rf+6WPnY3bvHwXTXCRhnXDNVX8yapAXPbQa2W
JfDtwOmhEHkyJ5BslteYmmoNO4OgIgt0H2x2NmFZCDq3rbfJh3jYlbjhMrSS30Q3XJqxZUxNJ6Sc
murN6pX1WdbA67RH4J4gySUyut0XMCma+9k5eb0jDKL5iFJo0wJfyvRi2DLIXudDOSMyNwrn//Lx
OSvlRx5zaDXooR+0jarQI9I3RPxtS4FrfxygwPiqNx5YTvuLQ1R+N6LOhuWW6ZzSBUTlV1EIPh9q
7Gy5UDD6FZC1zMhbW92bJOUWAcysHshLRp5S3Mr0KqY3prReFo0USAO5qDyLh/gVQwTfMJk/24Wz
VA6QV85q7QfzNZsj8JZyRObVg43mwOhgFlc447oN6pKP5A6tpLvIF9Yxt5AsGlFTpzU+aNTepbBG
TJt5ILE0MLaleCoBTnE6sKHL0JSou2sq18W9/NNKzYn3e1guDU/SijUxecObPQYc9fcjEfeGNILm
OvwA+iFU31HvLX1TroFPG4ccAkcw2vvZ2V6K2ziXSh8vPpd+4tIo/uCKcGfDgh167TP9APjcqPxo
umwJf7ed7SJuhFwtd9qFU8AaErqoLhSJHZZPJppIJhIepXxQXuSKTLot8KLUAiaJLncp+/8/qKGv
c2wUZQ/OqTrx9G5ykRG5OpwKb7Ksvc7xBw/qWA1c0sCAvY3CwBR/fcqXm+JnJxRdvf2fVUGR7nZN
qAJAJ0WW2hm9rrgtLK2MKukplNULXbsHtUtwgMTcb/hhKHHsw+HytFvbtcNje89WPRZcabnWPoQ0
hAH2ZbbXs9IvyAG39v7ySQp4S+IBoj+OI4usCoaZsFhJQGhtSMjLqIEAxXiuMl9u1CRxXhoIalVn
OqWi4rZEy5GjKOEZ+pbV377IKvxcWOCIy0ojCbW/GnWDKA8Gdrma9QtTAQG9IyV+UncsH3PVP2bS
2yWG0lCnGw0FaUaKxNJhhaiukhNlpcvYdIo99HkrMgYJ5c+68O9ldNeHINKy/Gd0Oeg269BSkXI8
/tVvEL3OrV2PEXtqF0NYtne0Ira4Bdah3dHV3JGHWwx7pXu//QYW/3DYjUQGawZUAuBmZEBZ17JZ
Wtv3ZOK6VPfu4tzyyRqVxB9o03GZH+87bOKJQfsJ6w5ScZw1X0umrKA7OYdYesjeTPDz1QQYwLMl
IXVxq7FLs6ymm6Ure845cC8yOL9hp8eUNE4IjJfYMTarORUejgfTm2Nq92zOarDFsoRmW9YvB8Wn
T2jJE9EcJA3xr4p+Rk7vga3vI79L2E4CikXPn4j6md0t65d6gmuipRmr1ZmkrgpS9Wx8tW8ykwbV
l667V3D8MFHF1MPPYfjxkcwET/9UcHgpWdyq5wisaEgwvDNzB8yBU7UJIj1Q/mfAbU+C+XDM5YD7
hRU4kf5TSBjt5OP9T+72PdS3RQVvURttCgN8nnnhrzgz8RZlXJgQN7aIShjUL0SxO/TTfPr3Mr4m
ID18Hm4IkLWvdFtCKqVVZMws2cQE58lK4YOHMsaSoZEAAgFczpUG8g2MY4JtLRLjtNr+35RnOTmU
h95dUPgYqABC4kqTmJwVD8/Gfl77UEhRXjkgU/OXGe7S3tjFGdaFXS6l4V+YiSmcsI8dpcCFtnmE
NpFtxuMwky9gIa5fZA3gBZ+hubAwji4BZlQ3zXjM+qJ6vTln7qPR5MPGXRgzoIG+fGxtRgS2E5Qf
8GtEYjI5yoDOwkA7Fgxu4qG5Lqs9yifdauSr63p5eInt+gd8oK4+KD3FGJgNlnuOC66DPzXdoApA
eFvp7EQ9B50n2TM7ISRvIcURpq0Yf9KEdNPrgm+fQI51oS/7saVME+uGCGnj27tVd6YYrA56fHUh
0Io7yJNMvAqc7SmT77kigcBS5tc3fpzH/xMZzxr9o9MR91WNYTY8oqVXCeYKn72fFtoNsTd1nJMq
E7Lh+Yduiq07aVvhfIJvXAdcQTxvw0PZZRJuqiZR1UaJaf4KyLHB4H+ZwUmd1haANqswqB7Ydxce
nRMNDwifVRKHMFc8BsxGg+FRX5fEn1SjLnn7mOIcPdGFgv4/9SPouHsFrbOF8rtFQ41L2dRVkLe5
GKrpH4MhQ89ncbhoLYrrxxWYLyDnBaSatypZzUSrBPPbC3dxhRt73eqQQ/9xARek/qpMd8CbkDsj
V5yH44ytE2BCXWEKnrj4LygHe8a4wRm0sjNqi0DcSlUvDWsPqDeqHCT2DkzILttzklpSf/piUiFE
WJJ6SmPtUb5YBrcHpTfgCTGBRUurZZkO1Cs6nTTJpax8M6TMMkU+KbMdmJX8W/IJTIGeg4kq71vx
Ch0+u3/YKPMR1c2WMPj6qduvnqUobkWucyT4v950QaVsjCpPj2BxtbmP7wGJ5SKOh/Bf6WumN5eJ
KGJ4+E5RdUAYBPMoNWDWAAjjkhIksFtt2vOk6XmU/dL6S2mKvQl5VFhm7Ah6yovIy1R0NaOea9gU
aUCKm89Y1EQO9nbJi10bMXEMOxiQQr6m40Y5VBhvMyBrZPVMZVFkN1RuPzbtVuIUCwIr13CZSjfA
+vmAiuC8ltSBZXHA4xbQ9R+XJhPXF0Z6NRPQzbSSxSxsiTE5V0sVE+4iEOeQHb2INd5Sf474RyUF
6u0gYLsMcpUqrkeuCPcMS/7T2fZoNi8A6iWa7skMogFst5EOayoyvun14ufB4qpeRY1UJGwTm/My
ziYk/f8dKsa9Tbk/Vkul8WA8VZ+2TG623z7rlJv22llmx47bcsY455puXRQtu13RQx4DN5ByUd+J
n17pAwoTZ6pU0ibp8mgSENH92uLNPdxnEswVMra7AX+fMR2zfpFptJqVQq2Uk+kO9PF4LmNPDHJY
Zyk7F1cWE8uBaNc+Hre/2h4nGgrqssGJWuWAHrsut7dest30toqDiJxXXRQ9TRxfKefv/cJvItas
E7jbfqMuy/2q4aFru3yquV//Ihm+WorS8C8zoZFUpaq7xkgtz6HCia5s/URyD8zCqXa8oBM9vrZV
ry6RqlyrAaMvL+pdvFdQBtDrolthJqOu6TN7daSztG3g64QDaTgIq/z0rK/1qj8fa+d+XHDfxM8g
vZZRlkFIrNGWG2iI4gQ5DcBdZi+pfftld6Ezrf28BDXfj9qDKCj6pnESNnLTkks29df0iXFB/tMy
ibmtnKd/fyNHG3FD7ThZq2yJZ6ttArN8Pxpq0RANFHQBzEiOG+loPbWOToqTRS9xpGv7wWCM9Ri0
QJAu8P1CFChO0rRabNq8QBMOz1tcwmi4NttY0mjBLzlLx3Ha5xmC4cN3zTP79qqNWmU8P3L1Z8hE
wgGwufQWwb6WJoVLm/+VYNOXgn5W1pzYI3foOwIkipMHc4hf3WyKVk8yfGU5PkZL0kyGPAiC/vdV
y3IGXCKRy7ciC791OTsqGZN3OhIdBL4CARCIUg9y4F1ZMrwTeEawQSAc863Y0H2TLEuKoXDKLXnO
+0L4ga3en8j0YD3vuqtDPRln2hFCnGs1x2fxVlPr5KW4ycyoTDb8Yjn+UU8RVEulZ1T5s6mnili7
T2+ql64jhV0sMtxTSDNMCnlWs5kFCumMaf07lJQJ3VSme7y7s1kKvmucNDWxf5Mrdzk0V4OuPzNk
c2X8KGBo71sE2KBIbdnwgvlrxGjNRYXolPA1FXGmBth8JE7vdqIhGJimRPHx/qIr7Ozs4el2tR4k
vo9iLepkMV2H0Z61hzrIg1aEFDNZ3UnkDbZ7+0FKBvXp4z8s9C+bxrsk/f47d0i4zT3w/MvlK9tN
MmFh4xaGzl9MKD5z9K977CCXpjJ/dVAPVB9k+URplmV1bX8xmabI3rpn2vjFMdc/ivtcxqYE1Qsd
XjWCV8LqXR0TcapEy631akIfAjX3m2nZAVwRJahlrfJHs7Fodz+zewGpd0hibiEO9Xy1xbErE1oz
wU54Izd6vdGcb2VJGg2THj3Z+Mdqas3yCJAfA9FR6K25+CFu20IYJtUPCeLmmdndIRr7cFRbnP9+
7WJDMIBCiksNn40x0Q0XI5LwvXvJu+0WyHdgrfhLAGsCgnUAPKAWpDAYQHaV/Ua1bkpbUIfO4XSr
fwRFnDoJks59bLkQUmxAyGtHBmc29R5vN8QGpha2P7Wjcq6HUE1X1nofRNkDC9O237Z98vm8TsBy
Oe5zkDDLaV7lpqMAP6Jiirhdj5c1yzzaNksv/LM4e4Zg7OrdJ5Is85dBXYUVup5xUY43+TAwn16o
zAgTyHyE/6q2Fs4LEz+PtPRg+igo1QwKWCL7kPPoSOCqHKkAENG6Z8vfU3+Y5kp70iVSEAFzM52M
mUaX9JRAnuB7gQSbZyvZkg4vrVbm1Ap2G5ApLSzsNLZ3N3XS+LYDfKbz0qMHjQSC4r1/lwwmHgSq
Q8ITc3ZrFwD/YalgPdvq0AymrNvgHxiNMNxSsPC3svJ30LSx7s17BXo4mEwORhhrt1+GdQ3uqS1Z
wYtvJm7GPSS+zZbzm/FmyLbERUC4MOvcxnoMaOrRhJ/HEdgJuVS+lHwiyA1c/Rqp6Qha3YMzuhsE
Bdhor2QhyUlsT0y7iGdV70d5gse6kNeOERqe7ksNAGw9WAANM4mfr1hVqBnQSIhRwQc1GRQNFH0u
euUJlg6+CdxDQPkN0K61hZW7QhgWUkjAmTSd7W68axJ9xAXTXmNtMgKXfAu2KYMGqHOToRgCxx+Y
JvCZ4mVJ8002w6g7S9XUjVdFKCqcspMmfhRts3hsfAzSXacO/q4tEVmA4fb1GR7fPaBIFJGjuS6A
/ztdQ55Dr2VtJKt8TDQngYMcdi8d92xjB/2YgQtk0uL+09bzO5RP0nvwNriA6s/XvnZjCY2rJtMF
UhQXxnFpMjUKGQPPAm/wGavLljdPnwAklODCqYqEELohcOd55Yu7zbYT6TYMcGY5dquaIljhHfnZ
ulE7Ci+iUMg5KMlQ3WEGKkaHJDKSyAmbFWwvwUfq+3F0GdrC/IdOltT7eIq4yw8Szi0wy42Au8ZW
cKusFieTG4ViGKqH2J7VDdUkMrJk5tksgREFy1dOEcCfOfZnRj3Lc4vV3bqGhy3B9gVD9wqx6uC8
/4Oj2r71JcBaDOs0vJvObN3fw0HC6EIFisKoYJqol0bRzkg/6zYh0gr/yeUNVPgZEXCB1HguxuOh
GWN0iXQEKQrSqNVAP1e3BTXSntPtfrBV/IxCFWImMa1tpqIKEa87Ry4F46xWEJIueIaSo1StRISq
n4M2CtZmswh4Gg54FBq7tJfVd6I2n5zepdEwUJdBDJL+OqtpAgXZVf7Idn2RPqipJ+pFt0SPrBTV
tUvhETfYUiiCokqhAU88+e6/evGPhdT1A111MrDKPkGnVxVL+0+ZnqtS40nyj7SbZvIQ9bJChf83
J8dcGf8y09iH6NGKL8rM1CEjg87ImIkkFl1iMu8iyxUkN31vacy+Cq4/cwcWq5GxWd1AMpmu1yX0
IVgBQkDYsL21RsMms4X+8jhNA49KEVzx5mLgch7u1VYPHr/81kaau8Q/7WrB0dsXHQSIfQSUrCxK
ekpXNsY1bh0E8HOJRTGkmlYgbM1KBhYQ8HwuH/pbRp0YPW9QEg+2TqLAV1zD7yPUKAzomr3DbH/l
SwK+FqMU9mxSI2FOKhGJck7iVK7x6SzaGoGsXzNBY1RT/sumyBf/rkk08JE1ezXrsoRjlOBveXJy
/Dcur9x6cF8aEdZNsZdHbOWuBWj3+Yu5iAwF0BMhnqm3fJKFBJswhH5pUk4ceRPzcobFl0TSWqIq
yx+GbBnd0qkmirS++26inBnMVX2vdnQPA3DHgUSnfQbZcpVLyxi1P5I80KCaLKNmdDjKq5MWwFUo
auwZvTAcIQbaZLpTY9mdJUgU/r9qiGYqNINxTNXxxwp4W7JlxXRLZSPqjlznv5IoBLruXGEOkL2i
wxd9Wq6EamfOgoFHa6yvQ32kDYfcu7BQouKwIgnSSfA8H4W2R18SFi1Xq523Jp23m3HmnC0pC3S6
cjFuBHle0xeKa6w4jGloL2N98mCUzv0dg5mw6tIzak/GoFDLu+8v6t1ATTyci/Sh2zz64IlHe7n1
ntAe/oKQjYmScTSylUgvbolqiAI4SCAXk5a32s7rZgmcgpgD8+WH+F9hNduSm2etePlAJDlf7Dst
rShK5fDJG5unHMBkQhzz7XlCPjw1XrjuANwe1CqPXhDhboB5aWFd7lBlGQzacfkZwNukwrFMWgUn
b0euU5waSpVINNHhFQGwjBinpGRD3IkFuZY9/kcm6P7BFSxLxm70HYQZIw79iRmsTiLT+y1vMBXQ
k9hfKzfbZP2+EN3juMutq67KiSgRpEUceYOPjpuUYdj9mMtvsPVlp7SSfzL2Kluh0hv2WuaqDsAQ
9c3jBHK5Uthm+y+lX0aDkz7pClfIFjRKZO16pCCyu09WL2PALaPFpTdi9hzAxuG05wsyiL3VtAt2
WY8brnppjLLhle83LKf3p4oWzVAtTtw6p4QoSnQvx/5STV2b8eJZPjQyLlBibSpZvOuk3a6miUjV
5kmjDsN9GuafgNuMzm8eD5mg4RUhCDjqZcbTBohw6AIBv5mhBtRud/yWpWu2woEiqdEDcfxuQsDj
FHnnFFUTOFYV3y42BS8JNHf/BGXz4TlVaCkud9CxJPl2eu48rW4Oo2CyUOrAQePsokdoZ0OG/K5K
RaiEQx2XZ0DXynVmA/m0e3XaV5myfGvwgqRMfu0gXTa3Kp+W2hlLm+w9gIvcOPwfiw6sdqpPaUFW
J31r20oE/YOnwnNglaL+rXdtdrv6uxp4Cl0rUWJTulY53bgvL5miXW7ap2oTf7p7diagBkoTi3G4
IqVEfIPK1TYXZjiHYNiU9zlQw6YtES3P61DER0815gr+w5vcNhGPpp58DYPcKilmfT0fO9asjlcC
llJotYviqEDGKD2W1dFHRLkWVIMpGQl7jY1BBFsOLSsrWFhEQgte2xRL6ZzJTXgN9HdNe5Gx4L/X
+C8X8z7NRBLPVJ34rlTWoO9rhVJgwtsu2/TwXkXE2wTuQyigogkFd1xoANScHTNRVrL+ovpCBTbj
2VeZ8XppyXtrVhw+Q9OuK1MiKX1Y1bbueauTi/1qZ3zTpCAP75mHePFVOvvvJula+Fs6VIDy6VG2
9QIs1IDdxD5tYyHsMq7e9ZBRz6RV9subhO8gzBkK7/YHudOnZDiv0Ljg92fNn/21rKgukCDyirwr
+qLkQRuL1EsCl+BdfzOhTTLR+ftFefubjtUH1tg+Ve4p4BznR2TJbaOXdRtkdjZtOIr5cY6Ld9HT
5lvt062I6V0yVGpomojZYwlg/Iki/Z6l7vMBdXvS6i2w1/QZmG7mwYpAlPE1I9/zPyYn1dTJa0HT
pV0PneuOJ9In/ga12Qg3j4YTo4UjpuSmX5rmoPI7koFyG9sTe6X9F2eU24cwUyGWV9J8y0eDx/aU
9HEtNPHOGkYonbu95bSd36Ct/e6+v5g9VbhQkWxm9VlXy0+xf62K9Z+r6jPGrn2azQmMuzJi14Cv
kgM+k6yKQGS1yiIw7tJ86bPYfMAxsgI3PmkSKVG1tKBpi4psOoSMgscLLhmosj13HvC398V0p4m3
exoEhuJ3NwuY3zwVneB8EOV5yeL0tUUVfBhrDRRAY/RogLQGfTvKGuP5lwlMEptEMUEru8fam9I8
kipeEnYFmnR/wx380VkGL00jt3QkMbOlsXtePlv38TxcHHFpskzYp2RdA6wRxq885VTDMtljOSi3
SAQyhmdhetdvjF/r43oB2z3pGrBxgZR6j77lqE7UK8Z1PfZxVLdz7zNt7G8rsoipiL9w6tkCp1L3
o3Sj/o7E8jkmDY6wHg4gngthsP59QEHg7wf/cM3521dzyOoGpcs65Bzlz1YTf0yrmb1mCU1vOslS
Zqntj/SJOxiDaVJ8FrpfbbPkjS6yKAggFXivXMfHD+3biqO2Ar6twcjD7zEfEnQkc7Q0ZxAS1sEe
oQTPpsYvJcspFoZ3P1RwxE5TTCF7spjzgQbdu/wrHejo5iqX2F0XmiK/aiIqvTjkn7OKS7j2fMAk
FdnVpSpPC8IxZ9hXZPp8FPB+PMum+mRYCHqO/44RBgJi54a9ui22msrPDJ/NFAeB8UndcNuxwqt3
MR/7x8el/5mezUkr9pXoCLjLjSz4DssqP0ZUtUNingKYcGim5ckx7gPWAMzHOiqXyUsRTqV2mbLL
DiLN9gVvnuB6ZMJSDrHeWLTdu4hkHqnVkf9ApVDFEg8UgkWYhJK4rBMipo+ORk5G+G5o1ZSxPfHE
ksnYsL72WLE3P8ok+ro+1ukkw3TqEvTf9vBIHe7CTDvKpnuaYj5fRcaLZrKibJunLx/RLP+PwYoP
Hr0a5XpQUoUR94ZYOuBK62gq1qPFg2FOGYBB0DhK2Ls58Vh9SathgOYM8pCzWd5L45LU7phadivr
NMbJMahNFvmIAziGQWZJb293Cm0+WS5h6Z9PfpVMOjPNL9LI+sLzBAexRTtjhU5zJ6a/+AxoJAr+
y91anZ9XqaiGh2QiiUH9EODDt5eHkc67mp5XJ3sDDIlTGV2ZtjKDV4yMnkPx1/jz4hgY3RTBdkjM
ZvFTO2NMOxNSL4h4vK9Q9YsN7t6dzIXkwv5PKvw0xdwOLYFoLE8MzXiP6/oSzOoPD60TF7U2518Z
UhcSwvGZactnDfQrGi/gFupb0VBlGkzjATsyYO514+CcQ/1KvHQ89t+Fa/B1WVNdrO9HU+SaDoZs
y6MtvW/S+ENXxY2W9dhl4l2TDoRoaCciU5xZ/LeJB/H2fqs4y3gEjTTDqnnU5ccuElHUhk4Csioy
LTmyScGNl+Q/wAPs8nG33ee6e7QTO2H5VYQG+HgU4V6JSd4WKE2R3vs3/JAiAZIFMBZvyYMvcZed
40QKrcWp6k/rNGM+7p291DZf3MQ2x3vg2890aGnL9VvvKFrJKIwPHSmZ6CnIQusdWZjFkxGq3D7/
UnxMl81dIFhIMJDXTXtaqmw4iV1IGy0VhBC8OrMUnWMPiMzZ4R7Sr/NjYfGSxexQIIOP3gJ27BW9
vEOZVPXLyy5obQh1Q955ZbUIvyk9x61R8vNNu3mPTtvpJ5i0AnE+7oUJEQJdYwMPqXezT0R46uxa
7I+35tFRSy1bEdlqmzFe72pyQifpJlGzjXOwPO+rz3Eq9Ms6M82YbCM7DhudTvZUhSGX9iqrrMWa
3ws/4BdCRnveQgc1JP7tWPAD5mgvrlbEGfdEJ11LerCw7ZOzOp6E1e828fEpTQ6C97L0pfcehPve
2QXSJBBDcre/KTbbflKBFkAFrlQIM10AP11mY7CzK2BfX0OdOA03lRjDbZ1W1Rfi4osoJx8qWRHe
ae4ZWu2h8MS/LppKsA9SXWyl0u36moZONS+guCbj/BVl2FiZISJ+eaon6BGYeaEkuUxKK4z2K2/7
+xP79v0PnCyWB/edUIZCVP9aeXazNrHsm0TQW0YA0jyNU/F2pd7FqklKrosP/w+OUE3wlvqz1ngE
GQy++yfWNyVfgvK8YUtohvQCmgidTZ3PvZbtSWEXja5DW5Bbrhg8yX82Xc26p0vRli5YMHe7CuKO
hc0yKytfADJjaGcz+1eL9ZuerXMCma1p1dPKItYADuh7IBwLMtaJHmM+9WKHKv8Tsy0Fo7LLTfYn
QKxocrWURthlARuSQ8fbYVhY74dJbfwYGLEu29w28ZhmkXRFSiur018oF5SpgmINy0WifaTEMfwp
Zu3TrszHwBAvYos5aFMGF5m860dUweFX5f/+I/434vL9t9CxDGRrpdyDbowAKaAwtaV9nuAHqKYT
BN8NRxU8bmuMuwU8HLph12e9bYQyt2/WtBdFL2S0SCdbv0tVivyqs5Asa3Iw/tzZiN3QbJRaPGLh
omuQtY5ucJEV2+skf9n6RtJmt1jbQMNcdX+gVvy+28yCIRfFP+1xXTMUv830NjC2/2Ic/BUQERn3
HERP3cKK2ElvHLSnbMB6EuxT5qBWuANnhMdFBm81fhmWA9mub152LsZp/DAcrkCwGVjEPnSnooQ0
iT3W97s4ByGPZRD0gN3AZJgvGoEOwru/+w5lvppIM2vtI+H1brU4Oda2fU9jPK9MukYm8y3x4jxv
c11GvGnhBnwBTCxsnG36Z1706fvr30JERo+zfFVzGOIt00Mb0t9itKK4aoNiiQgRkLzb2E02VhV0
Z1/r6+8VoVoQeWY6a9Z8ftRWPm/t3oxUh9xD2BtjpH3oFtBjDBLvo1yD4tEaFVOnb0Qe1hnYyhLo
GRevLEsi3LpkwSU5QbBJMErZmsFcVQhUBRC6x+acuqe6zyQTVEp3bBNaGXdAl4vnsfj4uj/xIphO
GmaZDZvu3Od3zrpIYZXgayffSp5G1Rsx7uBfcczrFyLgYqbnsHGzfIC3zya+0e+rTuoxgqehoXwA
3SQI5SCdgw2mo6GxXKcr0cXpYxOO/1uI2vv9VwJgzE9ky9cUqDuftwvubvygYpwIe05QFluUaOS8
nNeYKU5PQSI/Sr8PacrpRwGONKD/gCsARDTRqaL4oV7j5gE+N/QGRyYfU7SuUVXmWKvchUEuSG9Z
UxyTM5UqrDOZzKO9a0juBeSeBB6MbKt74PTLM6yAmkml1o9E3b/aSfQDKPjyKqrA1YEQevLfiPE/
xhWkPGXHKi4ANK3IEAtm3sV0axsW0DzPx5FgnEZqkaCLrd73ehX+zqBHEkBsUnJsY2YGpETel574
92mWzSGwYTXcHx/VkOtHcRI1nzqwt/rTGkb/1ArFmaEGEJ0/mbIkdHx359k6Y6m8LpHXfPqwxSZn
uLt7GeYBCij8uKA7ooc9DlN94RyOVmqnatrLXsRp/RR0VcHLN19rDsoamlrG0Lv564z9eIRs+9VV
xiAWNE5HBbHHp1krjuR0HbWvBPD7JMcx6oRFl/R/eCHnXCHAKIr925/kVq9OBqHAW4Y3ey+xNlms
ZOhpc8OopSu5f7EWocJKVQRjUYGAr9MuTlQ5v+AF9HfRwU9xaBS5Fj+lrWeq0xJkqkAfHk0w5fy9
rJv8/g2PKIKG5MmpoB8v7z5VvwyAPzevqDY1XvYb2q/YRD2xnH4hGoa7E05T1qgvJ83GUmfYHb5T
2ebOdQ3o4rl1lilA2FbRtnU4sHHznr4rlYQ8klFm4fwG2yr40eEDMc2WNtlA/lSoAM1+OBmtKe+X
LFyeb/0DRuNQNsYI4Y0o4EEguLh5i5raqB98vw/4GdGtg9IyxUiCja2G2Q9HnW6Kl5c3utLSpCvh
Vo8gjRkYHMwdbGT6YZfOgLvaTQE9V8hfU3NfpteLZDrz0liM94VfVVGxEij98WEmFcPPKnycgChG
JQR9FGYVXpcxpVdmCNK25ul0jwWdiOVnIE/z6ceaPQQY1j8DNnPhzbmYCd45Cuft+Y0miz7fHkrL
R+zr9HeU8n1SnTI7F0u8qETOUDDVgzxAdYCvO/OTRyAA797ZYzS+LngqRur4M0n55+t26Yp52aJ3
j84cn9jiZtl4/mJQY/wHA0EXSYBzFju3zRXVhC34u9XVkqp9A04Wj9gXV1DJ+3ucmBOSliDdS/qA
YLWjLFccl8w3CwB2Tfvi/rEP/0IpsUZ2KJkj7PYoZPmT/VudmbHUXeaZd7bCWdXnO10rVLrUvbuV
yg4DSSsb5VV84CBuoYNItXKJwwfRN7T4x3BEV1S0D55zIGKeT5EWxzwfMNjErYG6cMdsKAPneJsZ
znfGbksAJkZvRDAnkfoDdP7kaT2SjAj4ReOehSBLed6SPy3OXeNoWV5hOH31BgOkpMcqUcZ5YpcU
AQTQjpk4grd3Kw5OTRuTM2nHIC1nJN+PyIqA9OC20WMTCn9/orxGMV4M7z+3NIcEGm7jDdMfrIcl
uupMMII9YO7qs/Y9ArUetO/YEan1SkZ0bIbs4lc5LRxIE+3F4rb7Gc/4y12MBgQkPMFQ9W0QiZZ3
EtL3c24WNWR5bX3PdAdDUNW/VzMKMme3pv15L6k8F8u75lwwx3DaVmBCDUis6SOscS27OTe7A46x
AymsRhksed/pa7YARIEMmNF8Vjl2y+IQKHsXUruRkoKZGRD3utvFC6/dB9rDk/XF9AyjMl/VNVtt
F8fgSktDyc5EvguMuQM61tp5AIRZjnKW9Y14bScWnPjO3O7JoPmS3nsVfOk9szkAf9m/AiSSLEYz
cWgTmI4LQz74Aw5LgLUxvcCeUpohMjZ8LWBUPGnrHdMZQ5vvn1qp0c79jJs715g1MHk8Ha5Jr/JB
UI5hQVHsPYgct/IFkCWCRU9ZHkv+15C5Nw+tnxIw0dVGXds7RC9+8ue0NGo5TXaweVMWdSmKWAmO
em3DnKSDvQsFKrrt0ecF2V3yp90YB4EldSbyQynKWDL02mBpdFkBI1e/Cms1DGZgWn7D2XuQDQ7E
zjJkPb9JCmB/SVkOKdedHFMw7SFRGwX1WrFrMv4WC09a4ICVPs6Ve8rEnduqdenoKDnMIu9/6JPE
pXqULxevm+qsNUKmwL5xhphuV/pYISYOeoGZyYtjetIofBAd7kfEkwyrPR4AIS1v/tLI8noSejQh
p3zrANXP1FIF85t3LWMp/c7Wcdox4x+Au5LX5uy1wiOcpiUAAlx18dTOSjlcJxT0x7mmiQH2mO5R
+0w8SEKqzs9bKU+lODHYPTO4lJUa3It+Kdn3Hvr9ys3kwn0Le7bSKXnt/OK3RixpjD6lVrPiqHz+
ND3PFNc0tjPHgTglRMe5VgxNUzBaT3EpkxEoD+iERD4NQkLG4RDb+/oBFrs+SCXzUz21mVk1bzx+
vrXZ4qheeFN9r+MC7L9bJGNox+3eNC2Y/h6VKZXz+v2WWnK51EumG9/sH6dXPDWN4V6hVitA8Mqn
jKLKF7Ji8ll1IwLPzYgeZx0Za8yRIP/dvlV8iBB/z0FvjcfSw39Tj3itLEgXdldxYZWBid9jtL+u
V4Gyn6epe74coyPuDv6GAGtm1g6JGsgvJ1zTiuXKCH6wg07LCXE4W4Hy6wkmUul11uMc9ggSPB15
G2Gwf7vvRimXXChPfQSu0zUlarstl0EpetEPbU7VYbuX8LQNtfBKGdH2ZoyL4HC7k8ezGthRCWy3
MoZhPuiduFXdVfc8uCf3WJV6txq8mfaCBY48/oN06oAcn3hhcZ62Ywd6k0yOqU88Ra5zoapNylJg
LFAY4oCnBodr2UvrCw+kXUKe+sSahRimkaUbbmxhH9KGjltcmv1hFR+4nc8XQSCQqx/7lO5w9iW5
AGu+Or6ihrBUV24qTXR+ntX2utjbjSYxHExxBgKGv3G9a5ycCPq/dTuKtTm439b91hpifjZpJsSY
mvAydDUFRYKEd1kRiXrZoz7jMuFu9Ro3gJ0smiGEfA3Xub4emHcD4ltjGIqPUA+HvcPTEriNzpBJ
4ZeDd43/aA2NNysTbVVcwT/b9Cb12buPuqEvjMbiN1jBYh4ZuYUZ2NCT/gUgYC/v/LHNjSPdI0fv
RRZ3z0SPW1GQafQE/4X2U5JgfZFz4KeNzJHZD/e1FqmM6pchWB+/8u2tNm7Wgz7RNkU6fPVLoXIQ
jn3EPcdBZXH6Yw/0uN1d0fOMQhsGC5yLfHS1HBFXrSPpcJkiT4bFArSeEdtV4RCdmi2zu4KNIuH4
nL+sMRjPzmaqkGZRekAHQLhMG8YJ92/7e4+c9NMB+edkC15+hfoAfYFJA+/xchIwitTkppCF6Unf
SMJPUvwWNXl1UFYemnKksopgf4T90QKIHU5DDrTjTAZsJ6/LfO1PXRU2CacL7glXTR4m65j/WAox
4t76T+aLZ1MUoBxcMpER0J4QzS/rM1oKvYQSkmGYxxVDxhq2CsF76nxrxJhcAjlueK17KTdzcBqM
cwRz7EonWP7j4RKgXQseJwoHm2lAoDAn5LC7bRMJT6yl2XbD4LUiD425jneoTOUoaAa56BvoBwqF
chd5xOJtfFng7wOpPJLCGmrk9cgA19d9rjMpZX/HMGpqr/gNlQh/Acw6GSFAy6+PbMYr0sDznHz1
5Yo9P+yHAZQjinIjEJA/901DJR4jvj3q5bjCeAiORrdoV30+2sfoJwUat7nsrKqZX7gJZgiSyVEr
OhPyFpfxh71FnyHjXUPmJXm7lNYpsYXsUvX6G/Oe40KpYP5yJffLTwMsDu9ND5OEEcl/OYXKj/XE
vxymQHDlz8EVvduB9bUlzE8AQedSmWb0uiGMO0ZDuYS3CQtcDRODhth5PI8n/P7i59AgScpkgBV+
6MYgciMjU4RQ19/wxhinCQpRV77S7LKJb92/yuUMQWDoDGmAbsV51M2JtV6SqJHOK5eRgKf0AlQ/
5aARF6m0AtRx5o6/5Vuh6O4aXgkUbEgBLUoywz1piB+JaNlZY5oyxvUDXzADyrNYgvjoc/W01Fkm
1fe1r/JGF8/e+ig6KrmFLsESIHLSqAe8IKLI5QvIHryKfU8DbFFzcMd9eWinvqbZiXLyBHLShWgU
d/SPrM90AU3QUki9CQBDb5fWF7j3Rj9zmk5HII1uhIwn4tJsfOxMAHoORZmSnQW0lQpvJgi6k6Zy
W8mfbtum6pQO6tNIN12NbtAtY571ZffFXrY5trNPEvf1+PRMLj59V1HYSIxPCEupgxU8S9uUH2YP
YSX9fSgGDKeFTrs6eP3MMO74v2XxaXUQA+/BGuM+D5Dju/n/70+chyaRtdRjDZ8Cm1pywSMtrQne
cl+5Ujn93fk8t43Iuj7P94sHhl/9V/0QAgEb3lLjYIGDlVHm2tY3SnfukvLdCb8IVChjw/TXzTJU
tkbp8usvKociWGtN66uhWCw0tsAQkEWsXmpSNjD/OZ8HhnCoSiyOFwSz1mOy7OUGAi3E+TGqmWOT
U85iQHLSG6YxRtRFVd+cFuSfBYVfva7NKoNCrC8KmULc7o6g6dM63Y/uguvNW2dqX+3/5fQey3fY
90CnMN6Bw/rP6pgC2KqN4rfsXp/1hayzws8OKMN5ZQKp+CjohQrlclDPaetuJmwFduGz7JuDvwaK
7gbjiYDVknN2ao5qoTYtVwBjzgGvU0yMcF8eDsptYNnAB4070yYsZ2MyjLk/i3HhG+4yNMT8MbdO
EoE7e9OqZoZOeZCFxzgkcS93/HDD3IrVjIsYg75ZAIguDh1ixk8hqGgJhujhmx+MWuiTP6aRp3c1
KtpNdjo+N2ze85CtGnKp2CnPb3gZSD3La/iaeYUKU6sv0PIqAfHDcyI303pNft4kGFNSoacEA0ZJ
2WxGxPS3DrefnXKg9HJ4Fb9WADhenD2T60Y2MS7cQ9Onb2pGMXIq8jJ3vBmhWKXzaLDxx8ORhdxA
kXmlMRbXBQO6qwEz1NhS7KCLZ2v7FOOZgw2RXWM6R8RWlcMDY45LQCtRxcmeYd21s3Bl/rI0a9pi
ZdfcPYJij7K3zbhOEUYDjr19AhQaLJ1MXcL4S9BR5NG+xyE13xrvpNTOXMJZaa7350KApUcBvBkj
q+JcIvJHxRX0qUeLi8L0uSKjb6/1wKPFJBA7lxQSiTfJot6nGPxoEbv1vfweiS26ok0uN+tcG60V
3R9Yp0g9YDjT2uhHNBghRV3p16uRoicCxt/ZWefkN/5v/IlfJrNO64ks6PGHYZJIo5CJwmfZAaXq
/fRja+7tqZDTXc2uy8gzy7WA8E3rhSFPK6FrvzFvkQJBk8NaRq98tJHKx8/zR9uTR/HpZsfbWZrP
rZZgI02rgL04RHIWN0tF36S0S9XM1E2gIiBxez/aeKgezNQhnqPbA33+WodVcxiqflOGEhipyqBr
akSuik2EgRYUrXFCOmnBu+1BPN0kEEXTARPcIY7zuo3RPqCS6E3rdPIf54nsdw6UIaZ2WTrCfWYk
YvgW0igy/TZO3/6ghNVuFB89ffMySjPT/KULmQrsOUIiGHPhrEmu1Jr8Vmp7xN/l8n3Pa92cD4Sk
keXFljxnmqbuTL6I370ukn1ck44/nbRlbucCnMKhg0Li/BLjPFPp3cnVEuoWcCQLNMgkWWf5mYj0
9OnFIRk7Wzm2D0TBbu1KKt+JxD1OnHBsi2EmIdmlycSD3jnBqSXjofnQOTYxVwaguK7pCfyn+g4L
rbEhUrE9X9WnGFdYnWhXoishTbeCgQ5+kaYQPbv62WDcUcueYNwSE/ioJJZXshT05ttYleCv+VM9
c1+rKOq0D8O9JNMjF+kVJTrF9dupplI/6ZkGvm+Q0uaMGQx9m2sp8S8V27bFQd4TbYasPdB/XgoI
ZfGz27mGkZhMcI4NmMlDRZe3RntjUI2Z5wq1F58ypPjRBHC8mZVJAceFQidm7Q/531Jgu/nDU9AQ
PPhr6dSvTVrGB4ynSogEwr/JaS3BgD+eC5B9vfTWiJtLrQOaDqmxSrcAvU2nXKHhwAYca8/ukbjI
7Q7YNM3UJkjKoA2tCz2U5Vp3m52/L5a7NL68yZp4k22CKi8f+wBkh2NZOwhRBJ8gu8S+x/jFFex6
mGX2uip8ZHSXLi2I4lv2IJbyT+s+f2F7swngRlNZcIpSVG9k98k0nKule5JGQzLt5V2Sw4POTDmQ
n4TzDJDPESw9t8OG4oKS91U2QRMcrZBowOHupNMdWUvofU/vr/balX+Vq3ePkmuIY31IHuerYv6k
GUfslben0ZFnSLL/2GY3TIozerx7P9nM8SvvxBXkU/5h+oGkvIt1Jeapfw9UkRJ0lia6Iz19JZ+H
jrPrzac217xOl4+M4wWUv9Yk5DuqV0j2L6LDhOb5KPYckVbInQcLPukLdHcZAuEOPs16NeRtRZ7P
FmRcT5+QxevQjNA6G448IJ9s6bqeL73RiHofqGWs6HAPBAuOsIVUY7Gt/pOylp756trk1k4BN/cB
qY3iA+BE+EyuNOzaYo0tO676gdm6/gCoxzInjgBkhrMZVdS0GPzTFpiv4FRn/nilrye7V45idrYl
ESXrkJM1GODFHq12ID8uEEK1fpfbsiMB++LfqmR80oc0xAKzxQJv5AQuCEyBM4GqTpemu22aTG5/
ZKoMiKlCIq5fYlaBSJ2cbBUaf1K5KZuGmfCEUWr54FjOZUyAN2AwTELU8KFiPxYMAMcdFnhPh9FS
gX6Oe50tumyGsFxY2LCtMgeNxg5LasKZnY6hssQFAyKyP6x8eHrRb+rIB7yDB7jmtRcFYYNBA89/
t3Zjd4m7EF19OjwFd4V6WcfAThn0ypALn2sXNwdPHXpLmpy9uj8uhXZoI+/bEvgNkEo5m0vDtOAD
/kEJiGSEqEBDKZw6h0cQ4nFq4vithq0bvQfp03y+vfxcH9n1GClp1aWBD/zTQy9JdriH++ZsZ7wn
1w6J3Zldd31DrRqZWIkD56Vt6X9Zz1H+t2bxD3GcFtiJd/8gRI0B8qzGE19r0Latn5udF2bNVfIo
2IOL9tuq65T3LAPoc+aLSJvxWqPornZpOXw+anaW7JbrBT7J2svuP4vJ5ufL+3wvCc+vyNPv2r4D
S+nHHp5Xw/iLVyiySISxIGuBhq30XYQkKyiEzqu2pOSy1xYh/xTd7xtLgCPmFIuRWB7BC7O1cYcz
wOYgTWJlJePVhYeKkpCXmkK1KUfnbxekEXcANZDKwX56Q9rT5Ec8vIBtuVYsLXI1es2CjThW3V29
5SzYw75TnS4uuk+6PFBLsUzlZU3ZvW7grCwlh23y+UJurn7Zmjlodj3ckUDGb7V0g08f7E3d85ZV
4qwRzUyJLBIKCf6KrdjxViFaJ/kr4DUiRWp9aesDzHOCxxCF8y9gx3i1IlohETqhqHqmU9EeeTcQ
a6/Sgqs37Y06tn3TT5lU9t4UPcm2sH+EP/zxd9wxr9CErWYdCcPxuCWSDcsjRCZYq/u6p/trZkSX
tyEAa7fQgT/j2UstTXuW0VW+KUiKut+jOCtsbFHJY9VxO4YYGm6Y+17jEvj9aOYgTjmWlZ7Z9LmW
v783gu4YWjQ6gG8fct7N8jKqH32RL7PsY/hsgPAdzDVWrdt9pZRhh/3jPqXFAtZRI7C/kLeXqTh9
w83On4vBrElGoC2ua29y86HJqV3HnVGXKwCvIDJ3ALFcAEWI3+ngXxjbhZSCHFPq4DZzKSiWaqBO
Z30fBhT1eZpX3g2zgXvez4lDnTBPaOsEQcdG6Shq4eLg/QwIWc33wuPzvZ4q3jPLjQuQblvgyuCz
LniBXTBJ/HDg9V5Rb29XFFPeO3Wj83ESMdtXBQFnnb+yse1mRyvTGsbTMgpJsg/DfEG2lH66vaft
Qj7g5Zp8PH+HVegz13YgKA3i6XFjT3ZfiEIRolWkbKlmCpTBbFGhuPbLMJdPYtplpYX/yohr1qZ6
AnA/lJiw0kYdMYhzfR9DD+jWVka8oPWLehvli2ero1GYeQ4MSQW/GCS7Xxxo5+qfFGNag0xBfejh
MPEay5simhWBJxiF0csMBREturKoTDfrLGD7L6tYRlg6h+qfpitCDhAR18vf0cVqSDp10Rrw1OeY
O4bj3YW7jg4b35EYviNF4ejxe0r9tGnTKFkkSoHIm+MRlovzKM887Pul/S9rbMdEGQxRbe61uypp
PQIftUfZ0P0osg2bNrfdQXupidjOeKs2MdFBVSBIT133WUqIqYmr9xFhEY8xklfOMFAU+VFAiB4Y
9zm/EV0eJNhl5ehfS3RzESSvHyKqcuWhBtkzdgkU/Gr37rjR/7nI8//nb+Emg/Dgh6d7I2PR/IDp
I75SuCYO1x1fGXza61eVnHZDbxwtn8OjeNDym1nhRMNbPT6090gcCcd6+uCWCCHKbqPDUvf7VPvE
dZRPZxqNZn00vj2l0vU+c+KlWNE59Fpp8BgLwA1cWmWeDuby33bJhfG1moWbO0W8oqVHzzqCpHJV
G8zC61KowsTLrzYU/ZtVIvtb3uOhWiMso6h+6JVmw/EWV9jqUU5i5La1xVmtX2PW8yBtMW1YzLnM
3FHkX9kdVsd+RBHk8UXq11wrN0DRvmi7IgGelADWfZ3RbWMXb7mBCEAeP0cgLq8KKiIzSUapEkiG
wNQUIveVnWkpk24mFhvdZT+tfHgc6wvhwC4CN03UurQcF/JILM+DFLejujtYpzLCE6EbrLd6L5Z+
3zybekloFO9X5I3S7nIJ10AKwQyPdUZBS+/Tfw14U18K9A+atyIpycr0kvKx+c7rqkLcSB9v/T+S
VDTrzWlgzKEtXN6S/AK9n/O9BKdMrbaHF1LgCIgy2qGHfS/nbtg1jOaEL2dK1rLMKUhILFmh0Xxy
Kfi/5OwfjLCktZ5KBew53ui9Tt7Sinf301XaWiDxaXNAC8RMTX6SiEYgNesbWck5CtofNNNRCD4V
L6FlK0WcXobdMFGCiueA+lShMr7rLHrkXtwxkjeml6+QRJxS7nVgLMRgRByGTkxcsaSLb4Tmz7ip
K2EDx8ho/z83Swxbt8KqUNwBJrJGpSXII0kQBzr0o5vKro9PDoajBPir3Xszcg83uUwqXiF8L3UK
nTbnd9ONEI6ItuN5RwGbhX4ErziiNDXuX7PfClAktMSWN+xoICqTus1M1Nr+CyyXL02Am5XzqIYX
lRGolLOpXpBMZhRGMEbGSQvQL9nKUkufSiVuWc/gK1Gmb71ot0AWrEhVqOSYXkV7m3wXw3TDQRB1
hDhmtvHwzMg+ETwuNOyzgiYQkN2/YgozDNnELELLiFggy3Nl00bh0PZWFgJ0oPhhzddaGQDrf6J8
/rFITIAZNSE2uYCIozaNDlpRhBWfV2guA9um8zpskqeg/hU3/czuNnciTAaKf0zgbGMS75KL2rXQ
d9tIgPz3w6laebp1NyyBtz1UH2jR9kMPUQi7bywG0J4TMOo3M2qMQclWocJtHMAFQ2I4+AXVaIsI
at1kjPfupVM7ifkGRkiofTp9pE/zI9nXCqSHjc0NJ2wtr5rQx7RX3cAuCs4YM+RA5KaEWfOjyaQW
/10EVKe0c4WueqcLfCIhD/gPsgjBQjyskrRBO8+HvsB0qmkd7qNtSTIFPiNHCevjnnVJV1PDamaJ
Du8WCnwkh69DzQI7rdbgGCls/Ji0A7K6AEmXp4KCan72eFsbfoLbNP4jYIpLT0+jl3VevIqP5eHE
mb9p/p2RUC2IRWJvwz3i53Eo6h1AI2OCZefyQEY3/1/+NyZt8A/JUvmcotabqc54+QT3V6CyxgKz
nf6GD5od7eAACGWUqQQaL4SNLT+Q9b7ZL630L3eq1i/ivqGOM+y1GIAzJWszg8rPm4fAfMxXwETr
Wzphnp9WPP9CEaCBzRqjvAgIn9nPwTLFLGfFpv2aBWJwz/ymg6EVzOnj++y4rZWpM+o94KEBSpwR
QOVyortfAzlGQrUtOoXJQ2+gX5C0mYiboXT+yo0tuX3FGQoATLSsQmBVIDBZBF6oK6S+0QaT3LY4
DYRG+zsjEJR9TNP/cDxob0N5Mebj8Y8WHRNPbLJyYskn1Jfx5ebHuNEzt8N0cYaxBRQtNIiFP3a5
lCRD0pBTBB+8vDjF7Z6aONMI2RG+X1hCS/t4O8gLr8ZqQBWaSKkxD95gLldmSRT6I2qJYjSDaW/D
joC40BCe2rfsQ7CrM+UYIEyn2alFV/TEjHHuWX1N4QiEldWlD+xu1MEiL0xKcpuQdBCFTL1NavK+
n8sIqzXeB1pzi+APOm/gRW+F9Ia2rR+KGH4sGMjySSrU0nDtcOpnY6rE0BHQ9/nR2+yCtXj3dBZC
uDqagjGl128F7usclR3qcu9DFgTtNRGFiCik0wXVYf2KmdJvTiJJ/aJjMWgPUOJe8+fGCLQ81v71
T44r8ETQkLRnj2BExBcslEm8CzrUZnRooF0QVuRWoCAZlpv0ck5aXYW9A4q9wV0maj7iLvxquKf1
TNef4uVyiEAXX93CrDz8SEPUC+j3tXe10eAQPd6gBPsChddcMT1nklopyVVderrkDLXnIQdBlBsU
ZGfS6T/ChENWHE/nzJmxOK5bkiqSROdJn3d8LeB7FPK74I150bQ74WMxXwZEBuaEc18Rs4DyyXXt
P3tllqRciQL/X3qxDJF+/g75YX1EEMbgAJ57zVG3CmHH7WcrZrxSEZTiR2kg41Si+HwoO+VYmX0D
UEXsjzlGO42ZCh+4L535NqMPo3fdrk5lNYdB0UYcV1CzFXXfoj0AWA/RjJ6pWm4NtHtGm7vRt5KG
QO/YOP3uwxMb+O+NcWXEdG0G1vDB6aiekBXZVPagyfm7Y6vjqVNg/IRVSGnM4E/XeedmD2RedJcc
EEViOUwDqr61ETWkyuOx65fuA1eq4iunRx/Ii6680CQFtbvT1JplUqG45s7GE2doKurX3hn/5vr3
v6Jbua6XcnrPB7bYrmMQ3V5Bsr+MKCBRPzRS/XR/WiGieN8sAmoa4YCFRGqCKIfLg8Q5AW5UdvLu
R2wJ43w1gvlfGNuug1E6GxEctVcVe2QIxP+Ezre3OOgVyvqcWJNhYBc68QOJcsnRO1xHbHj9la8d
xhZXKLk+FwcTUqBOYD6pEdFcgd1gjeC1yqDMdltvtV2mw+/dn/BIT+RcAVmmT/7rQCw1D4N4PP12
r04Ya0ymJAQM0I64caw2NwqBgzI0Ou/9VF2xYfyUPzZpSPGf4O2ytPDoY12YC+UGIXuh25M7GiN5
IuDeTy5pS1Ss3FenoINwOMfcnE2JN+m4oW8AnMLTU80zxem6hlglhAdjjrGOOfmZQKd++t0/HzBt
4Z9rbW9ld0b7gZmBjeucfc/aQLgSB6CmoysX8AMsQeOQj2E62XUyXd5fi9eNTl6pqpVpJ6fdRbfk
YeQghQyl7rOywW1v8OoHX3tiD/BMvhDrtxNMbDcPt1a9JFVoSI7X0UAStMhBqHuopCWYUNtB7beO
ICEyORwpZFESWs7d/5ncXCE0hig52Ebl9ECW95OEA4FCvDq9Q72z07/KfjlACwimLWIXIftCNzAk
O/KpREhpRIss84AERpyK0VVXoqhEZuFc2NO3gbAl8bllEoMXDk60jilRDvYmSF/k4D40wuVoiPts
w9IxgSdk3vFu8ECF+1teIUjOX951LKGDTf72Ybn7BwE+d50HK4KckMIkcSNdV/rEuffB4WCSlt9m
mRusn/ESj0d3fm13vczrD8WxMiQkZ/wtooqiQePGU4oMBXZyPzh6QBd6Vadrhhj8wnkB0xphPwzX
1Mh0lQb4PzWinlTtfwXNagDxn6DNhS3U9frJI09e5Ek7DkQeRBbT2gVU+KXe+wRsRmP6Kq7TGzEf
nc724KFNkaFYvfDnS9P2IeeTxV5SGaQGpuYOaiqP9rwOKY7Jto78Pm/IDe0BVmUTHCB17DsGkgVj
x8fgD1qL4qQQiVYuAhWlPmk2Z8ZdXZd7Z5UhtkvXDg4yA9zaSGpTGSFFMGPcXKUS5KjKiMSDr/8e
E1KnDbGf0FejtXE9rHVpQnBzYMD2a611A6wlOSHwjcT4/7hzc+ay7IrJRZ/pqEthidwLYprFN7tD
KrBhx8zu202NnOdeuzJTntbOhp5GF/+exwfRpI0KWT1BM5GVuGxjf6CujqAyyZ46c3UC5pmt84Ib
vNNrzWyiAUTV9793WYCs+ijvidV5ZNi8MEVqnE1MwxQbumh7r3ZXF+hQgarvHYxjojvPqrpEp4T8
K83fHiHjGQCfB1PMQOBt4K39pm67IbqosCEXjKFzV92wRfYvuvJXooZfo6R26TK87K3KtSZCUx7p
7HSnXlZNTP7INrpXS1xpTly1sauNoUY9/I5CqH5RTzOx1lrGueeka/ZKBHQUELJqFcBp69hGyQ+7
It2CXUsSTsIuV0d3KUmcGV32RUfvgxxTRghUmUYuR8OIb1PlIw/0BALxhAkE+JLanaBWl5WsM2ct
SjJAMC9J0c+TMKVH2vThGVjiu9ZNFPRzHB/djctc6IcSyUfjoAOuqdS8coenwAzWLXvM2bqANjP4
zpJ2SW2m3TzNhYjVxibW7W4T9P0qq3dtmh5I/tB0wFLMsuTgmgh31dBLy3m4RQ2MgLiO5vTkvSnZ
glEj3HwO8r5hpAyH8Uc9HMkqIUVyircJe0vnd0ZArz7eEvsx1UohZzMSwzYc19DqUvQ7A/WgJ/oV
+4WcP2WQGx11jEENhfxxRCDKIy7LsdV7avd7iQmeZhX+RM2tAZ0KXLgQcef08BiTWeHxkRbLV0rI
KmCaRLFrlKuZo/IhSjvZmaFYwsBwJXRz2DOGgFYPwRv3/FqMEKqkm0f4CFM5y6UtSj88q/evwc5v
JXgQ4VLnv6ch8I1mwuvt8LU3nXBrj5hBlYoqbgTpRPlRl9/Q4SJ9Wy9HQPhyT+hX5xqU9GYoF45e
U7mwz7OkEo/iCAzqRweZAvnlTJIVxBbdYNICcKCEziWRqOBaDbW4zEqulQ1wb53tTBbfApitgWoX
PDWt7SOBPWuPnwKz28cKKPXJlwk8wtzSHCylAbOjVE2/SShBNo3atTmkYVAw57gTZEuSQxyc+Lon
lUYq8kfVOu1JNqSXTK0UrgQwJRr/FZM7cYYUFH5YdGmZ1/qK04NhqjCAI6smxUbb1h3KF7sZKECf
C0X2gfRRYGpG7yiOpTDcF+nelWl21Prw5ml/LMFPWmIi/VHW6SH7iYjffOFjz64XITKh1HpbACRC
6cRLZU0FD5tAPGjQtv+PHSi4skWcfAlsiHUAZs3qWjVt/Zq8o2QI2w4R0K9CpelaY+ViZkunAmtV
NLp40l9lybsbQdhLBVyiojCkbpQ1r7wUxEluXak131cbwnbjeyf4OhUYkCp6hulyTLyVzThPiIUe
F6gVkK7//KdngAVi+RgzhmTKnSe/DYb/IPjQ+2+/vdbYiVTF0vIUBzNsQ1Y8PK08fJafNhcVxu9K
i94PiAF9ZDgU7S3uAzS1gqdjdAqsxy6x43ihHtqLbxA/Rpeaz/h5FxXL8JMY6+CHICVTiu2ChTLK
1ZiRVcLmCcdKo55OrxoadSY857/yDs8xcnEAQDqbipobvj/VCRiEZSsoZtYS0h76uXLCAl3QFbCA
UnD0n2ULfIYvLpySrFAZy4YDG7WL8FvCOFAEMi2iTbsDMY2xMcl7Qy+YfXuL0jLOsVFs29UunCkO
U6cYgp3VtdGfgvwChqj0TSvOEJ+czZ0HnDO5n6ivXIKMgX8uNBNtIq/ULv0SoTKcquK3GhzXufSK
5AHJ/cHclqROASnednQHgIilzXgV2zC4fDAXE/dXvkHIah/Tr3X8SUVgfhIDClWtt6+KlrzJoSAW
rP1IxaAhWm4a+iPK50cgqpdA3huZ3P7c+lt4tGIhOwRIqm9X+HvQ5fCz1Ca2muanKpBdAAbsYkuV
HyrzA+e2MmX7KcHDvlGT12W8FpbDEwAbA+eYjF4eLs0VcGNwycuj6ss37Q+TGTL3rkPFPw6gDpMH
0eadvCvph0zVsznt2lkxOLPZL/F7c09Ow0/+DmlSZmrHeI1ojpcpvbDMPDFs/QzE3kcBirStnrtM
Y7INHDvaBlWGlMjWG7ivoyEf0ZSlVlEH7k6t2tQ68+kYcWa071HjSFM8lWVrdIUJTH9Ft/DZiIB1
FW18F7XXzsXeAa+GXjHgce0qJcLgg24L/WSVNYm3Kciu0PJa96wH4uJwqCRogHWA/ioHLrxsHozM
iYQ3gwQpg0F799gPHJUG31ik95VmaPEn5pu4y/KZvAMPQG29OplzxxYrsphp+gFl7D6Fi3BizXM/
bBgoPilqa+Ry8vjbLKdzgMP8DM/ZAdLvc8JwOT/mg9nzcrdq5mUNIzP0eGBGIyqR9fmbdWf5f681
AHzhPMcQxiGnUXxBo1nw2WwwPE/NwjI+K2C1THFyQLNXM5bQ2ffC93kIDBjP+pu/jhOFI20Y/ZiU
PCyVOte5iRJifJpGN7+fNWhqDiVm57+4+jpGao5lOiWx4XU5DPgKF+QUShs31mjDvUo/I81FRLZM
sx4+NLOBOc+OZo6/SxF9cHt6NtZRD5LFMDqcPmJdhE9GeXohlitvpWcKBOmgs5ZGS7QJW4SRQlOf
q1dhYJPtnxvXbtSvl/lGhcCNaoEvoiqvLoX4+qd4RoQJZqWu/tBd4gE8dIULRjHH9b3J01O1DPhs
Bs7kpum9dP/+ATqJZVxC6ioPlexWJ+/NdAWrW3AK5uc7eDIz15YVwysN3gKKsTmxHKvAUYHgWuS3
y3QH8PI0SOAz9Pjsap8D/3VyPqDlM9Tq6kViLIzIsU1Q48GdsEB3x80A/HcUWZxMUy7sJxUvGPBp
B7GtlpLBtOkHa5487e1Kd/f03EFl9tAYCXy2SSiW+HjLr1Er3n6IR31lG/GkI1WphiAhYXYeo+bV
PP8cQmNz4XDDEaVoxYaBAhrrV37/yEhb/h845h0/pOR2BbVEdBFVFgcynbR+vSEA9Z0PC6Jdf2nu
0KdILQBCpRLltaBHwoPMQj2Ih51tN/+s73mZxnO6sB16x6hVC2ZJzoKGqrEFtGg5lN0G/7Svef7E
GvrGNrKan3m5VitesvmEWcT2yRtPQzZBNyZlDd/XcVYiOrJBvk9/hSetT7Cof2XOp8GQ/Tw/Ua9M
E9CVUKbdxsjQfT0OhmcsIMB5xNN10ivhdLx9fgHcXvNiDMh/kjNuU+nBQEHaH96Cdf/SKOfQLPJq
Ky7sVvsBbAt5jSkthGrvmp5FhbZAp1gSJ4dzUXZgi/tZU5Ijxsxi80XIvIA6gLf16h8w5a+55Cqs
yJ8a4vwyALGC32hCSa75shDIV4Eq04/CGsdz/vBq+asRPaDbL+eSVb/LZZRzMPaTdrRCLKmaJ/lh
skEDP8jeFIsCcJhNUy71ayvBlqIOu6Mi5lm/9IPBdX1YCbOIy5tmDIV2ohvtzrJ36eAe/NHEwCcX
oNvnMgOUZNBgAFJIMs8xLNH0hawjRI4TRAmIWGkbkUPIwX7Y5cNdIQ6H6hWX81zf4aHaTY3NwNDI
5dT+7Dz760LYZ5s2uMtD5hAvTBe3vJ/Lb7IPcALEuwIp5OZ2gZKTuW3g8yKh0yJEivg+rkmLwrTE
e2ja49s7giLgYSV5WG5ILIb51d5YLHYyJ9HWD5S99g73l2xet/5xpb/4+Uf45R6hkH2g3a6DC1j8
wzwXV4YfM7Pj5FMiaQF+xZN7RWuqjjrpX0TCYhTBvH7oiYQDZfo3awIrDfXpCWl6rKhRJJhy/GjE
oB135RWqgMn2GwQhgCJe9C5fc8SOorq1Bclyt+htK7MiqRRyjIlzUHKHx/7+y+n4HwYVKPy0q3Wl
XtLorW7zf0//tasyC+Kc3+jvMEKiFBzxbiCbFFJjDGRQVyhlyhXDJzGU5hRi1KXdscwqQFBdQ6Rl
UG//EJNaD56EdeIDMUTgqsiWsWYwWwSHIJvQgljZh/g8CbHiBTF8CETXNlbjgTWBvxhRcp/oZ63n
ZYCpbZRee23wgqmtZJOFprEf2vBG6J7qjwcyFlDYZ4tmfQVMWVgf0KyojslJGSBZUMEDekKRVOSc
MbabIeSOhjFLno+mmeHJvss9uLvszCE1GCyjhkzEkokAr+OemMKn5Tyrd4S9AjGP/2bpd+zOuudq
PUulACUyv7jCaMVTv6hpC8V648c7yMO8ppow/9pPKLhn24ytzCm8eFBxIj62VD94FrxgHeGjFVwS
F089GrvoZh0ch6vLJVy+hZOYdqbThokOulscRzpb5MN909Tpec1XQ89foGPQuKn/IMOy5REby9MV
PR098j/GoVPmL3JlrN+lvgCHyhegz1OFw6VDcCA554wGWm9Uog+JEL79kdG8HPtnH2xYZTKJi6ws
pCw38ARhCNmbj2KgrcvT+U4ajNdgd8W7/JcTUMmCeU4KYOg1y/SFeGDOHTQNQwA9mntGRVnJt2cX
EQjceEyEVGNdYKY7BE2qyyEHT1MZCybxd+Uc0INuGqQ64IyJQr+UD9CJtXkrGQq/vO2vd3v0ik4g
yv6ypKQvlokrtBHaJwJYdZ27nusCfaIZqArHwuZrMpmvvuLUHUjtlP4E5BwdxmJXhpduo4Vp+hL6
8veQgrqDjD7bnHtkAw8ILBWySfdleNDHplKLcwzyzZ84Ih8d17YwlVvZQDApFKOjUbYn9kBXlgBP
MskHrL/xyIfb0Ra9OND/tKoVPDR6wUN8KqJTOE4u27g0UkpEZPK3NlUXm99u/JMgcmc5uCgZ7Yep
v+s2+eaXwcr35M5o94mCtH+w4CWSI/L+reh71jzTXCPRf3c7e8bypNQTAy9Iupo6TjnCF4relzud
9aU69Y7O+wYEzZZQM11NT4SWtf7YfL+Ct/W5YRxk6o+rCok5P2Ik4LZ2n9A72amAkgUwxt6y5SzR
Eh1/B+EWrRWoMfHhEOd+XqH5efcJ2YvuczXfwR0s67ojp/RzyAjdlkwiVRkVrFQT7Vc149jmoXSA
Zpur0Nj4G1s0dp3X39Ub5OkyT91Aa5eoYQEsLlTElcgrlpu58lD/16G1SgzWdjzdRKs+7jv5QgSY
74ex9vlZmI5HRaZzVi5BHtX5/OrJQYtDK4kpBVhcYvHouMKhiGKVD6pchDY1lM/PP+ptfuBd/n73
Oh4BjXO0uRQhmvpcpp2zs+fiDBana8CnaDy1MhREevAyGfovJVoxOAjJjZQ2xSU8/ljgQGQauOpJ
aAkbt/OURXytPZi/Grs80ImavWD3MeOxhrrnh566qZfqjsCBCv2n8NV7DXzM0aKB5Yo/nuyR3oSD
RCKhyFL2qgpTAsPHRne0itmy2qCOYfngoZQYOg5g+dwKATVbx3gBbapWHukFHP+isUDF1bVbavRm
UkEeKF7jkizxb8tPIMd0r4ude9KJhurp0dMiMb/LMWlA16cUYKPpqFY2IiBJtqY7CrkScuBVk1AY
qLxL2fVH+yA7Imi3VWS1d5gq4MUI3A92O3F9LsYBmeENRtMt4wuxK+GZiQjmWeSNUUnkak7nfR4U
UGR85CSzllCe7UhXGvjJQ8jvF4vpyexem6QsluRqGy2dsYYlkipaNi6jTK1i15ZyPdlJ7vow+es6
jTMhyCwAk7CwSeQNc2RcygLZCIbm/VLavzC6HPjqfGM3JjWq8NshFAirb1RMUg1/O0TQ9BJgCSUC
4u7xxRe32xm/Lbar/XxRpWx7AnkwT7pRV+JXoXKnXIElOvuv4HSpBnQZSOL4Fe0SMqfXXUfZgRzq
Z/Iy95lOdYkEYHShObM8Uh1HVWbxyk0ssKh5PdqRdx2pupMQ4kut38uBKEujDScNfVpZT8udSXhG
VaEIWvxbXj+FE2QShqhVuA8eN/WJ1yhZ/nqCgKYMXWe3+0+nDJIWuqQ5ZJk0tG8MFNXCgTANtgIH
DBkhtXgqllNEXOvDHXoBnO2nKf28F0eRqEU099bYkQvg7ZHfBmbpBwpi9fwQ6b8cKZBS74XJavqs
QEga86s3C2q9nAfTUtfhBsxMX/B4qUgQS5f0GfUqYzafsq5VNrEZywV2y7a7oYfX+lNtC4WNJ9TL
T6ZbuQ6rprOek+RZIm/CTpsTeTM/nP47g/Vf/rYovFjJUH1dQoSfeXUBQuuKXadOOMWwDMAfFl0S
BK0cfDUwlqV77mYyKlQytCbyN6UFhe/DTWud6VBpN1O21ELC+/aVaJQIKZiV6DBbHYkaJbbP+Lrj
m2KUXQ2Dou2XmoY/WARHgWj77ASf/5JaIGMnngUiQdAiZ6NBKFqr8G4CxaltmWTxPNzeMryQjmCZ
W81hX42vCCoXdM+opXLIuo+zpfkPBD6hvfcLzDMMB7hcOIbCv0tNRm/DeGPnasZ7TM3yiy7W335S
5CG7tEd92TRrHu3hpve8lJcU127gfiANhgSDNihswUnYtSqyTHJybULsh/SgSPyBCNY4dKgqaouT
mB/AQ2NsdnlbuWyM3I6kSxYCQOQqjERHCWa8cjbzVhdIozUw0fHT6Qtc2fQJ3OnpcS8UYz/fmt8p
rNAmmHODDvbsfSEffmS4DomGJ36qhiJ+SSVFnHpXQtA7g1oB99q3XP9HekCgogMnuQkJmGw1gsth
3LxntxhjOmKKkDYRrP9N2draI5r5WONMoAsaxig2aM6STPJ169nH2NM5KGvTu9H4SQBrrpi85iRb
BBJwWm99SHSsL+aYi752+KAenJfZfswMa7gv/PBWY6Zof7SMHGk8pgQ2TURcVdhLk6DGgqd6cNoj
raA8cAmAM74RLXcbH2PAd9Lx6I+kScpmcUWUKh7A9awAkSXLnkSo+aOrx0zpfVaWimGQcruh4beY
nWhKbPo3aBHdlB64sljfWATv2k6iYakt757TUCiacolLmhjeOjj4muo/r9jrnuzwYWGh/XqUr7ab
f7fQ/sgzbLUDLFk2PmtQq2FbZZ/Nyjjl//0FJdmqiNwKWs6Q/Ao/NANL91LFic0Jo2e8QX+oHpl5
oZWqBnowAbNKZyiuD8wjZrHnHfg+6LL1hE2WasQanhkcdxUDoJzIEEf4hNP4zuyfkCUo7m5HCf8A
N43pIAWq68p+y32G3FqdYrrmXXh5VnjyExx140DpFrAlS51B9HxRCUpvhErFNa0l8fm0SiHU1qqq
FLWzaCeV2w+ZOTij2Gbs7Izgb/2qMDP+6c80MvMw2qdPVXmBfU9pmCHp9dNRf4EGsnsenNawQe7L
eWkKO/QZBzdgZakGy5rqe920lgN97jxsj5AUfDR5WjZtMX4Hzaviy+FZ1Evv03BpZMv95q1t6XlV
sWuJqCR4qGyu6l2gX6xvQBGyhMcOog5jk9iC5rR4ATkDpmICTfrWk0q5GorKHJGb65K1nQNsvi6V
mp0H+mOEoS5vnTbIXLjcxYXqgXrYblVKDl65Uo9ITXZCA8gyQHRoyX9RtMuIeCsTmAAFLXkQSmv2
7yKNV907EIhmHvNbh5NjL6CUabEN1GItUbg4jNDmcf5YQ90uGM0htd1OZOWnKX1ramNDta4BYHl3
X6ULRl2BWv4K/D/FZzB7yVxtP5fVCGqgeMpY7/aA7hgGJTgwvxc+cigmSW321SKQqEaI23DRvcYb
pl7U2Ju0LAga26MHQuvCMTVzpoKgiBZPuFqx26Ch8iq2FoKYIzW0czpafQsPyLhJDZJBMbgkeVOb
b0rXQF6t4E7PjFfb6aR6Uum0byWDg/WXqiZBxdMbkWHxMXl/gSrgiUfI/ObJgpX317JxTpGHQNa1
HvGn/oHJWzIyxWPb/XR9cCCKU9lSR53WHz7i2tdfCu3u7Nyd2Yru5OZffBxvCQMN7ODxjT4Hi1Kq
JzbfFqWOFr07zkn6rO2PYr94OlGWhh2/MTx6pDCd5XFAYVRnSUd/U2vlPs2cwLeu2cnx8tE+SfBQ
9I2N6a433b6Lg5tQUYhP6h5ELUxfgcs7zrWs7jpF8fVbQZIiFwVpLsJtTR3LsOMb5UgHHqwfE6sv
fZTPA7QArByZFEHVxFNceyM1Z947rN67kqpv8GIm4pNvKUf3yuuh3og6yKi4S1/j+xA0OcPJdgdH
nPNBlgQVXGEMXw09EqmYVlbn67CA7Pl7DqCOmIJasiXPGmfxl24otNyxy1cmTKOPWw+Aj+Lxv2g0
U4NWG+ZIDCuHY/KMnYp0BsnJSfuVzTSsTB/UKOs6noVgOLW+6N3JfrgV8nlppRVFqWniispLYdEx
riDKzg69O0SM8uTTHC/FqfOxPP2Efiqbl4iT+jDrXzkW2p/I50PxhNUUuOZdxFzo66hpXvDFZAHf
kgANhnqw2bjqIlazQ9dtPO6JjCiFtYZZHTBPfG7FP7MJK3jKNNVCSqtjsQG8HsuDQkmnLdc2TMtS
L+pzg9kXKLjJcjHuinIRN8GlQBLlMqnrPNRKQeezklLCmCY6gbJuA+YcoYNgYvbX55cwFYGgsE+S
Wzy5GjWeuNfxX8DBaMwGaK6Ke4ITCsgUmAZmg5nZzt8Tid+FVBpetf8mzwarQ4ACuAN3BhcOIUOD
wAbRsq9jCzc8+KhXoFj0GbX25CMvYMO33lq5NVp4jOQA9fzPTL7bJsUpUwPLkuW3z1YVyAu0MrXb
eKWbEGV8bAhWd4tNI4AwUkrolyfBOqxLUXIZrc7f1ML8sErkCEH6f/jwcBZTX65rmxKEealgnnl3
KN3CuO6g3aF6LLbOLjogp9FazAOhwEnii9bum25BouLG4OXZhLTB2p2AWTTN90D4BildnR9XM7dL
n6BsbOLPlnFi1lxFzuIKUM5deSJYVjimMz3FK/Ys9cv+g2xpo/d3ouTu8E9zn/4SOt/dM1coYOBP
/dunTTHGZhrxP0HfOgCctRRt9zot4gpocLnpo4rYh5use5QGtXfY1ikDYYj95zKY22uJDPbaz3AY
zVfFWaAkL9H5jMI4tyNfphGUUAY9Y34reAguI5GUEt8ASWEz/yr707X6k5w8gwZ+ujvu8BLbzy59
vigBDos9eK0zKaSBW4KfKMTSe+yRsxMugvL6gG07dhE0Q+UTEDrZt2FfidKJmFG6yVGOp9Y9/CjJ
0iNkek0HNDF7nP8YGz4UNWikbuYF7RSo6cpYxgGjMThCnbxcLRXBxEj0K0Vm1rBw1mgCe2PdVSVD
BOPQv5aPqAKBx/irIpJw/IMK2OhopyefWYL38b4MYUZlmBp6Nh6uEXRUgGdlnJnaY6r4E7Z8MhRw
tV2WVETx3iOijoWquZHjIT10z0kKx1A7nrP0JJXY8rZgg/RNrWKArBppv2EUFdTslj+vWzlQq0xd
fGIUXQ9uYdXpYuZNFvho1pWe9TNovy+kKxVN/RLzxc95Rg5JOPm1VUOSPS/roo8HjaT+3HE9adqy
3SRP7QtkEjvxlFSmVNtCr9oNYPpyoc6j/6M7n863+cvk7nG2sdWBWyAljwsPrOPJGLYCVlNNSCs2
0nUqGd3K4cL1wNHhQh4TjXvf2q/HWyL3as6kMfmvny8XXHmhsMJLTNoefUgVOJGBlAbCYLrhHiwf
9j9Xd/BqOmTYfsAafamjvhooPAzaBNuZC6VMVCGVuogowAf4Hcnbh6J+J7zA0C0nbrIpsqenPLrn
z/PJjsKbHwdw2biz7KKjlHakWaIzulNS2kgr7Mn8cKjSSA44TlFyNkI3T6HkJRrOwP9A/ZE1h05F
EX2DUKONwfQMnEkVbrlgANbIrx8PVnncB3iiOgSSWSK0jZN6wnItLF55MNV1gIVzr79uybtzCHAg
w6WXXd0bv1VMERCm/JNCXm5CaQQrZt2rmD9MRRzlCokddywEEXxZCaXh1sluGhFOtaGgRSJkeXYQ
0/4StHUyX5JwquaSyMA83zSISJGhinVtg2epPNez3XSgjhCLhxeBCmzD7UXFk+nrX0UPQEPG7/hx
fgr3sbXhhkyDXcDTnb1rHYXVCW1DN9fUqAu68y3AlCqx+830Id32yP4znKK77umrKv9xRoRH7W3+
Zp4lX45t3/PfGbOnY4zuit+WKkYCwxYg1FmRVVvZpzGfQLPreLRbZS7TIkVJFiBa32CeWaIP5tXn
xx+8cOROI/TzGAOJLW03kZPUY4PlT3vXODGCyDNMUYqXetCV+RECxQlPQ6+WYwOMi/+erzpj5HoL
EktXTiJPH8jDyySd9P0JChdyHGPStlKPRQzZbk7gDMek4lrVLcehEEgbhYWXdIEjfIGs/+suwQ5m
Bm/657wsU8zFVW/QLSQ7kSOhsxgG0DDIQlOG6993zoZe7LsZX06bETknXnfYwXxCA7bXggDqBeNu
qDjpFvzfN2K1HsjFLgmhmICdn4SLpad6v7wTcX/nFtTYkG69W9mXqs4sWaCLTQsnA7MzBuZoxa0w
Rrrq0fG6hFucnEMFbjM6rbWdWvvyOafLvbi5bKr+4Zg+iSgz7v4pVajnpYf8gDXfWquBQPvnZ25X
GqxnIGq1h4wsWS+zN8rjCVTDz6A7TRzh24dwTK3LJTxnFcio4YrEan7S6vokybMCUyXH3t3txm9w
OeMKrlgZj64q0GGrV2XlxhuPZJvFM7R0Z6Zbm1a3OdGk1VRxrOotarEEjsk5dEWGQrPGMkhBZqQ/
wHnovs4G49ufgd/6jNC5zkv86wGRw1NdC6Y+NVcG6ZuiMXMLLSVALXD9YEAGAXHcQtldqul8jzxK
sBHMyrhuFFRKS4aF+sQ8/pk9CoCF6qGFFSIoH3fvnDwJluV9FfvoIagdlhiFqrlvPjPVvYF4wTyP
DPN3O8Ob6WZCB/xeLrUEJ+r6L3TZsDwY5KDLAwHmUlKN7fzBEZeTyxIGlCEqcmvHR8682j31Phgq
ciIJaTYASWLW8cpD5D3pMzBe6s1FD/Ljp3y9mUgQ+KCNFYZ6OHVkyxcV5ymQBcxOMvEcwy8HH4wQ
V2RRmr4zVZ51onI/F/WM2uqG5sAlaMoFYdSLk/i/LsUpgUNzbk0GIESD/m8QYS9cCXV25y8Bkb6O
HpQvccZYJFGrSM/+7V57ebnOvcxXuZP3E/4WlDNO8/y+qNN+GRg4z51mgvqFdFdgzgX59Toy7PSm
BBb0Fh24LNru/LhVfxSeHw4c7krhArQf88gj/Fk2xbZYz9BFcxvhH4hXty6oaQiNXTzLE80vvwfp
aP0hTFkK/lnPnFjp3KHr8vW2DeP0h6N2uQX3Aasd0CSAoffFA7JwBW+r2Vd+XdPDDoDGjEkbdHBy
nmgl+RTWCYE5touaGcz18EjNBqjWXDjn/vItawF6GHeWfPZBr0gBFAT271AVrpH7fNKzkIkzd0rv
eQVxc7UjI5wQmXkGggZ8LlH05zZf6HcD35Zb8lRLga3LLWVN5Z2jPgLyXA69g7axKs5qTl0xhq8o
yKgleynwbF3JbEOc46SD39m0FMvsYYDhoIU5TUzv7aRkFWIoXJuPIKSZ+pKWk9iKEbPNtDmEdXoM
327JNlDST/8IR42FgrrtelMuKlR/ko3zsccsdOYdj+ORYLpzVgrsNmb4/RdHotPnfNGuQAWY/yIN
R7OqUeEd7+fCdqqyUNHjqUB1dyzez8vKAlj/hhrEk4JO8/MSU1SY9aSmkOUKawXt53WTsIzG/Smz
ZzoS3I4sxSxporceRAAl74YrdU5lhLeN8aVLIfKdriu+M1DsKTcBKJtmKE9kOQ/KzlSTJ9AdFTrL
7nWYZ7dwfoKgbRXyOT4/YZ27PfPoqk6XYXvw1wVgRXxL+nofgDYvWB1RfYq3jIHDcZcUs5af8FJz
kRisKvfSw/TsU+3kXvdbAMBIy5nIZyCKdfj05/UL1k5mjrOg5sDjTs4XTkdmJnvkbEWQ+9GzhDsS
xsbT17oIXgZTYwEch9Bi+fktw2+VH5wHbk1KU/H8/r/aVGQ3TxKxhw2rBXMDw1XDhrYGDWAzz5Tt
Gb8PezbVp5PxCFLTbTHO7UbY8kTWoyHgLiFNYlXSIue6zBnq7FoSD1irdG1UhnleXkbZ9ctjQLNr
bpIH/Cx7CzkY6F4npGf3MdpR9mC1W/FaiOLoAh60piHKOZm6phWEgZWz29ormI0IhdRu7YiZQv8q
IjixuqFO+sATk8H6jtN/k5lm/G7T8yvMKPMH2FVyfT7mhpUb5yIsnGCebC3Op9WeWbiK7Nsx9wmF
ArhvVRX92OxG8YyeNXGJG4Y7Ffejm7b5LB3WnO5wMcEPevzV9oXhOJN3/t9V65poE7a/gFWeQx46
EbtBc5AzedXcWekNyU1boeGTpTYAVMX0asLrV/tlVrSNp/KD08/thvJOC5YOn28eHjGbNBGURfxE
h/zmiPowmOQZC3U1CyohkPP0KqaWQaTxe8dycgjj/oXe4wNR8ZmIN7aUn6zw8Frk89y45sxDbyTa
CnEm1+4lAw3oLF7G7tXIcFm1jLZViuxEU2KSJ6F6S1/IyU9gHT/P/OKILQIZ88jGgnl/oqUV0+6W
W0r/emAxXhzBJClIJAcAsobU8VMKczs9OrsXHoI8qn8GleqGCd6B8fN05ols7kSyUrjZ+eLRKZUu
aWhuFNeiTI55Tg4/6HnqgwYIolNiFj/YHNzAc980od93mslEXmwDFamXGF8OtW8Qafe8KmIq/kAr
xQPCh5YHH9syp0wC5u/zuN2Udwz3pEzrEhWgReCWzkKeYZseHSAEBnckt7Vgy47UL5NMnW8o/+Ck
5TbhTU2BibrOPw+MGAEyzvZarBYr//xZEzdRVTPZCUM40zOWyPy6CgsO/Z4g5F9iVnQtAeVyu6MY
nJTJau3Z+NpfTGOl/MbDPtlA3RdHiIInAukfcV+IQk1KjbuDzkjShzMpL3LCA3Wwf6Jw6bSVmNCu
2+hdchFfafJf8QvJ024j0a93CyweSqCx+5ABz19CMf8NKbDTPobTUwprqZZ7CpM6663kl7eEi37o
gcAeQIriFHI8xsj5HO85tGfLXdv04PH0LN1ivQQymLNtQrsz/VbI/bKeVLEvZFY0ugQ451bhFHa0
7/CF0dhqpgOWmj2fSrJ2/DAj+isy3boqQfOut2Cc1cAgobRhIOgsLv5cGR07JahkUa8TpsA06Ft1
VHooOqpvpskVFjd9Io5YpK39Tscb5JOFX0hOk+CbQJHn7ws8GlOb98LJjymK2suvENdiEAPq7ayj
Yrt4x95QFOnlexq1AqDxgBx0i9Y6u6hPjf3HvC5fj7WH0YxkG76YqzWROLZ94cJVrNsK6vX9EEu9
plbJ6nUt8YtXORNJkKBfDkiig7T2uTV99xKk0kgmxo4eqP0sRJ1ewgR+qt7lmFVN3L5VyjNF0xQ7
QOybLaqWcPO6mTzD+AazndVYEIqgsPa0ATtxFaNl65V47ZNJHRgwfwx/7z9ypqNo6GCuch0t5Eox
oDeMATl1E7obUTOZTJxTOfVZMm+4JI+dr2H2+Lt8taHZlstB+iNPVOtHMiGSd8UwrwH3G3LDFEAP
h9DRKx7CvfW5Qh+/C69nXPekb166/+I0Uxn9hmAehBxlyeccRnvE3qVWd7N6+esqptHy+ZgUPbnL
JyrQBpuG0Q+vgX2YDzBS7wo+yM8V31GQblAEdwNhy9lVrtkU0psbP3ZvfbSjmnl4whQYuaHw7hzO
H9bZaxE48p+fosbA1Pjd3gf1dZJIqKfLJ8ynWWLvzIfaGA/ftjSKvngua0+u6NTuLom80jTnrFEt
zAIaTI9dF/BGudJUmeZYuvm5/reM/T60EcgY2HdRwaa++eH9zKLVTPgc2rMcpJ9L1ZDE17OqnUPt
XJg+3Hiv5nXvv0YxtcbQiph8KcM02wqcTkx8Z0ShfuTOa1l40PaCCmpD1W4h3mQoh3i/bNBxb8zO
Z9UuQzMt8VRtXUIZUhuu9q01Sw4ao2x+KziSqPmQqg5ImDqjeeb+p1vk/j9EFXp+Kv3mDf2bpglv
n0K2A9XhVHb3N4l4lrYBG8EBxGjtxJl6bN0nEjGIQ7P0HURKcyDsbAwIrVyEDPdr69pSiZ9qZZDJ
PYR+yMtAUzCEasbl2710HCcKrGIWuSrH19+kjvNVErFpzgYjELn2rBzmHQjh/Svx4nKRQNpa4rSB
FUgTqqJGR3edGnoWXsYK4BU5N2OeFKMLPCQO8aj0PXX2qJbC3gGtp5rwB4VZDhDEHy2JhtVpFlmr
Ju0oE+t84CmutRRqPJ19vreCkoAt/508rWFbxxNf4sw+V/LjPc7KUNnhxaecy4+o+frjgaVB3HsE
Ecl2st6Y/MCfuytefDX8LNUsIFxq0OUzZ6Fb34CE+vtaDSHoGFahzCqowXWN6IOMrbNkKQ3IfPrU
D2/CgzptJ63o4+MVIx8Mf5k7WfhCKS359R4iCqrBucDw027y0nUoTTpYL+nvNxJIZA9SBzIxmUkA
GQHC2aygFvDmD1h9vMH5yX+rKdzb6ubNFPES7LCYQvx487SCNUz6pXZ71ZUvlS17jXpZTUvHhmCj
+ItdBVD8l2y8lbau2tZS5zy1BphRZdK8jfU4HP7S2I9cCs6/9LFkBYgRaFy5sT1JZWR4aYZiSYvU
bdR+qq84oJZIKCX02gHi5nXx4WpzGiT3cldyf2T8KYY6pghQnCA2Mlz6ni4HGGrVqRB6DY3zBSQy
34U4eqJ8ZLkZxawY4qBdycsbvOPZ5wbWl+nPsG9WBdamCAUD8Wg3V65EORfohY+11zCxJL8cDN6p
i/X61lCCIKjGz0hGaWyUMuCl7pqfdTAHlxYXqlQUP4KWIL0XpaE6c+EelPbSN3K4ssMW3ISHj3t+
s8KeiRfixJh+iuNbrBuypf9DYzLeNhs4lMK6FECVJ/myIT3CfWKRVAAb7NEqTSIUdE+bhDwdmgtx
WWTMBvGI9WPK6MWzHmX8mh4B4/KUQ+LVclU/lQeauheVJbv8uXGAQXIfLNuJlHij/PUgaVzIBXOG
ZhQVU/ghxqGrQYMPoWFVY19pms6xuKBJSaB271e100DqSORLiU/jwljS3sTUVdRT2oUyhjRP3jDf
vkOCRbenNMkkajZWLZ0nTwA2P3RHdao13FNSY3yoxe6Fxah2CJUfBSSWLQRZ5A2gAbl44gR/1PDV
QFtoanYWJ42nyYMfG3g+RrVOWmC+o3JS2rDQN1eS8FBRcu5MqBGaQavOe0eyS1MaNjeTFSAwblZ6
+r6HGa165U2ZY9DVy5w/O/TG0ZUyd7bNFe1ctf2dUbTFSqFi3QjEq+LEOKBxqgzCpKpWrHFm0mak
r6s7KUB2UiawWbNcAiKsJE82jLzDgRAdOXo6b5+7FS0svcn9aSu30EmnIeHO5yQajOL9EYleXWzr
Re9pE9Tjb7kUUMI91pcGXAHuTUKKJ+V4qo4boHaPAWOeHLQOCmX0JlQJlXYuvBcZRScrmyzXFUcE
n4dk7HDF25+txVH9rqYh++V4xmixvWWgJlU2PFT2hcpmqpF7uxgovXjq63IvIuSLafN2LteJEyNV
9qRlRAE6osQqh1vUGso68UteGrRBhr5WOJBWWd/fs6L+EpyFyX0onYHlwTy/PXrw+U7NUWJneTZE
ofzBUqbbLI3mLd1JZpq7N4LqMAzRXFoYokt8jLCuztmB/NMGoJ+ZbzJ4jT5pN3JMo6oFvorzr7G4
5DLqZcs/v1Ja4DXLYsQv2RI6Q56wXvTgydg5eQUzIfd2uDCPZPxpw2fWWz2PbEoGzIvimigP8fa2
F23CmkqsGGulY5TYnjVrtmgFXGJ+Sk11fhmzDwD3q+NoT3IcA2s4iKl0wCagX4FASWMea5t6R6X5
py2EtLNlzi5JPpwOkH6mos8agBvgUFMmQwCHfVazaW8nyQ6EClndxb3CYwSASRqElsG0VhOjich7
tvYf1lFZ/ml6cogxUu5ntgU6I5a8JNCpFLd1t2+qNvR4jf+7Kb9nIpGvy0NaqRuAE3Lcycnvadrb
etSeXsWVFfMVakeAhzafYiyI50lXu7vMI+IKlNGmDPpkp9dnN4j684ZzJPEwbLctOry8uOqgq3r3
G2VfBy6sKagy35dhiy/18viV7nMGuCh8TXgjRBCtabsIdtv81FDGEj12jnoCLhFsSKmdgObAxzPe
Bf901HMdHfMcm+MW7BWUEP9UBbifZeEJRDPpZf8LabA1ShEmbpZF5BRI5Wtt8VlPdiNVy7npVGkY
dEaLKnZz6A4/GjWoE4y97LO3U1So28CAtXBz7kX+FppkRAqXTcDo4wwGxuDT/ZNhac79tU4czq4E
y0tG0y4UI4bVOTGc0LPfZ6JlIePApLi5Wq9+P++90Y9gyStg2bITsb01o3SiytW1Op0vKUwYDb+k
0Pam7lTPrUHBzi+PBf/npFTuUIxXF0psaxdStvb30proRQb5yndXC4gPkg8mHKtLK38u7seztw2E
mf9Fu3nV2Sg//UszUq8PxU5CKYDKnIgTH83gVtFwM89wX59ETx/GSqUqFSBDSJeY60y/tQG0qZTm
+e5cqJXTF2gXEwOCTNn4HuRrWbZ9XBtMrVD9sC0Yk+CZ32Q48jg3K7/fkyF1MEcIcvfkOOaG0b+L
QLZm2pPUMA8BIBlgZEUj+44r0uAyv4ys+wmduu9enGcYX1b6B6a032o9PSzoGMlYfOD45dyIF7qt
GCJJF/3OAWkx5zcLsVAnb+DZKxApA8/crBoqDhGVo+oO+GIjFKnYAptJ2/RNEuMx9npoZ1WUYrPX
3WKABlO+HsD1v+AFC/kA3lMm53SfypYyQ/JjMvrbQzAUw2F9YnrnxEBzaRVLCskNgHMA6kLevdHD
kvRMaLfIDGG3uKJvxJisZKD+Muy1Mdolx7e9pSaXXHOPx5xRW80t4t+wVVpATyTUVSF5KnIykL/q
6V/kUgZS/yE1e7W7d5V9mCM26+4nRepGLCMoJgdQa6RtPsqaAkhas8lyGBEtvE9CluUDfenH4ixX
6labitUUx2+DvLgQV9dMvwPxbMQm9SIgdZ8jzMr0cjjsLQszZElVBTWtUn/GswBFkEDPDnLvE/on
HaCRp0/jpNU0LaKb0K84JPEJYwWChR3DUb1hAmgT1+GA9ejPuMH3vUYmMj4us3Y4j1iit9HD0aPQ
A9onzwkhJVL+Aa1ZLtU48A8py8d4giSG9ThMTK9Zyt82YtRyQ1MwHbXFqv3u5WEiBdH34OUEOdsa
z+X2/taJScUhs6NNqw+hIODDUW15uwXCFyYJfZk1fm1WY60dS9r+A6gOD0WpzhVOQdtqgpoBjp9C
Hm+oGkXJCXv4SeTFH45ps+0VTcrS3qpPhRoEXJqRy5VhVhnOFhe9Z3x1L7eU/KkXysiQfSPHL2Qd
jllwzEvm/qB7aC1z4SgvuwXS7XbXmkgCjpUnzHMui5Yh8wVZeo9RBg4ZhR3BLcVbjZqg6whr70LR
58uO2AD9kkiCMQjpaXmgltoA1hilLiTre3T+xYzhz7eKPQM6+Im7sp+Nqe+j1Z2aHKZ8uBaBHJFs
cRmTWEIcLfw5dckq4kfK/FUhXi6yH8w9eauEC/HHoB3pCqHIKtmmRmPUhzpD5gtOCtHf5sl/s/69
c29EPr/W2dTZJgwBey6QsHSkYgwRPJpoIKQqJ78GW9b5zQARmi53zsD8y0pF3eggsGYdeJuIl2YB
jBD/WkRC3obChRl6EKOMq78QNAVE+wz1Pz1bKyVc/I3jMloeY0xdqLJw9oUaxnjZW0Mxu1yNNLNh
dNq379iWfst+cxT4f+jJwvGjze3p5KyUNAb+X28+0zy7X2bdfQRmIz3Zegguu00/bXMv5cdnf+TQ
99Q2HnVgd9N2ARUae1pcrhskrnrvJEeRGRsm10vTaZHpDkXCBzvnXQb+yjtiCroiCVs7JKWsn3NH
j31UdO62qK6csYmZ+Gg0fXTCEQgb7fAyP0DqjF2f3AITwuWR8aqvkF67LOQDehkdJyCF8BChbBSJ
xAXZdw2YSfkTO4Fw/VeDAIvnXvYlhEdGInOi2VsiTeEqYUCRXLIt9W7HoP380sB9tscNbO/MXKIZ
WFU4l/Av88hu0NOadUfeljYL5KMGa6srnjURaNAQ6skDV5LSbV5TGP79BNRavNi8zVzEIOPXnwUF
SEoJLW77YL5xija8soUAvbbxonc9vDWUphiLJHwoT2b1w5NlO2+d8/wpfyi/CzUoDSpF95+JlRIp
At17jkPw/r77lBLMuybXkHFG+IC/OWZKIjUHxTBhM7PK/e841x2C88AHA7p527Vz00SLhH3g/h4C
RTI7E0zE/Upn2bqMR4rJgF9TA9l8ADmHAdOHCt5rfzu2HGnvid17WvzCjXEKY6emnIC3Q1O5P9yI
ZKg6WjkijcmyD9xcaNO8BWEn45xd5ViGj0mzxsvrJCUuzBVUuo7xZ4A/qmsR/u0o4GTlXMHZSpvZ
Xyzh5F0AdxJYD43HFGswUogF3Oa0Kmig+bPATHAq+yTvqSTm+u4TkEO4CwCPw/Osefx8jg4KW7Hf
Vo8J3jpXC81Ktiz3EbeMWtzYQhZgL2Ub634H/Qe6WYbxIQ1WAIkVY7mH0Y3CSEj1SouIh/vAGTyo
yh7pbUoFKTSWBraQseWDb9a6YeCylOVcnt5c5zqQsa2LSvLgxcCr9ghMq8EAEPq64KAWWzxf8R7i
LFxGOi1UysLLSrY5pnvKfEF7Gsc3AReHL0G9NI9yuVZC2/fQh3rBP59GCUbek4DyBWj5aS6wsak7
te//xk5lr7vVHpfFSFSak0jRR8ohKQHyGjwcTREE6aW4+o7wvmxZoJGH1YkWd7S6ZaT7bif3PQ58
NEzE7OxqQJWddkakqVGfhPOFgOiqpNSyh3KPN3nBhDqJk5MbvLPh21Vylj2GRqsxBUs+Q1jAVgiy
MhS6xQtbHql3lE1NPuCXBNN2CTLNhTCPdQbQqpEkq8aQV8ntReGbjk3SxzC5rCQ2LGuSPDoq8pJ3
gbAsJh6dundWJ39pxI0Bara8VLgycAViiiYiNOaLOc1l4WEFlUVbznp0zZfIAjQpmsLDA15ST295
BEIZwAP87VejC7+AlOKeIjMtHZp11a3wNRFvbHEQNGGueFgpQkbmpMrIYyQAQ7gkwd611B6ndm4c
V1fiM7Q6lL5lSp83lY1ilw3Di3Q/gmqVCwkr2ulLbptRcoWL9EOp/Wd4Tmr+2i3mq9ymby74CKdc
C9zStLFe/SxDCQ8Aeh0SB6u4q2sUli7csVZL65BAmUkF3/Zj5gczO5QcHrUOciCi7x7nRfSp1Ypj
4Q/K7IgnnMajnjq+6vsDMxUgrtEygpT+rqKi3CdGZ2YpKueoiiY8XILjl0p5+jp3rnwgoOzQauBE
JgrbzuVrg/0Vc7nKjykeVBn5398muNfzLe/hNnQRH2fHqUU4HSclT96joeh/rhVqguA20W+HMbs1
Si78fNDlx7RXHgJyFfu8bSDNFPHdkhKAq3VM9RBgbpXs1slsJNAdMK+ke+3xdRj5esCwcOgp1YXk
7weVeL7oQRwU8+pUXq0AE5usAw07HeX0Rh+mB7xYYmFxLbOxEDLunSwgS7aXLNbgeNgDCHoPA2oU
jMQm4sbSaQqVeaRl0Oahv6BmrLyVXJUYIdkyuaTFlwVsL2EJFCDwG4a90ZrMtZBR0xeSRrV6JPVm
uBd377IQLSFWEuF6nV7Y1arC5xXgc9Mk83u/TOEMkOcmpwAIATA/rHr9C0fBpcrMT2ZBhLXtpDgb
wu0a+9dkA9+FEL281o1wgqZhwDWnqvp4I4bNLSPnh0bF/AM9LUnDAtJcXz8QwUT4Mt2RgWFJ5P3X
cXpOPKNr/q1tDxbelTaM1JGr/Dbxzn52wAGUrD2g9GZqSoK6MOV9e19KHQz8jZJqxRWn4RV+wlcU
BiwFr8f+NjnlX5XmMTOuxQq5TTaflv77ixEL/qoKG0vD6mK5mhbiaZwrVS9H6CeZr8bMOD+GaPuu
fTjJzgP3Ug5g3b67WZdiWvLe68JG3mL7/bnIBqjofnn2AeNBfNO2dAAZgRKwPg71i7zElQJxCAi/
fTgs3tgtwV2MJURbBwbIC9zDBzbyCfu4xlTUHn+mGImtpSIdfXNXprLSpU5LEtYKrjb8pjWuoQWc
Vo/yIB1Dtvj2ussIzfcmTRFjPKxkySXhLmDg1s31l2ey0xcTAvjGd4e5JfHzJr0MchncNrXVifdF
/Q2ESvy0AjXY5G9Yhrgr/RtkucuPuTUC+TuWFDW2PdbcqmZ/o8b4iEDt9tTtJC5PFIfXU/0bJKyk
tqUx65iWQrGE280uijh8cfkqz3xES2h4ODlwr/cPs1H1i+3Ug5589L2PTzPX6+jHQvsWtt3qQ5RL
dhax9gc5XHezLehYTTEbt0HPYi17p2C65P6jhSdX7vdQyyQmnGT+x2uiOOipVolE0B0HAbP8f8jZ
mg8BTThNpgjjcelHGgepQHDWVNe9Z6P2ilGjf8WMmmv6oy3ceXkMsNQxg+IMJ93z3oPFlVDj7lPp
kkaZl9d83diR/Qc2ywoUZc4zzSdm2YPPtSC2L0sQZbxJ+9/j8CzIvLcSfJiKwQFOUdwIcoZcNjEZ
2g0YOaB19Rj0Ew6Lj1e8keVJEbRjm9aI/3uAkxlHOd9GCQ1iQN5MAZEKZ7vivPxOeyQ+sdkrmx0t
gKRPFnMbtYaFHR7xLbTEFibnjTSJKA1k0r5lggTs8rc1JxWtwlDrQlmufVNhkAjwGSsd4SGWmKfi
5b0EhZn/zFqxGxj0bLjWkEi5NsPhgAJbPGll0TmGzjazijj2EvRVO6mS+t7mxQYVTzapa71D2QSN
O4iGHlCEaH3ftit5FqoNjOlpWqg1vWFYdx9XA+QnGTDhMbuvsGGxlVnd+jP+P7392bOdiENZHwiR
5/aq32p9Itv3xXrkVovMaKta+Wh1UuIaKLlo6OldAFT0xnS/0ajccVrtK+OwN6H4ZMFW+7ShA8Z9
mZPK2w2o+TpV8uKNTfvXwt/A/spklaNGOisAcNrNBIP+tYQBtkQ7K0n1RehKRV2mI7KO5J0S7t3r
kQG5u/0ptOgbp8a1MA3UqYphsEPeXNbttt2CDx+6QR2uxifGd1ePMhJu6ab4aucArQo0jZRv+GBu
Hw5V8oM8jpXhX/gtk2aYbXISpNGqhW3Be6BhKhEzhJueWztzO+2Jt8WS4FiKa/ep6NFyR57VG2UM
Y5zq1fSwLZXhZQsOwz08HMtuL4pIHiwJy0UhNOrp46Z+OX2h6xbS2LM6jswbWhb3UUwGt4NMu6P1
bnzTFEJcyy85pxqQ45dqSd2GP+bBa3BZtrImK2H/guSkE1/gtkP1gbxcdZCg2fjCerqdPBilCNUv
8KbcKBOomGYun5Nc4d4kka/8zaIyUm1yxxtuQi+wJc+kkoeq7euBw7qbIDb43/TGeSlph7iy06gP
WNgKooiLPaMrYaHdr9THNQ5sY7eSbDOa7lrAILZu/p0doCYz29DfUUqhQGUB83M0NNgm0K4YGcnD
ZoG8IlSmDvoaAMvxpJu0tOMmTEbB6OM9iJS//kKms2dXJJBOryrdk9VxyQu5pLTc5EmIGiQVstgn
bm2jPuS+FGvy/ptbbaYIoujDtvKh1jeWf3moZTgnpnC/udvfgKzY5LHBuQHWB4Sp8EVSV10/ffyp
M9GSltwFBlyaoinwEEOFagKjHxHSwE5M0zKmweC+dZe9M+YhuIxxlURJ2RQkpXne3ek9xiIGUT4o
I7jOm72rjItRI3qTLSnK1iGEpa8gPkDWEFeJ0RfS8bBpXAVbh9DiMcO83vv7vlfEWxC8Bs465nYP
SSk4sMz4zsoZDx61e0SFbJ0viUes/0RqbciGZUyxBPUb9gqs0kYWO0P0lyNcaMcjwgMNRxKYVrx7
F+0YcgUaPydsA78BqKCF2i11kYmoCJCozQvm7qzr7ZWCnEd5CN+pveFjj16BOfHjyaSLzNmmGfvo
pdq0FjMe2BJKVLz9+5iOQ2jOI4P6VQs5pR18jMc51HBZjY+2Lh9zF9a0uOt1tb9EqT78vq9hr0XM
IXGYwdPWG6+0d8tZCxW5kTSRsu3pmskQVLRUNoYHlnvvEXG6t/3ublB7DF4INES+27Uv7UXyl7U0
slLsfcjzU4h8CAlPkKA0t3+TxtpxGVAuUDIy4/QI3fKvNJyjj4A39JJijOW0d5p99SxNyy7imib7
V1GUtb+aj6HTW1Mg5iYO7NZRvq49icAcftrX2cUH4Q3iqHNB7B87Ga+8HoVYwQehyEEu1mu6XmGT
XXZ77tXlYxzSle2A6oYJlJ38lf7XtAHUA+ZNfYVAxxPhBDChlUyxVcytU4oLu4eRPARwtE3PW1ld
l14r3+wxjNfxnX7mRoVPlGCwaY3RSF8Q2zV/o/NHr9lZdYCqZcQ/0OEiwL3LIb55BMYe4sbVFd0n
uO0fzDQE53zSkt2WFSlZR4W5/fccARplQeFfhzOmh8txUeZ4f7T9yhYuITDgqgueqk3VFEhVLS0J
/c5TdzvXirWduFMnzknBsjx9AfGzdS+v2UzEok2q/JQPUAT368yPtbxHFreLF/92beoDXZFB0h6Z
ec85pwaewgNl2/Y0h15TILpkXz4ExR0hO5zxJcEwoShvQNfM+9RKEigDPjRA5Hsr8WoR8WaQgs9c
/HVKZLBuNNs02J68Kplj2A8x4SdmpQdi5hONx3o5uqoiNICtQXn/ieTPny86wMjBcV10AdAnJl8p
1/cHzSUMTIVtL9Y8MntcjQIlQOFjO40V6nFT0dOGX56Ap+KDFSmapq+fG6PRRd8bqnt0pnHY1KDL
kuyYZBTlujfjY9jmkHNsa/N6JRVmdgvMMg9SkrufyEFhHyIm/kpbHqznCiXUOYH4U4iWmTU78dHT
ULNEiqSHofe+MU90arfHuoikY/EcUqQD4KhcPpd8g3vN6sYd8P3nFNJyypxvQaY8FjJGRukllrBe
wTUAk1swUnDV4mSnIL4uJyEaF8BC3zksxmmHK+C2XkYL1ODJtoPbM9a/nCge5FhTT3gsDhaTgUrg
Y7ri8doJQEA9LrMy/h8fzwJuDvpkBbmLCmuSi4g2bH1JncG8WqoZ3tPzbkEsJ5o6WvabcvSyhYtZ
h+6L9csGowXvjz+8YE4oQuCg4rj7GysNKoiWzJvkiGQ7ERp1Q76tWkV0vJFpMJLGowXvfgvEn4DV
znIRbh4MFlKIR+A11Zg3+Hd18b4WSe/WrzLSrhqVCf6EppkWAPX2YHS5iiZnUz7PACETOrWRLJHq
XjAeWiOXjBCXdLDxfz2lNloNuoiVLo6Y/DebybmXeF8/gQuPx3TAWtBhsij59TjUo6z9r6w7kn8r
N3XPAY8JaM50o8zvsDSvfCnjxJx86fchHA0gPZK3b3b+a4WaPZHac74kc1qXHu0BqOA6LU5wXo0N
qUM9lSa8kdM27NVWnsX7bpiYg9z6K2GG0l7adqMxWn6ygCUru1bb4sYXYyzjB0NBgK/AaGu3vext
7tio3kHUXbLr7TcIOHQCQXdPxtT+YXo6FgcUm8jyOy94Nh73pEwtKI6PHRKMtxrSlcV6UVHZz/kw
Ph9+uoxaoluPScotRf+W9uBQQGVkBSKQoQDaBsbmOEUYGTOVbQuq56OqIp2XtliLadwViqFiniQY
uRb0RCAIblMz/wuak5UUsTQPPijZT84AZFHgcRFw7y2Tn6smOdPIhilAO9WQEtpt1tMWomPvHXnq
o+f3kzKmv6fcPyQ/x2l+WRDeB4X+fU1wtFH1vDM63D3/JRl6YP5j/5RnPZbG8MNidt8kFGIdW7p9
AZ21Nf2lDGi4j5HmoHkWxdxXYurgDtUXf5SBsVe5h0D341n9n+GrgGbK4XV5vNQBkGtxQYWWKCO9
Zk10/Far84yGRtkf/+iTmO8qPiKfxGHIyT9eFsaXSiwffUKqtd+jzHeruNnaJ4EKekUkNCYOcaIo
+MpJqwwm+FFUpcmCyoVfyis1QSvOp5xwos+xljkUkHcDJcK0wYy+xAcoJZifn6rZuEL0itqzrXCN
jaauHGCuf1VFsW2u2s2fNbRnOMSdK2oJKRc6nehGN0kzxXEDvlMc9so9YScV0ryJ/JIgkYxo1Ihk
bTPhRz0aG3RfIle6YVpeDGzqv4UwGB6tfXoUXomCWHN73SwlS/u04pEqTLAtsneyUQs/FamOIjgI
xRshLImTZ6UPqwxEGPaFUo6Z/JpJCxfOtjudnxfo7V2D+nkhCY5oSNpjBEbOvvjVgDZKttkpX/jp
dBDdqCJWIKpgbaC5yUYbEqOye1oQxAHamsuT21jUtBcuiUVbcvwy1vaaE7kSvYIGyPceKFtBUXj7
UMqGtmfQ5n6bWFV3MsoFOYSTbzNowkkzsJM54D60WOsfhbQySzTix/kSqpUs8bGTl35cBDRgvyeX
0nr4sQYqk2O7Izvz4uWGgziht9za02DMAMx/eo9j7jITvqvfZcaY3FYPnaKiXPX4gklyc9xbytFn
MpAtpE58Bj6JYWfZse5kJjltuZgiBcOT2fOlmyFgSJbGCSCk/h7S5vKVkhJNWNMw8fl/knOLciGy
4lWuFd6W72+ZJUeezFGmg4z4hPrHT6T6qbo6ok/ZkXKyhBHGAeVri3MDaW/fLUrvL18IaGw7ixDo
8CK2uK5IV+8gzq0q8Mem2kyuXtENXgBQEc9iEKsjCa66mVGuj7MlU4YSq2bLfBjfT0J2Veub9EYV
DtFsKTsORKowA3YhHvY/duZyV8q0XayxROq6BqQwHlKcv41fPiWu0u5oSvINOKGBiEUZGDMjH9wY
MSlj6Kum6aFXV4q3hnBUML58uNpzGBWWT0fIVQMBnETPcNr8YUgXfkpktbEgelL8fPTZhrgbKi7K
ts69zeDc0Dzri1yXSSm/3kjlSA4ZkoaH6btOYutRPRnJ8pn4O/KmuN4YRZbVZozCEAWup74GNPdH
TGz1QdfvOLu4ILTIZNkK5FMRKDyum+MZUWOTDwsAZhGzZCgkb1UIIGxefeINo6g180YeTGGJTSbN
RjhsS9AfwFxuR1L2am9ltwDVmhFcHk0lqt/4IvpLd6HnuujH1ZjuDME+9bZHN6jFMBRJdQRyiRen
Ay6jDpiQXkJAMB+lMhKmquLqJT15D5fKYLRg1KmWK4H8AqgE+RVXBIozVo2SH8lwHiw9mJs1S+NW
gUKGzyktM4T0sVcM7FtpeL6+lD7Vs37SmHXE9I9L2zfZVUdil9Jn3gGfP5+TrMQKFaM8BEIQgSwr
DBB0FV4Ig8HHmpWkABkcSC7SHL2xv2Qb8ueHl/iPpQxUFcsfpdq6ML455zBUJRgniIGwz3V0FUOm
9tWzyq0qb83nJn9eRKod/7M/KgF7mWLgjCLB5K5uspOLdD9vAjGbnHhK12PvdXn8XPIsV7Th6cay
NxqdvljxrT3dXfyE9Beqct/jSEFhADw1v4PC54fZ2obFvghIMKJkgCh3w5bglUWYL2CqixM1Ctzu
4DTXxvyQgVeglaR5FuZzvNlfAyRMZ/o7iQSIaGAAtBh43Q2udz5Yq/CeByNL99kw3MZpArPZy6Dx
ohCEZHYOnmjsVpvNgTMQT66bQswZ8EpMLdmRCqIUFBCrm6XMpGYzMGRQdtRiPNlyITR/YM2zufa2
tkXCkYPyHrZwe2KV7qx8H8tUYIfP04Ka21HQPl6ZPSmSsBpvmm4xo4nGdxtvD0we9hvrk/ToZYMj
yaghjS2EEUBRdDbvRXqejetMoPtgmh9Aa3V14YyZ/agsAjWqXs6chwmGQncSaJ93W6UOEAUkyk1v
z5Gw6Fp32XeieGJhiBnFsAhEe2z+8GyG0qtEAmWnOUyVevLUfcpXljcaZZz76KaRZ80B1WRn5yvY
ZaGEYLZOZZDV2T/urMB0huCqPLy/s6yLRkNbvnfzVNQiAB+1yo2CBti4AjucDge6fvPR5FD4l8Tj
3t/TvrXDkxGxUsJvYX+AK3jM88PSRXeOqOF6/5hHNaqEGh5iKhbbpw+eCXsuU0k1WWf2OgST669x
bw1kyUba0BT0Wke8eQaljNo7s7PiCf8zsqrRlqIJKn7k8QFPeENHhvKWBJc3LM1NVsW0jPPXM3pH
hsh05RUR3Nz+DEKDN/s0cJSIBtfwM1Js5lTTiZJdUpeYo3a/xir87r70c7w2PIFMYRywcMy47JHn
zqmB7R4LruiJ0EdWTl3aT0ki0DFO47+BxSeVfKsicnaksjatamzWfamF1+kylJFe1HHqdp536ZM0
3oGpsmpTd5qZqvE3U00WBrWIGJFfU/WbI72XtLdG0Rm68Tcd2sq9v4guSBwwb9mKgyvWk+YRhJXg
ibQerKyuxzWTqXKdDONA6u0caXZSfEAGMuwpdL9duMXrEHQICuCles66zoRKqsMALrqjxtwyFhc5
xtcUlOX/qnkZAe5NLY6s864I3NB6THhoTQMEvMNewXmwmhOEKfqlGK30KGErq6FFlcqExKE9sVKL
e0kBCPRdMoVYEzTMd7gwLXfTRJPevc3O+EyjTZqOejL7YeleizmbhC/lFd0CRCn3epIo9OGUVFlB
HwIAo8ky2sE47jrrfqJ+6Um+j3tdYOZlKYWdiTT1HzAWexOu9e4M9+VfeR0moV4LNIK2BF51creK
uAZNQA3TybZIINYkTa0r16u6RdvVOIfB4M6HIr+Uzpjet39W/2dqPir+bTJqhtBIvvdN1fs1wj3Q
Y6HbOnFAR+Ffm8iSgaOecukknanEKKjofxxbgtKsvNvF38X3I56IFI/83E1IJaGZG+8a4vmFE4lO
ycjxhepwoM7j3a86b6hyffAsHdrskYEp42ffeiMpodWZa+DVmiWRVWf5Gyi/rrmTPokWM1zFGk4B
a9+bExPDOJ2PYYRbv8RoLxLvh8wHEAWH8123kvWUWMQ6pa0tfFxw8AInAg0CjrcQ0cFycLytgpGN
F6/DoYl+9SwLbmIGvntjgj1kacl/GdRJJRQ6cDbJnLg7hlJSEfjWRfM53y3+WgYqpldKe1wB9vw7
linYvdMi3zH5hY1qKCVYSMpMpPzQTrCCBQ4Rdf2BRBPPQ9dnCwDIpSh6Km3iuLNN3kGOJi0bG03A
a3wn0WYoFspQ4WnlWyQ8futWCoQJxPyv97QPBjFR6RVJZOci6MA1euKg5Veru0TcRRGnOU8FjYFD
88mZMoWFmuQwgrZ7h8tnBpFoLJRdmUz0apa+3DIKKWbvS1z0z57vX3wVtuCdzJTqUFWLuNX5xf1+
lZnAJ/34cUx+nV+dLGiDNNDHV/3TCC5bq8+zXx4EQ4iwH+bPRBGiWEFVdPh30qKgX4WD70exRx0q
Pw437k2be2DxxHbnbLYl1s80KYC8Ztc/2he4XAlAL2Vm7ea+7PeqSG+tJjHYcnwhD3KkaPuQlqlE
OZgj7JENIBRTzG12/0fKr78m8IZy19gy864is9MVqvWSWDB/ljCu+SvTa0EwvzIWEAGTqljhVtBn
S5Co+THHIs14ojV/oJBgc9/4uQ70pdloyrUiR6Vfzd3Jfk8fa/q4yBZzWgsSeyfb20cTEkJGK2BJ
8ObFPT79T/09Nxt6Q+ZRBZnZ77DFCTGXgYA7Ls2r7kAN+1gS1eXST+4FteWkBMMHGG5JYs6dF2VV
DbPSuQr7qyyPH2op+2c/0mG5X+J7G3tPI6HpCWa0m7OUiGelvec8PmRlQqniYoR8PApaRAgNNPPT
S3ZNlypD08+jx5YQUGY+yGflPa3h0nD2tm0ldWTUJvCQV/voDDwQCUxoE7y1z6KwF/AkSRDIPAJy
syuWXEBcWohN6bIWhBGgZtUgsS79KyaDwZSNmoVTXdBQtWm/OkW/PfNIEvAJsOkiCVX+6tWY/82j
pZOSxc8Utx45SFmnEw6a9rpS+zqpT04DmZymW9GiFWM8ivtgSWguVoQQiSZEr586eChCzH8PBpMJ
iTra8Eo405gSVUBmqqZyQABQc/P32oHYQ/i+woxN6ldUpc0wZs+zRW6DiWIa9pIKIo5aQonocS6z
RBX/zwxJ2VAUDqg4diWfeJ8DJqwpePlPN0nl6hgw7sUWaFMGfuNZWjV9BoFmH7vh9GNsYmVD+7fk
Dst4u3vmo0APwpF9MvwA8Px/jago3RA1RuRPTTX8Yw38IWp7Ci6raOH1KuYO9q202OcmBPvAfEUB
vvxPG1mcIwO6qamPx4XLSgXkjvSpb5vweW9yyEd8pcR+/SgQaAF+9j0UCsNl8B4Ue+0ry6heckvN
D32b9mPelkl+lisXSjarnAFj+Z+ETNCPSIdZcpKvSVGRlhXzZ94GPW/a5HNPizRbD21EcjSGdwoI
H2VbIsRVWI3p6QkDa9BdUqQf2AH5fbnnnYvwugNVTxZAcXwWrfb6CkZpK3j3ZdifUkzIrMXPkUvd
pQXtQtwUBYsKA0ss/3IsOCoFKBJYsaqRjXmOdGhNkz8lnqCs0D5+uOt/vX7dmeuIKHym+nsXzIzY
HLPKdxq5UfeIuVacJp2Y5tueKRMaczYpkqNqzKdqdnlGoV1Vfu0tCxtYIrT1bEqlozWQy6qtijBs
WZMRHiXv/CYxL7XpgoT0oKjdE3+qh6IIZEXOXWSQP9hTC9LiUoUM+LK+hJu/zbEBRFrbXQ/1DZ9u
tPwi2R0peEUAOvJcSMhfHinyFoGsWYSW1fOTLkt/xQmSOw2tyn7oPp9biWUKZZz10mUaHHCpz3px
BYbxGrXhBr5xOR1UDzyhZprQ84IjBz/EVVSTkZ04HLprEdUiyZho3JQyCDEgLZyDuRj1zK8IBsfZ
JlroeVgfj9HChXvBqyJtnXjlgM0/YUaBoBQCZUhTQ/PjqHxPySFrgWkXUUd3X9dMGhrn6Yud7p8z
vdXNoqyV8tkTrdi+bAAg2uhHFJUCU7vg7ftGIaa2SPBiHDHVPzwIfP4m/EO+rfv8GT09yIrU1lFj
93yUIaqGfb/j2Olauo6WcrgKyAdXRxDhI7mjoghL3xKvHSdXI9kup0Pl6x2vU4nrTRvvLRUle1EI
oyoiaC5jAgfKFhw3RXng9FiClLS+Fr8RkTsFpYVWn5fP/WGEC+b2ueqyQ1GGve8HhzI1P8al9Yz9
3n1VOo1g3IfK5EsKTF79y8Mkp/xFqdqM++/oyOVv9xfyiX4hRKWC/vfzFKVWn7raTzXL69Vr3vSe
bUgIFtuuZ3VjC0+WSmJVEt9X97SKAy3p8Tz068/sCkaviyhNPU47pVyoPNsB7EvoFMgdqT4Tu6hM
b9Dos8A1B7K6U3ckpP4KmEONyINy0F4d9MT7uGXf2V7kIM/ku8qBgSFYOeIVZVIthC/jtdPfOifg
QC3H7Y+whHmdafD/o7bFN7SjUv5uGGHGU82x885F/I6boqcTYPfPG3+y6YZfEXx9+pxklq9b/yw7
+6boXa/Vb3AYL6v+Z7vL2Zr03gn7kutcE5Rc4hVQ6jG0cGS0DT+70PzUHoi/2Il3OMMV0hvBZVVj
GzEXEP6Ny9oKpti8bkCYBgFhI1hurIGXFTG3KcjtO2byFyt4rqGIzfgZkohSWj/Bbw0xtfm5cJ64
FKAOP2UUuZDVJ+9GUioBMJteauRer0lw3lymZO3n9SOLMzCimMtl10D9Onz+Wmwb/6TB+GBnrIhC
Ex96hdvnFRfv2xHCykKMqPDaHK8Vq648tE1rAzlK53ZFCl9463eOqR4+ef7Ps0+cZ29b9ZFVTLkI
DrARP5C5Qs68WrR2vBCLVJRQP2CPeb8YtkyXGVpz1Amq1JsdYtnt87QGwbiZRLrb0wiSkvLODyN7
QLC1ioUXM+2hmBNSu4ln7NhMhAZF3lqSCYrHgQnMwka+BPJwzRANwEO5OqILZ5jGE5hoJXomUDhj
+IfVAamK9P/XA5zj+D15hbqMmDRyd1d4I9pgc4+9WMzTh6P95jBt3W63gNhetpYYLMa6d4duMuZy
Un8uxI0yqOclGNvSDyyoGu8/cVNNd4hj2AHMMve82OYeq9AwXy9MAXfRA51FN730gKaGkYLmafxv
epF0jZEQJAKph0mwb9Zg9F9LobLnnhiuqr6k7TTppSi+2QfluLkLHzfEHjiiDSmjYh2EUXLJVgoX
WMfovL1WTB7ffJiDUZ91p7LjyGT7yoD1CWrCVEnH9iu11rI81jt6v/PNTVF5sWbj86NAmniOAsD6
4m+tJx7pfj/7CsBwqvD+QeiiGpjt6xPvUQNJv8wa4FH7vWQD2K0wl9PQWJhJz5OTPVP5j++M9dC5
XqYS8kIsmc3E08iin87nZucvZXhtuJvK193RM9p/sxJd5u/6ky9fgJydXmA9t2fW3wlgvxJGWkYA
8WO1FkGd5ysz0SeklhfRBS3ZHec/WcgAa/I2Vh7zL7df0zCLkvXizdXPINza1TDYY3Yq+PcjIIDt
hTHFUpF8v1GbisVYiuAAH7r1WoxSgFsTHuvmrJiu2zyMVIE+kdJS5/cs3ovozI05e7lObVeGbHHs
0ndM1/HC8TY9c3huNaVPwxVCoVkrnuRvXrhmeD4CZ5Ubh0s+4umAguck3NGms9gHrjLeeaVMd/co
Z+AApLJhG+BdhIo3V2NYfOYR3WLlv/BeIZm7+wsp3mX50hKdwUzStDQk/nQwGyHORUqW2k43DTY/
E6axdkkDUFR6CvhIPsdKaiTzlO3EmJoIXYQw3kDIc92SBj4ZSCGYzpGh9bboot9R32LU7iIMUWV+
0RzGqJ20qJR6DrlnMHhOfNCjHdBP4aHuJeYGuj6bDsx76tgeCr0RaxeWf+NE4DgLKN3nLQ9FHu0f
m5k5R/l8mXzh4lPc15IM9+Wx3hd4MYQAIK6StkXvNWhFYb66G2fMrd+DqaC9k2y7a96z71Fgh8Ph
X+97I1TNhWWAU5oMV75Yhg2sKizRRvKB8qtdQ7Z0umzqvK6W8KQcWK+G7YRJbNpVYTSLQclCpz/r
HAtFYSup2j2JWZpc9WnF+MQdClNVRuEQVFbBhU3Xvdg4ydm044x9Y5i0ax8SjifdChlyAw67U4aA
HUc+jhqSjYUTVjEFSCpwk84B0ws9LkPby95u7FZjA2ZOf51ne2G9uMMo8GNaoQJDzF98aBvatdRG
W5Wgq+u4mItbisoTCCHkwGq/EN5gX7vmxt6Q4ZsiSglxxAZlVgw8iArBY9iZ41rId0cDzu5fi6bb
M1lV9FitwrrWv//D2IhD4XuRIhf9b3mX2x7VouIWX/WIGTF3avHCY0AZpaZH1NwGJG2yKoAxq568
LJbw8ZGvX86u2Kmpo8xJPraALcmVcqsVO21c5pkmhRkHyOOta/Ste8ra5fqqqGoCaAF9d5VVk7MN
nKL86eSG312RnpXXh9p+tGksiG/Tyc0oMqMy4qvl7KVHEMATYKr8nEt49/mb1YZk0FyVbg/ObxU+
9GDat+babu6J39ybyDBJ7ELfmx8IXO3pojlYd1AFDjnqCYYU6abEkHgFXQUb/BOGqxIUouw2V3Kj
e7EyEAnHU6kP+kajuntBIpKZHV+Fj+SIx09LZpPefrW13iUM/IgHR77wk3VKolpeUUT2+pLoLzbq
wceWAE8vvMXUnIe7VXUTUJnKYty6s/ZoLmrq3HyFJJaKYpBuEsoHaYa0PkEwReWsG8QJxKS2PVwY
EVXA2S8Gp2XveiHd+EG0eOZzUDndP8rZ2sYMGKMAa0qgG0e+33etLVYF8zMllpr0mmSBdSdYXqtH
Z4k8eQmAhZ3mdHz6FRLXOgGhPG6thDFcJLkmXBkKPMKMStp54HhzwlL+yUdW4nwIQMwM776ypNiP
vWMoGLv2vs9FkDjQ6XLMBXhje4uMvj9A64OnDrV4e04OB1Ate8bwjsG1Dd1rUr0TYhYUL48v0s1d
N1HDMlxnB6zSQ9pwv0LtL6kzXw1XHDFo4+IYVMxKl9m16nOiVN7S+Tw1QvcWd6bv6MjwrKBUQsS2
XQKbgfT8jNj1W5EgdqSKJ0Ur8TMEgo+Lo8tnM0b0zgqJo9KQ2PeKeAucR9O75LAT2a8Jf4IFOYP/
TSdOn5ExCDHKaQWuYVtk/lXWxXBShciuNG016eVDLjW7N00Z62AF7CAuKRXdkrs6t+tXLpmRnOXB
oSXZQuRrazvrfdajNrpOtKtLmjSwhTJqr5IcdExwliC4nXChba2DuSAmm9gyHGyV+fKKU1VwcQKL
7CP93iFEu1YsBQPzjZ2VYM6dwBiE9VfMLmiC4iHBIcvk5uGvOpVwwQVJB9yCQ9EAv62m04b+XRBj
wLu+/c4zwrQ90S8ltJY4grZQzY7RjvogdaLcYyK4xRUVlXEw78oF2rHMI/UNYZxsLBsTq1SShJu7
BtV4n+P8utVY6eAl/B2e+oRO0Btb0vwtig9VNGIHMQDxdfrsDnFD8n0m489m0sK+CmcLcP0HpZbz
w/tpXWZeSYi4g9D6f/++X/k82RfmNymnJgVlrNiwyrBAuF9hZxWhSbyEwVfSteSQLX/GNtDk3w3l
j+rFd1aNFRuNOfUmPtnEeSjbDcvW8PUHWGf958zkhl2TZC1eGqR+6nv70phZ7+FuLiJ+Wjb5abaG
HIYFtERFrUGjthaPo+XX5+kXu1f08wpMm76ERKY4YmRWG9VFEIMwSTDVmjmK00Mu1VxUCS7/WwbT
QNh1w6+gK4umq83nGbs0u8HPJ8cxHahTjZJL6ll+TNi5DY2tQynjxYxT6UO4LHQcu8JyOTKSCppq
7tPfe6w4YUKF18m3vTt37oKO6uRNujWSsZmdCmRQ19h9dUb/uBcYy6lAUrpZWP61+Ek9g8YL9LRd
NkprzwMwUWOhsicn3XcnAwgNXyTrUgzu8SZewkyqM1ahycUc/1OEkO3H5EWrH93P16RDb5VsN99R
gccqqPz/8V9BqxZgZyJX/uKzloMhNfsjJ7XkBOPcDpDZfFyXkQwarSQUURLgb8ZEgeqZOsK7A9eF
mO7tVIl9QaiGxaHDoBpAoA5yzVcmG5PAxb9a2eypbejiuEUsOOYCGR6bgvehvfeJum64Xk54+Cto
b3Xi7kBtFi9nFC3tKnRTr9P/0ELzPH6MJCFckwLNRrXZJSLim19Osuds1WBf2yd6Tb9YZZ3DqM7o
RvT1Sw84mvO0ZJ0oq8+7AqWQ+1MmLdFcOiSjzgrH4RWFX5/JHT5jdj6JA7vvgarRflGPMQ/r8o6/
y/uTiHk07uUDV3X6bikr3PpfBNBLAZLp1oJ1V7a4/aOJV0I2R27VXC9yWc+o83/4QY3ql9TMeqTL
oFABKjKmypaqOTfyZ+iVuaFq5eT38B1ME44aZ+DRVl1mGqMISyhihr13KedEcs72a1/Ezf0sA/DV
UN8ySf/1SxxA0tEIVmFCBNCijRWiWQUcKIe7ZhstaUi3vn4NQ86754bKE/QubJvuLfjRd63Uo65v
rHhMXo9wEPy07cB0/q1QRCOorYpPASwFr4ojwcqSrGf07/xh477pL5fzQQpb5uVDHmtr3eR0XZMA
QC4RMbmyVRYEZsQMRqaA9VDP7qubGR31KWmy7v82jBy/nHaQAToSJYnVwF9EXU9pg5lj6CIMAqn7
akF5OXsYOXrjDhHht3VGarjE9kOxBETuplWXrDStvmsbBGsAhRnKsoGJVCuo/gDxAvh6QsuSZuQL
Dz6qkJOSEDelctF/DiAWbmk22V6jERr+P5GGjQ5d4Rszvkah4Kn3BVVGnj8feI8/fIe/o40uMcyO
tCsI6PEnzYQggOZkSUmU/A/AXLNN+14+TUl+3ZSxTG4Pqp7V8JEM2kyHUzEnRkqKNoWrbK2gdBp7
9HdWAZfTEYTZ5g9gJS9J4pCrU1X1DmlCo8V+xylVZCjbhWwlZyScs+SjxLH55xuRGBsF75oevPwN
frZ/Tq7IyuBCATfv6HkcRM5znne6a9vHjkHYd6NXF1t3ZICMxIGeWe1jNiEEGDpu/35wKLDkKpGu
1Ntuun4Xu9YClr3lIOrUrDdPQNnK6o4hVwFrKq55D/tA299+EbVdhdf1r/Fcu4ASx8Q5B7fh71M+
q4A054V2+acXppgx34ukn1ozvT6c4k0Xlb0FGNbtilV/W8NMzsRelmnQX8ZgzSuVpwsW4cj3ViS0
nUzMyNFtb6+8AoDLGAyCyCeUNvJ81aZveyHsyWuE1UgK+sfKr7WeTfhGBHpNBxe/de1/nMHWxV+R
PqDCzLukdMm5f52DVg7FKPrBHMIH2AAE+UQ7dAmpVsQfX8NqKsT/6uJ94OnnEKkxGl1nIZbeCHxl
FqgZGicMZV/FltFryhI8GA5QyoJpUZZhFolgH1B7rQVHXIfUVUnnp8itzciIdni1hjY4giiWpSE4
SAgLrt00NCtTnJ1ooR29Sel+kYXLoBhiVwhjsYW0xsRFmeublfnt6miB0sIVgnn2nTURteljqUhK
GDb2K6maL6hsBa0RL7zXtrQbbZeRz1KZI3EYObg7L9khEzrd4lev69XIR7mKsC1ksom3pwF+NkAU
bBM/1n+HdDHIeljCfU7poaeh7qWFA0nOCbAZzAahb8C5gGlc25vQY+aR+3NiW2kXqxFbwaINvyOU
42ybmioxH5F//bL5n+zltoXjpYaZN1kDSfBW/nsQKo7THkJJAb1jGSP39qtk3i3jloGqCwiAFEdP
tsBqr/9GPGDU4e1hqJBPRAZP7reuEQWHR69TApcLUe0deUUF+lsSGtdVXIUlnoVGSFCKMoxopHvx
/9Va/anfOjLZ5NTyUYksGRyIQXh2Sx64E4yWHy4kqF4bil2lp3E7iu3c88A9XcLwq7BVfqtenPL+
7mHfrasW4FTXG5ahTR3Qmt4pagJm2LDf5tRqSMlgaTKItsmCKE1Jt+cmbt/iiv2pvyyP9yhUTGNW
S0Tr3AP/2ct6VBbmpa9RGoxR0K+arzSw+MWXHPm4JC4g3V/2IJOhRmeIlcADGz0ytfd7bVxA69iZ
ZDV7rrd8zQdUUpCkk/OBTj6ADdDHCTKkrIkZuD+Cn8Debto2K91krfZKQK+nEUAb4SEz/hxPGnUA
5YqWk0VeJMpPZ6JDYfW3aEtu/M0O7akw4xQED5psBfo2vA62Kzi193354QzJ0PATWxUpPY+cOqQI
0bsTMyUumtyNKDMMIZhWq306uas71LvtR/JcLIevUl40uu1oKVXWvessd3WAXS8PH7Dw47WEf/D0
vHJVp6jTOR5y4Wd9ycovhNBS9ueY07kUefeomXS3/wDwxvHOhnR5myqMiN31Y0/e+zBx1PLEdIO1
xC098lOxGV9Z5yxqj9+sTwMMy/KbZQehrToQ/SSjpu5J6yQunyi+MX3OgTZlnMLMUF65H6fbKEMg
tEHIa092UCvLDY46uqCmhDHvY91Fn2xCQxGRjuZtN+fhwk5suu3Hx5aal2ZCvFQstuR5UvH7aFEZ
nwmlNuVl+wqkgoqsas7RpCWjPUbYctQpZoACjA6xb3feQunt97psfWeYpolGDZah+YRMFFfBqy1a
s8bpI22QrCIifxiLgU2tIeuZVLri/oJx7hmnA6OCjm7t+HHpFjSyhkNUZdzIIMEOhEXLOi1zHa65
kpDqJ8p6RHiVbW2nNxz/omJ+r+FimV1YqiKJes4ZzNxA7FKrI8yIb6oWpn0hRIwciR1H0y9LArr9
ee4VdK2B9dU9pvExE79yVSl94RmEeTDTMjcBSGb5PccqNriE240DeU3m20jp/7U8YagxQmS0doET
p8m4lwEknIFOjzqPG1YSTxCrITffTF8OwUboPW5j8Y+RtS9maKho2SW3s/QC6qvfAEcOtgM4UZ7K
h1HZcPRtFg6gcQPGWm8v/nJD3HVSp+dXyoFV4NKjn/ujquyOijWkfkVkZ//EmELuBzD0ZKNd/jBH
vt260uIRB3v0ZvyfUbccNwsAAzqXhwH0WXRw2JKSQqGdWA5ZSHypQoI+kmFcaMFAUeqijz3e+ULj
wt2BxilancWfnt1BvkCXhX/UnNr85BleNypSa/d+g/i3WuvVC86j88ztgRnOMz2DTKvUTDJiyx4w
2qPMz1HuTjmPca0eelsq0ET93XYul8AomOJJ2NnYrM8z1MTWw2xMB0WTI0d8+McZyuXfPXlF+9Kq
L0QVkSCKSxT1VkMNkjbjck8RfJbATnvEDukXJEoZMT2up0925/hRMivxlyiARBNbRDLudfLPlMXR
+4KkRISAiPpSfyLVxDImG0N//EM+FG1jqPp5aGi/Do+7nKUaN+1IV/2izPZCr5N/qpWP4Yu4tATd
1S84p9exOzkgfYjZBbTZitNWOTA0tSINzyjAlGZgADmFYkma7LIxlF0OB+VtLUgDJQDxKaI173QH
i93k9jRYUSzDsaHYx/xfIJokfSr6iYsaPsXN7X6k7xmN8QJ5/prrsJVnTwbsR7Rx28EwCQhRYU24
r4P3oNIiFb/rn8sjyQWXgJK4jGd3guSSsWu5Hr6ALYjGL/BA5rflCrxYJFu0JUdZGTSZlVY/7f9j
WxuV3YtvdzmFiCd6DWK+pQ61bm3vgd5z9YqPRux6XkyTRD+P+W28YpUdqeMUw1IKr0mM2siz77h0
XRaGlaoA9oRxaLNzPjjvHmA913ykxxefEVbAYo78D/p71244QyJADwihOgO7C6CEWaJJzOgGdrVa
vtKyyCohfzFCqWVdg/o4TJW3j7lMGCNuzM7HqU+6/5RJl1Tm387euJWoL09dzeCpiicgNBcfGMnG
G6F24chsSHZwAeqvxdMECMHCQJ1lHPYyN8QdpU4OwGEyjfrpAirWXvUn+QL2+lFWgIae0eVtrkAx
N/h9NtZzWFI+OKMoYyVdlLP7gxbgYNh5SUI4JPjbrSMbtKvIOCSq0//TsZ25ealZnDyPpgxZsRtQ
jotpaTDWpwLum0PXrCZ9acL3e8/BdhiLsqZhCYGSMwFTWJ+2xqSC8LiRouju7LnanMKI86srk1o7
IMqsXNU/jM+Qud0WCHduaCXDjvYJA86iW8dHp+1vL8t0dgyKWTCykf0BCfks4Uzl4wLzohOBKB6C
SqCttIt6FfypR1JkF/V+7pm1BAHuMHDuGweOKfTQfa//z7Ij5pDypgku7VB8xLKMMi9f3gLrzt41
OPcPIsvMwtyvlQzAioTIh/6i0rv9pxR3ahdTw/FfGBKqjI3XpQcgBPeKPsyA4vvUsFKgSfM3C4/I
sSiwwY+STOfGxbCvwnKMiNT8b9qxo4joyWN20pW8GiR1DgybqqWwIdbfIytGS31xsTlcOPhxOMUo
+olzp8he2mhSkg15PILzscoQwn1fK7djB86UecsnbasqiXtF4AmWxInGiWkE71ugbXS5ei97ipnH
pe5xJNOfzh23RpawlGLVvRYZdRbixjUHbTUzn56VPBAem+SaqisbBSA8CX8UywyEoIitNuIOg1qQ
ipxz9zl0KEDjBgC6vCedwFafRkSs6d6nXLOOfUb+AteLBe2UkBT9MgAm2AFaCVR0AbB3FDwSP2Hn
3T74s4q/jAOrsbtxJoU38tfF7ejv01sFJp+QbBHi3SlsSIza3uNe4b+hAHxH6kGvh1b7MQ4B8ElY
cyzfmL40j3zb/N6CX9Iup7790ph4TGz/zRsqrgebCyHWNpXIdy8cBthb2GQz5GvLY2eX4cC2lrkH
ZgzIrIprrZL22lRtOs3nGIIUdyj+Ys0/GpXrzcdU0Be5OkO1jmU9aw/wIfFRE5DGIc6xg6pj0ReX
vKMRCXPuDPvcsFmMgmYAr5l8g2OkkjZc9+dkwk4+1bILb1kv8pQbLeInmpY+q2ygV+Oe0PA/lUH0
Nx9f2B7XTvheQ6ecuCf5HPg32zwX7h0WbroZLxl4pztZqeVaP7MdYJzhBp81jwpbZMm9VP3khTM2
WJclt5UC64vkyd21jpLCBEOR8fQtENgNo2oh4NyXMkTCMuvx4jK7U0v3GodMNbgVL6iKOLOWF9Xz
y/+eEQUggEgf7+XPeB3Qj25PHrYIL3z6df9BH/5jYa3j6x8PoaDxHfPstT6Pl1hIWMqfTDd5frFj
+9nUTP6vs2eZwlZFjW+b88o6eDRSv1locLMyegn8KD2td4N+D/W7Kp0JzUOtgdIVoCUN+/l0sDov
gfUE37RrzGzVAwKIZXdjZJX7ejn7l+3x7xjVjqeYKxt1mmFPSXTJNSJUOa92Bou8l+ZgQUZCDkdP
DQAh24eShBwddgxj+k8xam72k+Vl4xarz3iDUoEZFt3+0qRPgH15wDBUAn3e+ZlaEJo2n5E6zvp0
c4+VYY8q6rYgwuCxvf+6m3zifIeoNnSsdJJqRFBroo2TJv1N/y6+kbYUB6peqiIU6paz7ICNKAvH
blc1kG+3fDe4GtIUVnFzUBrSwIAx4Xi96FPcYiqOBDEG9fQEnLg0qC8RKtFhLK/L+iQftycB0+S7
4TJFDESHxtzfdnSAGwfG/GrSDeqNeGlwSNowI1X48h3uilKU2QR+Ec7sXs2VRbRCOGjQSCuyAWWC
y83UkZxoemzpxBq0IDUC4RcNGsrziMfFHy9CQ5eVJ3yGRDMFreGX550fhkV+3Hu73MHYmxqnidk/
rosH0DyQ5UlsCZ/pNWsJ9a+AqIYQfDdaKNn/FEgJdGAvcwWVXMnSjeuQcYaGgKIIF6AhOB9K8JqG
MJYNDhjmGcHAM+uhJb0WjHV44cOmDUpca2R0epBOm58xXINCIVrvAFGZ++hhQ/lW7DKsWPXqGEA0
zs5H0Tflq3ECNW0gw0HBu9Bfz2nbmolFBWKryIx4hiOpzFYh7OdUE8izA7huF6OzVaEBGRwbchbG
2M/GclHS92GeUXjA2zkltBU82CoU8i2e9vv8N3VfhO5rk/80yasSZg2UsgnxfPJzTQIwx6LJlg8O
mHR3mHDdGyurXTpku8kK9xthotglmAdSY+eyUGa578sErKf+Z7RJ5pkv5eleNCy2gMHl+1RGHHdh
AA4lUzemSuFMzhyAhK/dPMUlsmY/UX1U+CJOx2a5b4bC6T1b6GYKhCAKcmucKmkffCjbprGOqPk1
Py3PGM3sgLfFQyS+erF7wyxMeF4hkC0/Q/Wcnw/+L8VXsMzIJikwZ6HMj9CP/MPv2QLfgPxHwEzn
rN/GTF8fzYvRVIeTRhjaoPVhU8XdI9SYO4DFNi8IEQMsaFV5t9iD/Alhx1A/6X/jTeei6RHyswhY
rARqq7JJ5IbCvYhrHh6Su0icXAs6lBTbuXj8D9pp09P8xXGhFGH+agDU1CcSR014jAXUwWMNEUvG
Mc6KOmxgItYSzomHBuk9rU3YIyL4qeEbkMSeyhjOHtiTwwtWer09K/PC1qiKqQie6K+6HBngGJh6
egKEu932GI3BokWa3lm+lUcoZipsqb1tJTPvMJdA0A9PhXEh0U8jfmzNFtjZAIoCk3zmNPCKNlyX
RPcUFc0TjLUVu81G5UNqmZm9sl4dqTB0TOYm59Y1xiBMoGHUj/wO3Yb3gzBL8bk3XVtNGTtCOn0F
UG/MNZW7rGdYfM7pxo7LuazUF/+IEemVdcIUHce0NuFqXm60w3sCPKicpx8odjGgRt6qbdEduNvl
fq857/hDIFdPc6VnycQcsrPd9qb3gk14pLUkb6KV3oIp7jXwT66Wwgm0/QcQvuOXOR9eGm1FMASa
EcQhMxsmDp1P0/lZ76imEitpeLgPQhk5xihcyTgV//EXUOBg612KarOLQCWenmgFg9nxTCbtin9j
QoHO6Hr8GCDs8UYf678BLhbO3M4glR09UNFNORVUqHBkEICmAl9j0bSrRnQSKq+DixrjAUsINKns
yogDRI+87kcl22Qcm8SbSh2ycPK4wEboEOBDaG6oigonNuhxc9s8BDoENFvcqsVU9JaqRVPwg00E
9muiFxnuamDT6ukuwzwHzbSWm0VF+HlBmanPkh0NbNL9UfrH9qS0oxEOTKs58d5rJvKByLdjo1Yr
+5gUAtHfHuT++iNJ8d+WIUhAK2g225xiOAvXgX2uY+8QWpLpG8t/GCgRvDwArvg+j0OOYan2isZl
BC4Eg++f+x3+JgnXEGNnc8xT4ZgH6VAFPWBdriRGWU0P4uvXpJBrHiiOjcwl+cZyxXmDvLFHZUQD
l8ojmgBGz/EVu0YexhBV11Wr3sU18HdXLNj0pMSYJM+uZGVeskgs6K7DDZgAHC6AHy3ZcjFZPMLS
o+KdoBI8asWUlhbL6r8k5shXYDNu5B7yGobuqlLpbwrf4KdA7MoX5U8aM+coQPu/TGrmKmazHw1r
F/ed6RTyn6i1NsfOoA4Tdj5SMCVYUrhJxplV77AzimXjx7ag7yfXjaNewMM9mCxzPTefo9TXlu8g
l23uCDUiCtglm5HOKubPK29OGsb7WvscCsgI0K0uQBRM/O60mv3r/Wpy7Ni9AKdbPVYV/p1sr6Nv
VYpT7R7kxRJJLxTIAnVwLYynIEHiiQsSiFgbUZ4pgtO3ZW9O9esCFrzPGZdMMTjeGQZJ3q8+5n8u
A71F4g4Wcl2oIYegg91NWCwMDFQihbcL/CkqfADtvon00jGOjjWf6HdFEU4wnmlwKG/yGjqIP8P1
N25YyRLBqYTEgDnhcjrIZhQHE6uMiO0b2sLWCHGssTV5Z33YMBqAHI+9YoFbCm8JAZ6MpBsWTMsR
Eg+DVoePNXXXSKPpHKUA+Qv84olfcjhQ6t54g/4jC4OupNgnfv9Admt7u4IClRO+Bu8AWLMJfBPn
T2tBWMXucHimJpplKkAt5uUJ3/uWG+O/yeNWofbKsJ0gBFdmkzPcbETV9rwIR4b9v9d/71lCEUiO
myaiUUS4WUiEtl6QI1qM1w+aQd13tSb+Y+RV0DWmHuK2M22oj5mC2IcdOE791flLO92e/FPKqQ3k
wR5qg2IwQr0LSg2MIvoXOMoPQj1+LkD8C2hgCZlqvg72Ho5UJMfS9/F+vEpCOr0maAMRMcFHh/VL
tE8wi4vsl2s9MX+ixL39Bv95UEEVt6TKfjI8h9qcmEl0Ww4QILLOCveAXk472Fd1SwTgzCS+QUYM
VPydR2R5oqPrQXM9nxrLUUHrmLftHE8V288A1fPiIFRzRxRunmN7Nzu8aN3knXprBsyIzxh2Ba5v
tqd8yKSY4l546d1z6LfCs8thfv1iwKowq5rgU3d2DwppmC7Em2PB9wjoaL7B0ZX20PCDB9uMk6lO
X3xjt8guDesGf6C1YgT1fsavEOD1S7jSmYMpTEx+z75dPiYNkHmzS9Av3Tdc5wUWV/NmMVMrXOhE
CJ5dCgitdcvinF4Ch/z8OPO2gnpjad2PNlYoZTzKoUm49fyHSucAOaLCOKzTMX0ppeWw8uvPCgjk
aFo1koC6k6mVNNkEfdvioQxysjSMNgoiBjfawLHM81kkw5Ek5ydGRIPDmqZd8PLvIjw3ByODsDjg
+MzE3RPAgz4MHPBS/2EGy3/rBkAT56fNJgbApRDZVdraYu5adEsJQ3rnfAzxYhbud6Tu09X6by6K
aAz3DWga4QrrBYQ57e75be8bzUtuRwIJfotg74gd5gQkuUclHmkZg3PhGKY759zWpSyrATAZmvqN
zz19zUpR8AlKwBgY8342+vH90IkbBRA3iEThLX4jAGLwU3n0wT/xh3HOQyiX/85Tc4E4UZ6aZ1G0
TO+ROPGvrzU3BP0liPb769P5C54zE97pc/gJYLRt9LITYre53/aaRVoMC5o3EfcWAq1JhunHZkk1
U2u9zOUayUvD8gVy+BEYQmv4vkeaPyMEMBMxjSSMSPzMdi8RzNsu1ZWbrMbMhVLFmOY5dXfDSUFc
KVooGNtCYBN/8KBx2EuMWrwxOgZwaDu6nZ4pC/fwOAbe81AZTIKBd/eBPtrscPwgVZjepwY60MD1
rMd74EwJ7OZKdEvnlgRjUYIsBc2Ax8QffJiMOfYl7qLG63/8fwG5680zYqm22FYU4kkLkHXnbdPc
6VnQFw+F44UZ3coWN6QPGXQBafmbCBT6P+jbeiznvtHDny4IrYlpG8OACLrfQL7wYeEEG6jbujB0
TxOMMod971ujF/pbYF5kWgTW+TqUseoCcFwrky/rAJeFpdKGJfX5NLVFZN/Uqm/Pssby8MaAyJwm
+MtVKPmef2mRGeOJvTVfu+Aew/CH0bLM/jZc8ONqn1giE16yBREhUqirqI3fMIprhs1W9igqMH9b
Nc+SVkkmHUXu0NmvUQV8nRHNVHCCG60UcFYOslx6HeJWjD63lkeEUULXnmO1jkjMaM+neVcUENTy
HjNlW3ZLLMwQUg/RKqq9BW3uCEfUCtfKr4phHfiMNXxFHdxO5dfWVK7wwjymfAc4L2GBFpAoY62A
V42gdBdpuGYt1xFi13G3fcUd5FLe/GsgX7NmhvYtOvHC72lry8A97Ml0HxnFeoXXx+W6o8hghbrR
8X5vkytKaH3XHbxbC2SGTzrBjBMwfY3uSTwUMdgM6ymKb0XczxyWUN6xkS9Kveq8TmqqkE3uDHnF
w/P62nDY9PE8hcLBdV9D3U0i29mCoZNn8gHeEi8GEPLiKBM6JPSt2lhK5qAtDWbR4nZwxnUMEPIE
VAkj/JRjunbWv6uZcTB2Hu+cPHCrfLHRBcPGbjNxiIQ1/TRqStxMExuYtjqQum9ZOrdZA4ufe2+z
O7GwKsCOF2MnP4XXDrdVdhPRbK4XYj4a5/lua3dQzjOL2ZFNt2mYDCIKjOMz3fbUVz8eeUiMoe+v
OR3pYWXpT8w6x8S+vFacKfKWjkoxoH46atesv79ym2cASFoGFUIt4ux0RCvyPZKrezotCeL9z1q3
nmdZOapK0uAlyorP7TEq3OeV/d/01zo1dVnlnmx8SCaw5EEMxtzlNIfEnzb13UzR72Ri3/Iby5Nu
h79iQSSUhQXkUVwHp177E0VED/ur5sjMSngMTuBAfRnyIbPuAoFBmXvldv9UhIO3/UIJ5LaWGbJU
u/6/jV8oDW+ZhXJ0hwxFG36BF86f3CdMf1PX93VzrLIOYbDNMyrVogOYSZjQigWn7T2MGuz4AIHe
ROviH5rRyqh6bjsfmwwt4bLUK8kGCjmzDD/c8TAeL1jpNjn0lSV9rqMVr1E51f1y9jbNHYisUfAj
8nFrcd/3SHTe/KqIxgMnUD+ndznoitdSG+w0BlgTUYDhaE14svJPsMNI3nn4k1KAZwdILFxI9VRB
PERLIWevwtJS1Kup88f5NgE3KVNypU7nHAkZitlmpXdfRNWQ9F0FqOXzWCcQgoLkhJwQTgsHuzaa
NI49LjYIwH0+MuSLRQXwr59udDjUM69GwMZx5jewb8cWBSYdrk37ALOcpDXCkIyz1RzRO3RONGDE
CweHp/qurqtVO9EY7rTUp+y7/qCZsIF0ZND8kyz4SzFmfCzmjIg8vWD3GzsGqErXglAvF8n7CXme
ZFdblsBdOwF0hwSU9zKcM5N1ZXPSa7FSMvPeB+zuBdeETXoGWXWZAJCTQd3ykulvYZ7jmhF/X6zu
wHt2zYYWZy0wG/dzKOHGejXg+AgyhA7yUs7RuEKFzgCmQrP01bNzCkXwbHCVEU5J6mL79aQ21aLq
zYOsd4XF0Q3u34fv9KjIv4GzeWCMP/zn5PMOfHhXW2AsiGEK9PtAbFiQpFddF3wgY4vGpXahxH54
nDO2AVCpMwypploz6PoLKEM7KHWi7lF5yz5g5Jbyl1Il7dHkQejv0aWJRvmCtF38Qs0QkbU1oBVC
q4a9qBEjPxRa1Vx50irxbh/LDmRnWJolOWDPm8xSjGN6dFu+Sbrsh02s56NzW/ZBd5B7ETajHcCG
Va6CRjsOkzUVQ3ZCvzfNIYzyZFwaTIBO9VgqNH6xKpdXY47lnlYYpVyYTI9Ty13RNI1LkCGhwMOm
/pFEEsYktl3M5utovFFza36N3wiQzrQ+7nfv+WjJCBFuBbugpDhS14EerfZsmNVHmghbS859tp4i
sjONghmLeIbdJwpl0idQR0gg85sdrIz4pyDSrGWJ/W0zo0kZy/bONR6u9yxxMR6BJOY04981yC1j
N/hJPEZpRjwtL0D0ZP7LmxzHmgspWtcUdrkqoTZhr+Vszp4kYtBMECyMM7YH6FUm7/ZUDl3/dKhe
RKaesLLluv0NBI0dC3WVfrX0K2XqjCN14zTO2HUgd7mJkTSjgaXzlfBOJnNqbk7LgedKwKYBx7mv
OUUI23FwCgPq+HCy9UB8oDUPWPGlLHS6E5FbfLidLgZ2Jt4wtuWakZqW4whn8h1PVKV3gMaua/LE
DRs52F0yCHHLZq5jRHsPl6/0fEVztxXVpo+lLMLTRNVC7I48bn/hyj8l7hPuNhP/MVSOgmPCCFp9
jn+CxHPk4hKag1SS2RCYVigBbo/kR8dIP0PJBPu4qACNZRxFGY9hm6SXcxIm8isWCIuWE364hKXF
TFVN+u+laKDtXGDltTiUTEJCktTLl3L56oIxWjDAbz8b3IcnZRMzuzswWTlSKKzXXBwrFC+xXqxD
RM32BauDhYCpbXe3eJrXPWTfJH8rS46jOntSu5anwEWJqirVLZZBMzTJiqEdfTQgPfT5cqqe4JLL
JsVgNuj2EoCcMx8TqTDla56wifQiBbrUa0jFEG347rCtS/Y0PKrIhha56sENiVdxWWxyI/ewqfNT
Nf4hIjPqo4ic09hfLPDt3nKB1/d7O3Sy0c4UzvKC1fJsL1oRW7rVWbBFuqPxzGFzsueO0jj9DbX9
Zta/AqvMNSLWzBCOtVpKhOLgY9mSawBa+lmoxZrfKPNFCMsP1+SV4ertNLE4WdqiZEYwnpnZlcz6
T5XxOY3ZVDpBOQ1cAyIDZHX4RajfNZ2/tbdGE1Y7onuVpoZghExV44pTIDpuEw7OpTWBX4Su20Lg
OM16hYBG4R9rLY3LovcZP4N138vYGZ4Z8cLrUAE2jy6s0RtxIe37xY1YFnOyZ8/o3Nc36rU1SZpY
nWaJFmx1aVoHRjdDFy8kxbhY0/WX4nNM6TRovZdU3OEG+++gtRPHTvzmIK69dDTT8rWq9KCXdMll
rp/BGJHeXJz/E2++IGJxYpjhWVfjvdChZgxojRPg9ISm2N7M0EaeE/6polsNNv8c1pqjG7MoNcNb
LnUCIB7FStrKiuiBSP4nDxYsd7AECleOEN5RDID2cJgTEYBTJxCQXeAKqDeCzujpmxkMSVEs1Hl3
hAd+RA6CY9Iveu0TNf/V4eB1uxNpSKmwL9KuhcjL9rbCr6eNeLC9KJriUicS0jHn7Zdn3GSiHybm
mg+6WllPv4vDc2ruwlwe0M7jNi0hhWO9xnqEt8lOudwdb0K6vdkLDMAxMI4uOMzXaCnYsoKQK5We
9DePvjaJHXQKPwIOZtsWjSmM8Co4odtmchr+KPTkwKlaDqpdQRA86yTpTehJlprEg4r7GahP4HGj
CnclgesxYZacxmQ9SAYO9dHX/gmZqZFn+esL3vJF8AKUEBXqGlrUt99JjbzRVsPkHR8QSsrwxNgf
f+njT43uphrYD7ISs3fMLkYKLyoBqPuC9+/YD6LAyHGMRIlRPHu0/GSoTeQgCGhK186o0EyYt6oC
rUPObT0YzZOsFZVIq37fpnZJkW5VDDQdcD/aeWbLg4475o41+hhEoStJQxwNI/fJZf7eNTawPoL5
p3hQVaUyR1LH5rs5MSOFRwIYQuqGCZNF+7yZvPmlcRVFyHFJt5BIoGlg2oCJVRKYEwLtcz3b0GaW
EB14vewltBOckxs5ZilNzaVN2lqAVGvnhxNSpIEOv0Cs0/E+Zs57jALfbt3zZWajKKIemTI5un2A
DEexy1Ej5Ym/xXvdfGkYLX/bDUbRH5sMBj0yOVB+o+xist4x7k6r+3tXHi56aLnmq06Wn5BHyHox
XtZ6oQ2QoeIbl2nr7wIeVIdxBU7NRcAh/6K9OkfCTBaxmJeYk/vmG5YCYG9EjSADf3NO6/Yxz5rX
A5pgAJQJSC5PEvnO9vVKu7LA/m8f9h0vc0XlWKsSNp+WolzJCKjMzKsaXzqoeQ5dStOvIqHx6tAk
6wRJiPp9jICIxIr0/GpnceFNWWDwZWIEKTqP9TirEkq2BTRStP4ABaRmIrBO+r87Pqku+VHkeTbd
bLr1vLOo4ZVuagq3uQc5u4KGwK87GsQoVf3VfQkovJ2Rus9OIp81PwzK5W7cBayz7LGpQIekrqjG
hQzsCNmEaljlN6uyZPpNQejxVM7oXpgQFW09D/OqSkRFIKOatTVp3bnpBFBrL+a7YNbmCSmPDPnB
4ecdG6M5dXxnNXcvCdN2prIl8nxr6xtIyxazkdYt3lo7zAOTylFxOPn8LYlMJM6fO17cAbZ0YRGb
OQqaBasdGgKXShX4j9lzZg0Fq67BRaWAjAzPt65oO8+vzP6LtG+wwlpHCzxawOBB6EsDZYroX3lm
/s8eQ0qGfTL5wVAfKPwIwzvjBeEiEDNWlxjk3XTIjytVmb75XBWgE+BiCSy9aj8nWTX93m6gF9nP
BIS5L45zYYiNpvTAJJ4MydH8I5zO5HEsTE8ZyRy9vGD8xpJC6NOzAfiprqRBOfY8zzYdYghD/X9C
af9wgcaocqKP7lIHviKhdSl2TeJnIn8liFkfcBZ69/u6bpt3IB9pXxiXy/c8SmYspPfRU0UwiTr7
ZkqQOv+6QSzqNkFQJBFfMj/GaohdUvcM/UJ3PPVucjx4VIT3okk4DCYW+WTkLSFjuUTiTIRr3gHC
cSWQVcTMOxA8dhWyAveVd0oZ2jqizcmIrvZ9I5WVIsibGOrKsZxAZIWJqqv7d5AtQ9KNzjDg9sQo
kghn1/mqgmVL/iaamQpe5c/wRPHAyEfjY7FGjHrBDqa2JHRZkllrxtD8Xq/Yjgqui77Tfctv87yT
XI1d9UAZCGHXKtA56BfjMGD2LR7c2gxqLpZSYLhl2wmeSYOIvwPk9Akk6T8+vgv2AtvReg5LqfKA
z6ARL89dsgis66rC+UZzq4ff/aJ+J7mMkYBDSOPLgJGDLpJjP8x+TOn/+JFmZ/pSm69CppteWsXF
T4nZXEP92ZvKeOqqwEYy6/8CFlSGs9CS1RQAivvrSL3RRnHpLGoIMR2o4mILRRQp7J6ghrXh2WJt
9vvEeUOnhGFzfg7kDU4e8pa+dkwkZUo0GNhPtYYDprbmAXT0+K2saCCIEnzdTAvraFRtbJfD7cNE
cnGT1jq1P25jY0JOB4yqJ2Kszy6FiwS9dSGgow79q4jY1ga7Jr8CEMv4Ltp25F1jZPwtwPEhwdBb
cqYArYxQLkPLkiLLfn0mBDcs8CbGzm4og4IICJxhl+xy4bic8uHSu6aq+KuN88Ud7w4Y3PY01tlP
tJ7JYMm8ekVo6cLtXEd7MtHRInNToMVi4c64nEfhRN/fBsOw4i5WKV6IHEetdqzxpJimttUaLobD
quxRE6QzrdkMLnhWYVN+WLb3dGWhzNNPd3Z2GCqDFzHCIO34WoD1gUCLUhZR8gSWa+c3PiNlvlhx
hpM/53GKCMAIUG0NLK9TcnGGsiDkweN3t5pZ/NBD3+XB12yYnbj8qkt49zORRCgi4P9L6rfQJNVC
TGkeUvYROnUMyFoS2rDXXgtsehwh/hKX5fg522pGvPaxZ7ehz7qxAA0YF3emTyG1x42lB9PNGacJ
lw9FN7MX0XRR2V7GzI5AEi35bRx4o0XHO8GKNh+1Q+SaBBy14+4QIpP7ycPEF0ZLr3TYF2gg3M4C
XntDol15WFrPOHoWON2dsmrOKiBz0ZBIHeclUObENLuDjn1djNITnXeSYgOUEJ43KiWuGtC2CZyl
nCBhbNc48Q/16tV+dxWUtEHUrH9yIJfB+HfJ1RqTfDr8dUT+LWbftxIiA9/5lRvsKWxQKtTD0Cr/
gdhsvvoW8CiMS2x1gkzp2D/0RZKi80Fv5vPYxCcfdYQ8xRLpV1wivv9ZirVA1eYv7EyXxYQlJLNv
ggDWZju/GacHOD1Qw5ct+6B2UiqS0JQEzZfqtrxhBoGrZ4RChMcOAmSL2Xt6zwg9VMuiofFPLeAQ
VPKTks6Haf7gaQM/9MZuUTWwur3e0onEyECANMuS8c13eQuxkoSNUktlRJMg9z1VzDv5FM7Vaj0h
b5B6IKe2mMxFXW6rbtX2XQ1H0v7yO3IqfP44J7Q9zrA92FAzxKf6zMBfv/K4F/C5hM87Qye6sooi
Qc0OtZVieEA+qnFKRgDdvC6HpSn6EmRJdXqMixU4cVOvGlIbCoIeTym5jvgCrbM20mtScAuzR8Fh
o535Xrk/4cwgumxpJHPjb7jBLs/UPsOvQrtliggyp7iHZdL+4od33h3rdrmQQLqWlDGLc29KnWA8
pKsCGUfWi+ixF9hqGjWfpj/RCrRcMRnA8i11l2XZsqiOsvgP5CEPYYKeoDgZKRkDHK58pWiyhMvZ
71b9GeK75wa6REeIj6auqUH5hK5XruAszR4oPXXY98aFHXuEzph57SqFjd0M5nRsmYpcm60Vn7eM
2UeVkqbDMOO1AhkXKH11onS5uuKdVH44m9/WHZEXP9xXkKKMXmb1XySzWy4sobGVSw+/HSPvXD9j
Z4JyqN7pH9hpaVFQ3vemXofPyWCS2fMRs4mHkiFzoGBxbUl2zNzgiDZhXg5ILmiJ6iJ3amhWrVS5
L6da6vZiEaP8GiZ1S12VJy392HU7gCJiHTlddlDg0ikhnF9YcMq8MjzjZOjDyoQT/Op3nNJoi7BZ
mlzEV9Qna/PI+KaAveDBHMPFk2Z45zNqmCm5uFRc0ug3YUpemIAbAqAmmimrUmbXA0BB4NSrApPf
b0RdOLntRPD5P9qGWdxQFihGYSj1+y2pM2JV7V+JaM2BfeLGWh8ngzPmpDtqVLmBBAzygo6x4zuD
hHwiROHHpCmSf2hcbz5RNrpcHl2rs5UjmjpmXrNWNV60KzpbiQAEEgZpFwX79EXjB2Swi2NNQvkz
vjkF1XjVxoP4piPkySbhRGpShOMP3wheZMexFXdBUFMfWl/r44JhZDhVPIAiQxHWa56TPTI87l3J
TlGKMaEqfNSLRGK79WTJcWsL1IHILXfpsfWX0irPByJEjAXpuf4qpb6jPxWsxXGC0oxkzT4d6lIA
7OVnu+6e6ptXsGJqFeMDrkCzfJ64qxgMS3M/ytQpbQnPKPZ8c7CWPqmHBU+r7hq1Ylqisp+VigKZ
EKwL+UGLLJxOIoDs+9f8xnmMxfGMSVk5x0HigkvEa1rFu7fse00XDgyAJOhS+h8o98NKberyTNvq
LtaJ1LAMIdnvgVnTt+Wx/yNEWftxgzfVrxUvTDmDewu700JlJu00NgznV1Tj83oZSxSJ1w17keHI
UA8nQGvuHckzy9w236lwwDqz9CEBKlfrzJ63AgeruGcra6ivNA44jhz175uRBWUGH5sXrEyH3PNe
SO4zaefO43SmbFAzC3gOSevlOrxu7dFpOQh2VafLTpqUY3A4vVlBfT4xRE7KXIkKleqpuU4wyCuR
VFWR6hhTwE1ysgSa1rxu2gGbkUNPDN8pDvQxRQEoHr1UN4VNg07yY5sDgDbBcG3Nj/A4ZKs1du5R
VuaC0YR7UtSM8CcYQboyKQ2NUkSxIybWbshN7LCnv0m1pvGUr3mpv7X12g9QsN+Vw9pLeDJn2Goc
w6doR6CfI4a+mL7C55XAxyPNGoZHrNUkjRD5B2tOzHt0slNwvfr0Mykjpm/W+hDuUYLPvFf9Iej0
5wPWnZCpX9neiZxPYyp3LVmmZMZUd0DjPXRM2Pvyh2nKw2/KLZnmWX94MI3xA/+DOFgwIR1dKC6U
gmp+SzCLMK8D3adQXcV5qaAwDp6KtAbuYDfKIuMtMlquuJNsJ08W7Z9ARieD2KJG+7bNnlSXncNI
RqqyUWkN5gtdD9A3A5lcLKS0viA29bXJzMA92F28GHjSk/2Ln/Yob1HZBN+ysDRkAXM7L/uaKsiz
YXleS2dWBsY+sk7hfojrloWYln7rFYZJFfyhNRUcjGSzqXTEp81o5a+dkCI/Dg8cfaNJ2RJP+mpZ
p4BRdfN7TBYimBqWakXhfLXepP4m7vEyfNCuaWHucY3lTOk/2wEbzxzK1jqCLnURr4jffwDN4GWn
JwI/16pEFsLmeh0/dS8Jmsua5D/Pqlz1IGptbkzIid2/XafF8cqNBSEji4KJ6pm9vXQ7UBwXVKtx
I7d+9mUZ+TAwjJy6s2WL+BDM67CNF9vryZbT2kh1y9FlyLfHK3qTNP3hY8BfDcvO+gKJ0q97+fJV
VNH1XEwjkUh6S6qik1qYqAzmBn/0fl49VtgzYQFPxCBFptF+GmzN/PpOzTDrXdW3OT5cOxkEzgfH
8EQRN7XtD4NPoUmQONtrflltPUuiggeJ9LhE8XH0TLBoEXA3kJxbJPIux1wxZQ0sp2/ga/kpAdI+
1Q/3B/KopGach4tkPdgI0su898oChGdiAwAjlZB4DLKWvS+LhH8hX8QqKfAsJnYg33MbEwmK9eEL
ydhEIyc11ocOjbgqGQqjsoVm6z7s8KbTooVLTBZTkYGynUTMxGj7Nz8rQw6viUsLl2QtaShm26av
NpwK3AKxBgKeYy8SGO7Il665ey9kHylb8cskDSyBWgU3QYhTq+pnJQKFT/m46t/uWFx3y0Q82509
nR3QR5T9YBxVj/zpqak4X242zE+58izd8mvOTbyMOeL9/5M3hBBy3TQaQfigo4Hct9Aqb6kJKpgR
Mz9M+yunMxW1ofisiECg9eXieKlvUurzOYVXyj882qEu6/Prlo/DiEzOTTaEqcfGo1RyXnPCAUFQ
9b7pObviMOJ3/QxEw3no4e2B776RJsADD4WqukczkBCYTVbsWEOJ9vNSRgRiACRn2FIC2eBKrfqK
AaVS3qd8JRgEA2/xL/CWhpBPKmJiGqr/9axeFzuub3gglHj3uhnYoPMBFgW+WzfNqv3XiXGhuUuL
V89gG4bglXCxp+44OvzLOhehJxd2ebA9QGp8EX+mllNwQqmsfyfvv+E50Pj5HuiNPQV41rffBh0y
F6GQewerzcwRw3Kl4iy3T3YAzNSksz14yYzKYrUhsO2AXKkoRlzj1xMbUr/Y/CaRK5wmNWcJqNlC
uvNVXGSNILz+hnF/yqeceXJ/FHoJCmqtNbW0VolTbWtR10ePELlH0In0txkVl+Ojp7dbGpdUW8BR
jzHurlW49Ks2lqrw901Ir2hmQqN6MA8t28m9RREr4p0SiMN9tX1GSJoXBS3e9Pe9CtJr6wIIeV9m
7nU0aA/0X0w0ygu7humxOkj1iCQGLmZZ9IQnzx3mqJSaqhs4fa/xVwfXWqQCOsNs7YP1FDAF3uaY
0dC6yShHTBDu4DzXU+PQsL4r7x1tagIKsUuSM3OnyB5ZXRy4Gnn30lgBbpa6uRCftntAaoxw3boX
mJm28P8oS4mNBm7IxPSh6VeL/oLhio7u0nW4C6J6SHuELNwVY05towNCsOLdXml3WpaBJsMMv5lW
z9GGMoM+M1paayFZUFZxuG0hRQJWae8Q7YXpeXHIRFdt+22Wz1s1m9KMRXMzWuCcOAsQhqsXt8rj
u5QbaTctoJ2knAR47Yy1W+NbOSJbwpAIS21n0erikQVq6ml0GRkNzAlZgwn6TxEFOv/8n/v2zSEJ
eJhHETs3jz3h4x7DH0VT/Fl0oDV83bvQFt+sKEVPyoRRBGs3AAFI82JYrTpamRlv8sk4JeEYG2uB
6UIjUReIkzTVwqJJyXU2QVRQ7a6pNgCKGS65CWN9Rdn3wtHwVYAaiPjkzoWZprqiYnaLrAq6GOVV
kGl2tXiXysZf2RIrNqVpiCl23LZa19wYilDg7fIjdBoCi4w/Ks80x/KsqgR19YAWCnZ7kuyTaQMI
vc+FRZOQSzFxG3TEf4Kc4XRJOq0g8atnpT0Qo24mk2ZB3K7S5KBdNxC2kMQnNu820Y05uGYFvbx8
AzDP0Fwougf/1bjQjKstsenb6dklc3VcyY6KlSso68Lqu8dDmsd3Qx8z+7S5R/L0xeFAz+R3wUR9
uF48s8Aa1OLQ+j6u3qTV5jR1XikYs6ygysEUv2NO/BkniJQZ9oBE5pecJmLy3XPMqcqPtJbyYrpA
nf5QxaLpzGMwjM34CGPL9GIbdr2pPpUaP+kgQm1Xd4RlX86lbfAx0HrJI5fcCsHIl74lA+6R83tO
Opo3SSEzyEpBKhw55krjVOVXPatbmusEmGqCr/FxghB6SnPngGQiaFpo9Pq0KMMXqQO8rZSIJ7C7
K2wn5GG5snMiKetgPgh2MxKth64+ZTqkeb64PIQy3KrZAg27PkeToUCjWMQdJxdVV7DRL8tGU0jS
R45qGTFfHkLIkb+9OJcRnDfvRqctkGzXAE4tPBW+B7a9F+NyS7D6v+p0RIfaUcRsLBDIac0ILKoo
BlPrFNBFREexU2aZtBeJCV6viU/qdogTu7J0i8HoXUKUSN0hTRES7WGCUK0kyQ7V9P/myAkjD2C7
ZXZA7zZOwvE0a7u41+C3XUYs5+oNN1IpA1MrhEHhN8HQqygGVmRe6S1XZUjRl3aNcXg9v0BwCcXG
z3HM+mmoumGdyKI9OCjX0Ud4LXBClw0pHwOxxcV1vG+mp00H2JZyIE7VSUJyjz/etcHfozKEuksD
SGridCktsGFPmLqZ9Ndul4gnDbJWEAqu5/PbO5bca3rmorulm+m93gSQWF5jkzfm6E1od80E3DVH
Vb+dr4W0QS/A/RQBMAJGk2d0UB+emsojeQkEAzrG6EJ5O/5zwbE1E8Abx9l3vzzwO5IsUcuUhdVv
O0PQHvE/L1FXAU8QkwqXz5fWUS+F+uCYjFXvIBOlPIpDrZNMOTqK7maLT82A7Elcb8XLG7JqJwQe
0E8rrLt/0uDp12hGbf1ovrSDg7ZXaVJC2kiiZj0lG7No8L2aMh/BeVA2G1j1JAqZ4BdWlSZj0jtx
fPsByKr71Z/mjSxdg9hpjEwSu/69t6dsSKj7CSCLGFJUZKZujSXtxERKepgaliRz8APFVMa0r5Fb
YLWS+TiuIUCkdvFs451XKfseLHjY1osxRkwCgERuBQQCHzuKeJSQ+E++9AM2U6eXDvUru9KODMuo
yOvSZsiX0UIZ6z7GDYpeBXk3iDCeEkHFEnmzung7JhviYRaGbJDWP6U4RRfzk5tGEv+ClcKtfL37
6ghkcthE3SFQvnrzW7U52jMNommmzDJHLYRASzhitWgktsXv+hSBjLVYq1gnioSYbMYt8/P0Jsmi
W312MfXtQ9wiTv2RJ6joXulfr+EsmNwYuCoK5+7VZwvvylJqpsIpY7Lh9nDX2ZEzAyOyfrCVI284
GwaJMJlwPKdSteZfdDIYbA31xUF2XYUFnnkUsXF5p0AkCkkWn+1PLHk9re4qzIEb8Eh5KheH+VbH
DU9HbZwx5zNWJtNm+hV93x4K8ggOMr09ohYQ8snHaXWDuoBWXDnQ91EdRSLIyOKQDVy3X3K7u88E
8Vpu0B3MRCx+sxiVmWB4iC19ZFP8hnTH+nDCZcPItg7f2hDT1rO42YxHLCGwhj5xqI0iiMYXse5m
UKuslSgWiTh6/lI3iyw8XABXTmIFic6/io8t2eyOSAn1fq977KCMUc0U1SVWgetOJsmQZHWPaJQZ
0/CM4XtSX5SME0a1apOcEMylKSZh+Oiq+VKKk12xCcKfQSxRISISlpgXxGVmDs+2Wh97Jk+5BM/N
VnNcy6zW2BqUDgoB66h6lWTo25U4qeilFy2lpkHoCCT1tVh5uE4N84BQ3n/L7yNE3o3O6pwjh4E8
/xAl7bg+SBL+vgeQSUBnqYN0bU32Zum2qTiwMglEsbXNEaM2PlZNwyaZp0UxfKk10qmHyBrkk64U
ms1I+jrHBsvM4ownlcq0RLYWr47OJWA+Mq+aF3Wo2nxoQy74UsCMCQGFbKR242F5ZJBw5fbgHqpp
phtAYbWHBwnjqsB6xGcbfO9hCIloCpGFJaCIIcvP7jLpvRrNTr7h7w6WJXxlQKvhPU1v8fNccOpr
gIB6roBPwmu0NgSNIELpoNrgtWOg5Qqdb1KafrTtD/ruNZWzIla8XcuARXozlQaLrPfgWttjNt5t
20jH4Yrop8lomVQHIGlYbBAjOc4WSL96/QggGr/5zgVOXAVtVDpWYdWA90uf6vi3wDVmd9OVCwUk
irBY5fpgzGCyeKQuIJDNFcUup6d4kGyNp+nrWWqaFAVAin6gs8IXpLYti7hmpHwb3VWW5kUmEL3d
vS/wtzILnFjVS3MyoL8tZ+2wdVdgGOJ16XN/lu/W6RJhG2CmMRXHNBbmGknLtLAL1JLAUXGD2JRA
iqIoX6W4Oi3jhUycWIVP/fKzT51jkEyDKyIlMdjJEWwrSgXDwRLY910B+t2Mdua+UsA6xMmB0Lbl
sbHKtAqNdW/du4D4ABaW/nbVr4uHgnoEjtET4spHHMuJxhb9DHKOxOEJnf+vHz8fKf7ra6hh9Pca
llPnit+Ij5M8ZjaZ4iVUD3tmb9ljc4uN0o94ocBfqYGP4jSlLekPfZkjBqIMhzrHLQYmxYWauPIk
WGiixghaNNlwi2M/1KQYiCO2RdPHFHtKekIu/fe/DrNCZWjVfLJFkLl5o6NAoe/kkPdJcpi805jM
6BQIMfPYVTXFFm4HcOL06yLjHU+djjdiRz3o/1cp4wv7dPzPGivKkXJr8pNjpFqS3be3s34/8A+3
w5tOPY+JjOrRJx59mficmgF/EmQF3O7btwMbmMi71NCk3H3gX0YAn3VsNOgh3lWiDJOdY2L9HVj6
lPGr9YU8q5mS3tYBZRHrKkTG8AnV1VObjEESt6JDjRC0FCHWLVQqczuBweCM+z/AJ0NjL7488bph
CqIlvB3sSjHAO6EUdH1B93nv5WiUotxIulR5ejfl5IR5zA0Y3Divo3R3OLXTCB5qWUynH4SDuWCu
AA7XF8exYpSfhl80t1pMhEROgMxIoOmGWA7eUWiUD8PBEafbC8xwwAmriv8zunRC8Hva4kdznq/w
BE6D+hc59ZyTuJhqRpZAp/tMExylttS7n0ReJZUUYjFcuKswphW/ZtpgJzLwfrFfYyXjO8ph0l7K
5Jt68QFeuedhNpgPysFDg9D5BOg9sLDcp2t0pTXUzbbokG2SruXKeu4FiMpQek4LYliCckw8OBRE
cqGO8np2Wuj7aRklDBDCanKTMbK5vPDvkOz/Y8e+dhm6fTJSIeFag+ujND/yu7FR+LPJiMGOCYkS
t4NDXqgLwRszeagRZO3yrIuA6P7MH7LovW9ZkKmjfI1QtoIJBM5PnlDy6CIyDZ3sHTXd62MZHjbL
T9CCqi6WoIe7IGuGI2Q0nnrbWBYm20dJlRHmaHmJLgtvZkUDZi1levr3ehHiHZNuzOXRsro3D6Ga
5v7pC1Kr0hI7rN5iSwchejrmhDGZqkx4BpkiORD39wGrMjt8MDt4K4ApkqDWhy9voyo0+kMqTMZN
SDfd0c8RUXqrL0KUloMyZrNxTWVEdoyp6o0uu9B4gzZ5uHebNifL1C2AiAgNKRcUlyLO0RdQFP+t
8sMYrFx+5F05HXZnSXfnByoFjJtDdHAxFovU25j43gVMv7N/zGgqHXE5FfbS6YcScPTZFafVQUri
3HXTgsD7DHThUnzegeHGhvf0TQFDS06bdLx2AwoSBVh5XpnOF6iwmO3gFiRPdL6mYrQcQa0r7V1h
ViF0LFth/N4nWDa89mVyHJ9nUXTbDeIDPUu96JoUYQBGPBmLvSto+4k8pn0k8Yp2da/UO0x0t0WF
P7vjT1UCTRS1KT2ZT+jKOzbD4WN+7crLZHNJQuRUyKkVWxYiIhkc10XCRjFs3X7WmC01Y8fBwXbR
zGfC4vg8cI9eZfXeKjiy0HaUleZ3U5QlBtYmX2jaqqSDjU2hpzaXBBbipXNFyGdGXxR4NYBkNuhX
tAXrbGZMtjS3W+rWejn9L0RKWxOscUMI8KwAnANDzs6YnZPtZ8d83nqG8+vjj7McUxebJwUhbUJ+
uT0GKvHNPEREb3cBhMs6dzI/CX23+Zhys/FmbN/qFfl1RdQA+l23thfeyRtkLCy9ODYi+mgAUUJV
CBJVneKMUEPvlmv/MsNqKZaKxADn9LTEzWsIYnae6TiLrwureFjFjz7Z2d8wv2dHugiLk8ZUmvKs
/acv32GgCHCLZmGqH1HZgCX0RQsQprycRsIXd5lJvbbksiT9Gubnbspc/ia8P0mfl8RZwdX4SSx7
znpxv+zzra9XFx2W4Ol2JvOjmA1uZ9Xzb7XsSJOKOOS4IAAd0ZSAoO1wheavNppasf8Fhwi/3Pby
oKKeLzot43RxtYXoF5E4zJMdDpEhqsK5jvbEHNK1IGgsQE8Qew5kJy/DOiQfyekxN8dnsJgl79Ws
ekq/fe+R+SePA3W7nATHWDt0iLOAYUg4QNoBZNn9zYgDpNwZmw5DIdzdaVNSXODdoYp534gKbS69
ag2tAH0HQWXr5bCgUYfqCtxUMTjH9SWkQ6lBdXV6zjnVn0ZiOkXNxRJ+wiTIpe5SfDFNVSfatXQu
BZaZodZHw17Jl6XxKlSItyU3hPZvUEn+QF5nAoQvPxpuuWAT/Nou+UUaGH7PeUSpWWqS/A+4KSPa
eC9L4xMkBT9as65l4UfLxXAp/Tp7eYKmHBMOxVf/BFNgWEv6qwTk+YVtK6nhrIK3XutZchPjS7fs
YxuK1xNTPJYvUVZYD5M/H/kwMGoIPs+dlNNhS1EsL1nGhyD5Hvr2/ZbqIgX7DSHJ0QGEDX02yEPH
xkXqcWjYc4Tcz4nP0bBdih0gRoza8ROEBqeh43iyyX4RaQJ2VXyk6yhEADVD94Mssco/RJZ2L92+
MQzmn7rcbq4cbdm6rn/hfXWNf6ZviHR5jQD92n4/CbpCXyytbEFD47JfMPVdYBKTICrpltZSJ51c
REPzb17Xv64cckccBL8l4dfO8cS3KX6lYgPVNJjPQicLaC7lXo//rlM7m/j6MstzblMsr7254UfU
F1k+9I621MXaUVV1CmZsIEEx54MtxHOxlPUuc1Hre4WHLNviW+6NPwWa8oZs23rq+vrsG/NzNTM6
BQ9BqRD9yPxdEcKk7ouWh4kH4WkjSjke19nNicp7X+ocBj/vSz7Yqq6lOnGD3L/bKANb5euSjj6+
rWLKIUOoef/iktoUuhNrs/4lsCz5TUPAG78q1+QevzZ5GvvAckNoaUnTb5oJf2jFT+B45Qa1Xd1t
AwpiT///drv5KjLsQkm4bXandoqK9/u3eHKg17Zs3K8BPlwnrmoajxyLhNcnBnYq1qfAOX2uO2WS
ZM+h3c/76379t0Kh67jY9l8nicKpodo4+0tKuFpv50pEM+l6VxhUIRP9Vx6YR49HzAajJzBkWDWI
PvxczlJ0W+01WzJEG6HuS9Gr9HfP5jZjeecykoIXlOS/2dzSXDc1vQ3M0OOVzvG+iPgC9Numwv0o
rDdfMY4jJAZfD95CBD6HKXRY3YselGkUS6+1hgzomboVCxg1HZg/DlUWDCarNTbyt7QFkfCPusBR
KsN9ocRJSg2KPFQpA9zG/PLhlt+K5n96szdD/CHktFGKirYSXPQOfeFQNGic0IVBrfwaMGGxmnc+
05r/a20GwxlOrRsQH7JcCyDok2rpnxLoTdFZLUHn98zAJkgsUsF9/JlDy00eu2/sULrNAM/pkpAP
vUHHNREfkEdoTCxJt7boF1oOLhjHVZsN9AuHD9eajeY1w123B6leOGphyHVZktdzPTTYARqz095g
P0MjzUKNqeqwL1hWDig8iVG+1s2o6BxJGxWJVK4Aerc7QwR0DFX1ndrsJ6pJH9r0XtYKcYvWwUrV
ZukwmvPYvlJxu+e93vpbmT8qpVd2pL6DANH7jULFxZoC6baiBtpi9nCYbObeYlk6H6oq2BzWQJVI
17t54yo5Qu/arLsxz6JjhgBVEGtPZktqq2sdTKscNK1EEKSGIWrhh2E95g2Mic21GzTnZrr2MGru
Epm9hmWkKbJPgssRMJ7M6G9NV3LMeSSXP8RaL1MxXYgWbPNd1yotmPNWq6FW1Rzx0jRvt87qpy7K
amAAPUsGNWRaxVzlhHO74RVM3mFaCkhDJ8aWe8DyJ2V8IqlfhJ3zqRAs4EdQEc76VJAIwsJPNzLS
qpqdxuFIzIdNMAXjmxp/Ojl4Osr92W5gJHpafpMRuubyYkW1oAY9AdSGYp86Ey3GHWsJ5fDhNrlj
kb57XaonokyBdUv+mP0jtSpU2H4saSEwmH86eRvlFkNUoeTwnJnXTH7jc8wh9h2bVOjaycTczuBx
FP8PRpBI4oUN/z7GQAELCNrYnD4rNttkK8kZJwSpsLVQgwpilvzjOYBqn3JEUAwfyzqo7AOI40qB
QLEmubGMyd6M9c72OkUJstGqr+hUzzCj8aT3kyURzKx4DssnQpeW9qBagty1pfyXkeG3ibv69Kf5
8pl9TxeAiKmr6DK3yYIuTkVV49G+oGg/HLGKv3EZs3m2AzJRa97ZbBdfn68s+vAbXQ5i8ZKJFpoe
FaWq42MUAzqTJ9/eEXbQMaXPZNBmVYxA15x5FYPwCTm1WOVfYCVpoxW/SyDqD5ISNwaeW3J2AgW/
her+acQtnAYKA2cP1Dpku+R9Pl+Nu09Q2QmaHf2OKxqhRUy6syxUXyQo7B9Y0or8ZGdw1BnMMxv7
Qrqpa3+bfAsx5Erg73bUbfEVrlk4E3bAGqjxPWVlCHQXd5ZRv2ZFyVFM4QqePw/my09K1hTd4dME
tMuB6NYHTT9ZYQ8sJjPhWSZGmWOPAUawYKoij2y+B9frZ0Mi5DU7kOEgt7WWFxQfWQerv7Ypcm2F
CI88+XbAWOdCy7eCP7P53UxjMhs+c3p2FMQRbe7jpI5F+xwLGgpAsei3X1cLKdZtn7/eflg2EpSl
op5UISAWnNMaPtUsQQstVK/zCaHBUxjpMpmx+jVdV6kF1rh3MYLlI1TAuwPwtm6NOY0FTjcak4e7
1BlP0jjWc4Q5K5zil2Z939BYSyD7NtoehCXMZEYB+OgItKBAoszG0p7Dvph9klqo8ib6W52uMuVg
6dAV8wSGoIW5wBmfDYxxR5KTyDO+7rhITB1rWDWaJ6OsShetJZKLE7jwToTp8Zme09ftUTcI4ufQ
x0PlHaHVkbenm3nyZJuJrlzsk+iMYUq29F93f9CRIPnOvBACrVTG+A5wPLmW0UcvX0vkYqClkUYb
znGSLg8RxIJ9KM7CVz3OwD2zlmV+klo0iUvMWrpzY5H8olAL3pMWFWoKzUgocdA1K7h87i2N7WN6
3w2xrQ9JeWz64hWsYg3FweVv51L1h/2/kRbJtUysaSTRmGV9czDIuNiWcaMSLF0YFlzevMM8r9Tv
uvJmy3tiZr9ZPem6cwWbpgPhr1vL1I2Tj1YwU/rGe8dPfCadCO8muJgez0DjtSle6toplJoY9SOe
6NE8ASTT191NPga7V+OmWyflvIWBMGkMd5HQJ2X+FWRf9uBiWu4cOPGe9i50ZaL55UZA+lIDgwv8
kUDydHUxWUZhr7cZmmKoj8eKuJsk1cPYnPeMkHjERJGMUurC8KxS97PUuLK4bjQ0auFcnECuPbIP
6ekxrFTw0zX/vzA4ZKXzo6iEzGTcjNBuaYTh/x0gPC5ghh4KCKnf7CByDDV4xUS/XTbekV8oO5oj
iEYwei5ajKUtbhVgHJkEYJT/wvSHlvX4hOiDCTIaV59UGV7Ims8Sr8lR07p7X+6daXGozo+LjaB9
qspNz7nht3j2T16Su/U1oEQYbJ/hNp5IiXXdvRRLmZU1bJChgNfl/WtXEIVs/LmBavQDL02AolDo
mGIlTV6CXvlQikvCqWd4PZyDX3Xy3UtI3EI/iNR8jFBsmAm3xN3dmK3vzFeqa0+t5EH4V1RSW2uj
6ZgX0UtsjQAO839ifYprEiluYsEoIeBon1OjmtKTGgSsUFd0/q32rtV9pZvadOHkg+vP94wrey1O
X/LDctWcFu8sOmJVDshVzRjzodDvtk31akqzuBqyyCdXDNgF37zQVAOwYsFejxGdAHC2ZJY+XJvA
ywwkLFAz0uo28skysLA0tL7kkybFb6+jsENz8yQpD7VWmvmQdFnRMMseMehkaCo6FyUkeJ2gPvcm
JWMFgUfKwlBPXDCbNPU3wmQC54+P70k7rjKDZ7LqmzNKaNfyc/EMIJ/hbVQ9gMfjnHuXmUi1CmRj
7CZadbb1OuniXvkr5/cjIVfAlJPH/aG6TLkVQB1jDiY3QfDIL6lyzIA8yzVRTuIYmZnUXLk8XrXl
IfiasVPG0Q21nACxtgpXuCcQ05/vY/xWeqGz++I1341OztlUIP/LA5Tp/xHbp5ox0Q3UG0MYn+wn
YFE6KNC3UGJNY9+X9OZQRHU6jzRNXrIVrSjoHLEkXANGJ85XJ3eHOPX0VmfUWRTGnTNN28l8lvcY
gtV1bvJwfSQIwdb9+FvKyxCxTQGcW59SODDUCu3cbpIGOxj+c/j866LFrgXhKb3dKkmbYR0PlpZD
o8XMGQ2WR5RUS8KAWzY4dHqdz9mvs9nAqxnZEI4nIekKqnWoR/YS6xC+5e+MD6rkGKpISu+BStQR
A34gVnFe4A1CEZEF/3XuCWAegS7Sh6w+f3ERqbnnRkPNW3QwhsZgIVttU5U4VguwEv3usI8f3P8V
CIhY13xpfifvl0uRaUVati0tnrmh7Ecdr7EoXAwkOGqOcGCUl1m3SeCr1taezv219CMfI26kyoGt
/ULLcWKyHLzQVdOed7aA4D8P1J7LflUzmb4nIiqhoJhjSO0shZyOgThbQ+PTsaYNam3h+UTFniFF
fHSMDwHvhB0/8Gxufkb9igaDCe7cCqiwaop0cVpXNG4DycFqSn9kLI/3ZBCIIQa3fcKVBRlPvrcp
dUI/IvUsLMSABvwlB8zgz6OB5WOVhiySvpMxKEInNPY5j21meh4ZH7d4FwlxdxUGCZXqtb1n9dgh
I/lxcRKhmcWEh93ayGG6Y4Z7iYgZAaAx9SWiuxyMO6luTptasiMhC41qgM6jyEtqfedxpXZnJGNp
ti5UPShSc8n9lzcRiOH6M9uMZ7LOgPw4D+xXi0vWTcTcnBsIzpZ388JYOcCYT1qVWWxieDRXjWtH
0a98dsZ3G23n0LDIv5fQZaXTWGyXxeYHAAkdyxWOUi/cELQwZGqwITqMsNF7qJICNF1c+dqT+S4t
EVw2q4j0MqaIjstehsGL4aqrBJYx5ck0z4p+JIoCUKQhZ8cgj2dl0rzw4g/vAZPhN1GimhriJdRP
aaI7qPSLzEd/LoNrGDDkMJzYyqefEsn04NCz+OKVGQYDGT9v11ab8P4MhilyaSW0VXXDX01YiebT
U33Y7wdwkQ65EKBMui7IUUk7jBLWxAZI4QtPKvCVfF1l7D1dImP0nO5zbeqOri71DCj+Aq3hRYLR
pLUCxdwK5fRQeNNV3ALU9cvU518vCNWBqPb6ufAxkHyTohx0Y79vhT3ntDDGrD8ZkS/UWFc6d3e2
RuOwyaWGlwwGL8+/iafZtojBRvN7JZgq7Fnwt9gxY/NggUdkQ1//HNoHYXzsSI4Eu+ACfTkp6rpH
HtCmV6rDA0Xx9/2TZeqS3Yfq+mxK2XEv7inX/TDik1+ht2GdSIkexdE1fhXqWGv3gn4mYt2QNaAK
B9Ju9b2t0/v0KV9PJ5CvYGTvHBphb4XNJ+UEW3NSBaqw4yoMU1Neqi3VgFhDHXNSmR+nRTIHZ/3p
QAfFQwKYcPuwEYsbJthQPsqEEpDxJgcNglUn20szsxQuLzvfB/XpVT33QfYKAtwWpCj1kPYrcOuI
aCB/pnJ9k1HTrpXcd6wp1KuCNWbpp8YVeVxmLs4w28XqjALfnjZRM8xSdUM+1lu4cBRU0dt9GIiI
/5WbUNKLHxrPv51hPsMogrrTSUB89Uk9gyzKl2cxSTirJtEr1YGbsda+l1aFpzAwLewFHiWA4JKl
ekRsKyYPVzIaX5XS2kt5KSlAjaTDSeges7J9Sc2vfqfu1LeF+wW2YBUHTC0zvaMxakmGsLbHkSeN
1eD306a8g8prmDkTp/xylLmKs9auot6UKUHDANeNl/x5MSznBtSuMLUGam1D5mysler9Fi219FPP
1RHUL888vI6mTUWDZ0BoSkwsAUpLVGQIMTg5zloyd0GwFcu6VWZQ4mt6OoGXgWW/zEuSBdRfDGXB
cbzB1vZpi7u7VlxIUcLIepAT9ZhUj7roa8VjkAtnmAu95rly7kH6YklPhcnSfYg50SnvgD3N2ygU
533EiQYbIXdbiL6uSfjeQF0wBhr01ndsFt8DaxZkBlMSVqXwlAu3LAHc+84uanZ/unLddBtOS/+z
STe0UyBWCF3kTIgkWR+1ZoehpdcoVPq3e+Jb6DtTCcUdWpEYB0Z55sA6Vz4AVpg3PW4ZjinMwX9B
Rx79KA+EcICArZ1pJsnTZRct2TFjF0M0wVIF1t+X1y9CqIbkQmhFy3gkkC1TXVYnWxN+Ktzi3NTm
GUZ2ittPDajgCVtYxN1hHbMUQRuaP8T4Ghr4CCuC4CT6sCjQCdRFHjJyeci6DzFbAsXXI9utfpxz
hJ0hMncrX1u70Fdz4JeuuYZ//4fIJq/CdZRUCn6iE+G7vqiTgEvDR9BQYvi3RKiGGiSQ7NgUnt5M
nWPw1YOv5xF/b0H3lFEqn5qAGvZfgK0XrFGfDYFT1RBNwRdYHg4F3j01oRkPPpyxwIexcVywweM4
CIcSuGFDGYCruhTa0bDiGKtUywb/EN89wdjsmRWJQ6Qx4qJkWjSkNr+gy6USp/k8iUgXAzCfThXW
Xd2MAYagJHl/aCqxkTON8JOJcmxp1a4lqXhi19kC0m4RD9betXvmWrqilOEXO0GAWXI6NOLPov+c
fuEVJ7XXKUAWOh1FX7ERm/w+AartJdJ9q4Pnun+WFTTtDGiaymofFC0RhWlwIQJTcTPIbSKeVV7u
jQZ7mcGBtmpamAod4mSnXjkNev6Jbsjr4nl0EOTWs+NDL+5TwRYV68pCZpi2htWvtKAg61K5D/sw
ABLtRMQ1/ZbA6OuGJeWmxJx1L7La7uPYp8WTyxpE6215r/qZt6gVfA99xUJwv6CV+R+CSwsFAdtX
YGRMKGpP/6JlMLJ6hs3EszqWPbG5Dx3uOvUKtGVokym9NNdQvSAEmcV6CB9tAPE/IgYC6iwZFC8c
m6kuHBZoU6GQ/Tv1dEI/Qb0VbwjJYuFcwxq79JOtee9/bTxfnYuOdx1F68WVUWlHZv2IIQC0GGBZ
5TLexiLJG6wqDbdyXbymUC0o0ny4xa5WaDi8iB8jD86YmV9NWmOwDmCPEaOrIj5N2Je8Qg6A4fNU
EJoSmzpi8YO6Y9Q5zLJ2R/hztuyM003HIH3c9jJbfNOB5lnivkdFe8u6HWA2MpAU3A5btXECtOPa
X2lNgfeP8Y5zh2yY1p+bnueMXExo1WYhCMv7XqGwnIJ0cI8r/dZDmsRvabPTrQvbIemmqhAfYCR8
KTLyZzthOHPMoqmhM5b8vO9LTc1WWQp9zUqIzdk/LXAOSUN1x39+lnn2wM4Q+3TD68AO1rYEuO6R
YDeB9GD8IHnIUxO4pvOYHhzr6gHSx23DCfOd2lmxV9f6yrewc8abSLwed6ziz8N2pKDtE1CbCJv4
QLUKYUG4qqaRVfoR3bWypvWqZqFJq8GRx25b7tzxuTZd7PfRBedL5g5VOOHg+R8z41mIllxdBVmO
P2IYkAGFr4jd2iwTmb8cHCOOWzO0bEGYQ0nUYSF5I1vIvNaU4S+JuXqkmhAtWZnmVDR5QhbWLfI7
QVl6OaEpyqSgI6CMS0iVZTQWkBxsLi6QHn6FZOq+tskhCnzbtdnikgYVB8v7HrvQ1P+lMJceYdmO
Xg47Y7m1WomZt4FAk9JMSkUJXkdgmhmN8o4xogR918iI4AgbKOUVV90dMr7MB4NwsS/03zPZpGqo
awpOZ5cycQ4PiseMP/L6yVUNGmeQSyZAcnaEqsXQhSb0BcybjmmdEEU9Xu/fL2xqshvFytjtSszA
rvPDKY3GbA2L3WMzQrKBb9d2r6u+/QTOUUBPNM+0t+lzYaOjKyHW61rSVBanLcsmJHFQLt4+RcFt
oII5qpOOuU7anFMHny9Az9QW8d4GlkPiltS7DRw2KB9ZWJme0zH7V6mE+OQFr8snnFtJUiUfljOj
6fnAH+h5AezsCTJckyCPQpoW+5RXsg8kNBUWCEyvkkAQaigLPNDjPIHtxGCBs4YVfzDiem92K3A9
NdWTjf+mXMJkvr1s4EMcH6f6EoFrkfwyfp2lUv7WwHm8pCEJVPO8u6fttBWl/7zf5mw+JmjoFIIq
77U7Yr3ClAoYEvWH6RJ9E/k1nEo5nfKvQSMB/XnDuGW9Z0qRNeqlb1YgKIdDgmS6MrswmFQblmcc
oqx7ABqFtoxugLHFspwmz7ypbF0qn82R8Dl6c4D44tYR7oadc0p5nP+ei/cFU7qQCmp2+p8gc4ak
8mFaO2xtS9qjoPKkoc4acTg8iuvjEVOtYC7OaimpOurt/pzyk6Hifk6y5XMagUKZsLpdoHNmx1pb
6qkx4X7ZCVPkalvWsg1TOLM38fV8BcntUzqQuRTCbCDW0CCV6zCLwaLuKf+ZyF04eV5l6uF+2fU2
MBsgdGrpUVONFQs5E+16vUtL8ZVET6RVeaM14kOO2EJDV6frDiylPvrdoVL/fvP1l1NsxomGvUsA
AobqxczkcPx9K/MSHzYs+/dIzXebdks0n7VZlQEBy9ARmW4v//45oz+F5p0NLB1tMQmkcdywX/sP
Z/8UvO4TLoR+eQggoBU7xG+eqq2SrSQDeCeeT8v14TFDkYqK7W63+JiZqfVDz2ePVh1Ie9/jtUCb
HtFWqz3nVYZqQw8T0Y82bOxjr+hJw7nWg45fEkMY+5YIXKa9BifBWmMFdG8eTi0Np+VFNdVDKVaj
pbXYHxAwaElh5P59hm5ep3WRN0FL8qZvmqNa1KMNtJXGbeotf2q2GczAN7amvBLXpbarIgRUxpMG
iev1C0+vsCMsHHnM9GwY+N+mp2N9V8Ta0ZjofkXEAanmy/hjcSWSbijzCVcM4jWmzMp+pWNYtepj
WxICqtBIlNiYLLQbPrPkiT4x79cXVX9bzRSJ/NAEKnMwdOQmR3l0rJJ00UWDuR9nCgYhYhgKbFx8
HvpqvzgCO3NUhGL8VhQ130QK1D5xdHahAUG6pd+urzOvF7L1ZJMLwDmG9+18AkBy0HzOauP6fqo8
7snbgCMZgFgoYFU7pSOUSTxi8QSwNBg15AAMoZafwKy8+x2YCrrXpSJLvjn0ZCPQYfSKx4aV+zYB
OcPwBy605Y0ykl51Wmja4OnYGPRaMsVFBWjnoSR++r/q4J/bkwCKWtD99Qu3jqS5r/3/gbDZLkPk
jMyAl+xgeSXyhpkPeben7Zs/cY9tuThEZ07l5cKbj3KjjxkW2ObueNkkSXmVqQVxZ3ORxIK+AQ8w
I+ZVvLfq63gVY0j3ZULNbLRQ6q/dq6PG2bXis9Nxpa1SxFh9Cni7YY7sPrn24XlSICrjIJIQt2X2
8h1BMkmFOomWtCiTDh/5URZKYThaZrNMfDt4py2d3wMWjodU8/WrMsI4/mXoaSJZT2bXqPZUntdi
iDIAGn7rTxeYXWTP9fXYUSx2K53Cxz1pJNDY1eP2lKBo7120l8xOlcIr+l8IAJ0UgPUp9Id8NgYc
qcwxQet/C5tR1jKfl1abc/Ad3GwHnXGQZQofbzdTuygAA19wZUhcA+p6e5Y9y/+Rt/4vQATrzLlJ
tVyXCkvL333xLabwo4A1xKGurIHHBlodswG2oSQqSM+0NczC5h2kk3WgS2PTL9QwxX7eMwuXnPgn
EstO0taj+CDyD0S3mdVAJ3DnVopHauZb3OB6+Ywc8z2Aj4a8om1OqAO6+8HUsIGdO2to3Gk58BFi
Nh7PTcw4wV+G1CzNXU6kaMQSaIy37AsNYfMPxUH4nS84MK81LdeMtSDcU2S/vKjMzNsCRAEuAruz
BTYz6dJbXW7o9emF3iBIdh6EuqOKq8s/1FykFmDYstUmcFjS5fL/Z/GMDYBC+Pg9vq2LshJTfpse
0HzA7Bu95SJrAxSsfzy/G/mykyMYRksIF/DaaKuOn/JaUqUydyUENqo92QQaTrqa4nfIe4i3BiyY
0QEXhzuzZwRytl1ORTuuuKO0jBRhydLOnXQ9LxTB+G8DQif9Sb8pg+Ky7FKDT0/0M7vga6ji5czT
pidirEZnuRNkMG6PC2y4el+wNZ13cH7yK1ixvPOBvW5tnPFGqi5QoX3/6dUkCHBW4SRZUTQp+nmD
Wb+qanLM6w1IcjrFRbpenPdByKoxQVD7dcwjidNm3XkPt00F/0ObPyq2UXsPuMzx1QbmMIrqdISu
fR2nmgaq7sa+A8Ji1gJAWCCaK4h5IZqJTos5KRA9HSuy1tZhxkbZlohL/yegOQK+IaVECBdVRLBm
lPUfUVffWWJ2t0kNmOoDlUAbmhj/3O3uR8yLD+dpIVVb7voN+GTm+5LZqpMPhxHBvaPbahhntDhS
W6LlFeTN4N5dUwyDWMmj9guQnO1ZxUenau29z7nmmNW8/lY2kU03Y13Kz+GyttMCYLinxRfttz71
UxFP3dvFNgj3NTltJjFQNgcido8oDoweb7mIZT+G8qZTRIzrIqF2wDlyvcoTk5PBEbmp3a93gIDt
JR9BFMnQvyUspFWjUyEeEvXAwAbDn0/3/nJzodlIWW2B2td3uNhnmomIO/DTpognVgkv8KLqdV3E
5a/U3fxgYTLMAoVfm2NVsfoMRhW24FhF1XydjKdiEzAwDonu7idotTaKze44dW2Vc/2aYbzFIpsZ
r4KPJTvZiwMlXozgBOzVFVu8ayBaEzTRP/SSu8mmzpMm5fQ4RKKVqjIWbkytxj+Npw2SzRjZmOee
/p/J+vVMq6INiceJ5HIela5lm9oo/QqDuK1F5+OKcK4d0WjbdaORbphHSSjgXUEVpW7coAz1bl0W
AtRvRI7rUg/sn9PwWsZjdsTeGpcn9dsPdklYq+n+j/vFZz/relEeiCcPlr35RuSVHyI7fGizp6xx
NItuI3SX8Mc6aBV9GIbDh4frDyY0ribIq7qlUw1yrzfqYS6hwEuZGsQfb5Vgaartd+Z3qOO9lc8B
Evk+G04Z6Txb2Rt9gAm4Lcnw6FCUOZGPT5odQsY/RDucVKQsMywAytS5md3XAEmSbivCfEbcmkwS
BYEOwOu2s0MOctlBME9Y0JfIcIYfNficp/l6LIb8ogBfjkqYnI2kWD7S7CCzB17OtykliGqpVsxG
pYEolQFI09t2wcLFINq60VKBbed6ngEN4h2duZIwOPItWb69wKGGDV8ElPW4gzhutN5vQfh3VUSe
wLYdgoTzLQnLgmVfQEsUwldPbR6aaa27fCYE2Vump+ETGjG6mLe+M5qLMiBOWc54myb6GymvADlr
yQLzTg9WQqDCKtzWA6isLO//m943w5XKIgtSm/5jrGCpuKWqZ09nwxy7d/iHWxKavoUyLKQn7vX3
PERq+Op+XrDx9FEk1e3RoIfWN+9Kqg+GjJ75Jo5KkAZUkLpSsaYL01jaLVLeLOU5KQOHyDs+q5eE
XcDHMBjyiS+dnGyqI8qA7dtGvsoa6Y27X6fh6y411uRKRImeJoBz7UW2jCVU3Ji5C3DRcj1xGimI
DfYv35fntssO3udLaz4LvzDmCj9uD9+hyc/jkznPVfdDNAxzkZmcHwyzG9J2lhcT3MUuI2QtUQv0
73PjDAQojr5nII5XKOcANRw9zmabmWhXhtdPZ6tJaoby88elqgZh1C5n2s4iU32St+Djj7/WSV+i
3WcxsnKbl7OOwDGEIArTR/03J3WtL5/KptPB14H8P2+/L7Vels5tOSZ6mO6mE5sdm/U596vEYX7+
l/qshVp66qdTLqHvjV9OTVanIz4OgxNSt/hfER5c7e3uYpYHLRhhGB3HC1m6/JtQJhKqx68db+u3
p4CpvbXJAdZbGWURjD9FxpjZMCUvLG+vAxpBTzwhcMuM3swwutiwd9AcJRicFGaBndvG9zmERS/G
zXAXHNUISBvx2GsaVZlZECIyv9dnff5IfT/mpJschJ3PS53RXzx7iRn7l3OctcDvTm32kSEk+Gxt
VzdaUz5qBMMPdByazA0fgmlfK6Bq/xgkLayuW3KRG513QOBZ6L/cUVC3Sl8XXbKhvK6wSKhI8pTU
TmHlYIdJkZ8E7IrYC6VSSV09gAMM7A0eIHLHBfIdNiKRvAa8J43Ym9wJ3ee9GRwEZUVvg+d9Kr5v
7eIXhPJsxPC0/qRGjKQMtwaMws2CIlVE+JlTFH3iWWvduv1t+sb7joJWynWoCusB0fjZyaf2uKau
ASIfQ5aqr7M8vNpCjJJh7BCQtcgO8YTT5sEsAEKGbBC1pFPZl9IKyxJAPmYsKk1EcUCB5tK9zJCk
ThuueVdyW4fn5EIDi6ykPi5kiITI86I64/K+CuQnkVZ/tcgRd0Yb6IT0bCszPEBY2q+NEzHc4aVn
29RVeXpJRhlREaxqvGSSOK2RT2/SzjRg7ZSH+qWWXcDZK7Y1EFcRSV69QwGjxhScWD/2skdL4eP/
kcFaPfNjTD03yv3CchvsXSSwUeTnrYxrH58zXnKz3ee5NRxCIVHjvqCX8vF89DqZ8kGGZpfv1EAN
R6I/loGIEu7tpyNXmNA42J8mRDEPdIs4MQIOUrHS+u4dQdGU4sAIswOlFUwFdyeWoK+cDnXA2ctz
Kf53w4vobhh9Dl2X3y3/uSCd4gmFtGatGi3u9VCcclZwt53cPcCogT/wweNBpaxuGPyaXomgkDXo
vOGhkJAcKsYTQVRoFXp/1WsTV1LqiyJXPyYZC+nAaNo34XQd9rfd5Udmn8g8Not0Mv/LNlCwwqSP
2kUqH3IMLlkUfAfzUlkxMQQbd7D7IyPMqCZcvR4YV9tglxDuo/EYBJgnsgp4P9YzOdi+8i0WQ/XP
7QKlQI71j/DMOcaUdqdWWfkm0kOHNmF+xnBmhUaTPYPeBBHWBLLlXeZHO9aRtz9WCS0fW0WGEc7x
4piT43idsBXuJVliKjpxnA2T++Q8wqVas618/SfyHTLqaOSR8NZ0LTIwLH47cdtSQ7QM3XrYQZhP
bzAbng4NhDvc8hki28E3PM/f+vzru4K/DkgX6ZIf70lrO5nMwRclwwvZvm6XYwgIHDXYwjeyp1Fv
yOYg3VnRB1bEtSIHT93MvSsBmbUIH5lcjeTfkeHOdbL7VVhy3fJ7aw9eOD3alK9duukzXIBJmgfq
iGl8McJ35zVp8ik0sECz8Sx8d3BO9CS+lZHnBZ/YNTm5/K6p/jsKoWBL+QYfn7I04+0bK1zKfvHx
e+GdbKwAD3BUdUz4wURSoczGVDOHvZuDrDgWPlZ0NYtVHfSgJ7BRBop3gNBJt86qdw03P7qkUNMA
ilw31gce0fCNGKb0g4CuuWjFFkuA/i7Fqkwsb3VKaUDp6zGPBqPTdn19XwOw/sb0tC0lU704P5Y8
UXjt7tQ069/5xUEFc1UiGycAG1Z3y3nHfs9/5/FNjfmWK/3hp2mDpFX/tDC2ebzQVOShf+1vGv/5
ER9uThI+JA5NiPDRu1Mwm3NJD0HGE2S7n9Q/2xbB3mkLcDPVwLtIlgfvI0B2+VjBo0zcYG8trii/
x5iR7lPvt7ABjOtqnxrHk+SNp+bJIDgNaej8PpQtkJHqaYtCTVHoILc31MiT64xISVIbiI6MkzcR
qtMKap+Bi5mf2cNSznrDxZGyqI/arBoeq94d/aLd5khNf9tfVzxUngsQoFC4LcPIHIBP48PEEI9b
+v4DaAmsQ9+Br9eeX3dA4h/VOnKHvfwiNid8B5H62e+JWX7UnmOGV1me3p8+RR7uxEveyTMrb2uo
FDMXoiSVQf0U3z8RpRTqjXlue2EWF5D5EiRSIAf5UIMr+j7j2ft88t9WD/CafX73I3yhzZTAk+xC
fW4Wf7N0VscYOj4eSiUAt9YB/orEnoIbCrppyJPgKqaqqIQWTJHayFdV/8x/GUmbsMlT0DL5nXEU
A7+gdhln20i9b9pW8k1EslyOPQ1PSNLFnKV5yD5fHUDvyqA+qOZk6wWbBrAMqckp1azHSZNkXcnx
RVvpi/6YJDZ4bDKFtl+Tn9E2eozEh+7CfGWt4T7rSwOlZRxq85TlEZE+g8j0eIjLLTT2c98cHZPq
nIx52P7imyQIVpW3KuPBdtIx4jvODJADnZHtF+LKvtIsA2s34ZArwwNacSaQHAD/MLTWK1ukRb5z
0TUBvWouIe/w4fmaTUKwLDbYNPvJxZvp1TbfffnvDzBhZVBxIcgY3M9d/3PG4O4JZ4ue5kO6/yii
vSKGrA02WciNnGOLm4l7vCQ0dmelVB8zkBzktZYGGL5yex8vrYZsXsFL1bk6NkTzsLx0HUS0MqPx
mjVm3GCapfQj4YilhTCI03J6XHqWYj6HRpX6z58mIiNwAKEjw41i0KoppibiER6cfQShVvJNWXvP
Udz77eLiUE8L+Mr6mvRRUENnU3FgINNOmt1X5vBMWfMI0aWZ0Mdh3sl1PVbTrgEkBB72DGFfixxf
4niZC9PtzFPnozdak9oc8dFQf1pVOLo4e7LJ9Yyua4V81l7jkbIMpk06/aEe6Zjto6famLfoiuBO
MrQgZw1GUemTv5c6pJ60skm6LTyqga7XzevXfkOXYo6jrd8EHYZOZ7b7Ve7U/abOdjnHC7i8cvS6
cs+5PPJbb74GOuu+jn+1OBi6RSdjP/1p8eFp4sHzeNDXxs+pQSuojCQUIBSfBPpdJMsaWReHw8fH
iVk5cvk7AaCvfgxal8mnolX95Ya+O5A7yrOM7tcYqYnpKuqJ9rj3TTS66QQJpa/RVWmHyOSJ4tmP
vOWi0hVPheD1zCuHpRvF7y0ECM+hfmjKkeWQb8N8A4M4rRsgC+UXyh0/lrQAiB/jlP1kmbekS5Tw
Yg5CbjYieU4YuanhtuCGZt7poa9jhGwNPv6QjFUlSJxVz/WGU+aIFw0PwyjvhRm9adOO4xroUPbY
oRE36W1ZZmdjKHLZb5BqMon3c/8EslsoMfCFESYBGmhdox7/ezXTyCVI/2PC0VSbYnh7zZ1ubwlI
UdkyZSJ5srWySe7hNW92ZvhOC0A/nZxAWwO/V8xBmMlscv2v/S5vie6iCYJX3B1QouIu9LAzUGUk
QfeJyWfqVP+jyPJdBfpqxYCvoAL3/BQBrwue1ku2Xq0wtlxlwNwX3CxQMeb24wF56ZW4FtFdmFuD
sGw0Qhc7vgu4oegC6GvXhhRrmVl+zJi386e8hZ3GyVOR+mCtg3KAf56qcrH4Sor5iBIDn+l7s+aJ
Ut90ndzcdH5tHocWvH2zMyna4TirUoZC8x2pb4a9Hp1aKfgnDJlqhd3cSL4C9tCdIzmT+7+QCYVE
75lmiDZwAZ7be75YkCRpz1zseYoKGqBA/AQ8f5fDqB6414KH/yyHhYtT4IdOXdLHys5WRTQeqk4A
RyLELI2xCt0QQ+fVfpxyt/9cIBsle8PUSRIUcGrL4Lw/4jethU+mqijZkGqaNGnKIbN3kHK1+90r
WBHhQHvcJqIcUZ78yzsY3NkYBcdTcT48CyNwthZeTV46zFaucwf3jHLu3olPsg4eAZFndj/soOFJ
RejAwVp3r+9X/to1jKgl/olyx3levVc/BTCkgu8t20t+GEC2u3UmLy1Y0huAHeHVB1SrZNSH2get
bu5lvLEdp6x2snQhcHG7/asOt8/k5Mqg678UyAdPbSreu+JlYoBqgW0ipEyXDY+5BofBLef1Ei5H
LDzx0dnbtqUcr2sK8CDUeUZMZNgpontEekEQKywHZHxoOWGUGxxxphqE50Q6gQgZ8yNSKAXlspTn
ln9nDaIuVeKAhFsB7MRx48L+4dqC02nQHf9VlrqFfZD4dF9TDC2mK5uQZDoO3Zutq9HYPEQKiITJ
ZrauuuJD0z4NDBGSTf7iyQcg5vwOeeNucIP1TVP23O/zWhOKfPtoSHpdZ8EwYYxnsVhjYNcpNSt7
CYuGybb0hpFwVxBzFe6RWf5UkAK6209b0FUi7R7CyTJDpdM0cVcL4kje25T6M25hhHA36mXbnC61
0rGqWEaSKLVK0I0lOq+DYhYIGmwrw+cS7svGHn4nwqm7S3AtYw2HGZxbBpqUC02Wos+bg8tBRz99
mt/aKzt0GuIaX5P3mMRCJXjZ6HMZgBWNxwBDFAHpnuQ5K3ZF+L3bmfBj6im8K9MZKbQIdn157NoB
XMjVn1CqEpW+qdfTxrChHqUOB2IfoHIrMpidlJiB5RvtVnc+Iz2IYWaaDqiT3bFkI3TAE90d+QdJ
VXJzFGnRERf60udUIu0xdy+GEpBDVPZLL7PyWP0aY1y0cFcQEiJ7sPdn2z1pvil+y2xrK9qCab4y
bYwpt9S1mOjE0+/7iLtTD6Q9u0lZ8jEC8HKR8exqNwL/uZjO8fehJn5xq8GjLnE7rWebjg4QaCEx
8BmpYHF4Ksi6GwUuJxEppfuYTfcyLGLQMbPgIr3U84x9VpwQ59xDbvfsXTXQ+H505I5CcSwNceHq
JgQeyjs+Crh5Ddq5CXuG4VWfBXHWX/CszSv2sK+vCzn6cut4riA5F21Mpi+Vq6t4zNZqEPgq7bW0
SQCLS2tDCI8GVKIkX0gMx6A6X1psy7iQHEl4UDCjVrd97p6t6t1U9fKP36kMUIQxdwm7o04sMFna
Wp9gUk8W91OYDXjoI5henlC7RqbQDTlNaaNL+OhQ85frQpXxGuITpMG7/6FgFmjQZMfMWfmGOUBi
cYCZN3hJ1XIkF/mLNQt313AKLO2jeeVboaHVXbWymFKHkaQjVK0sNhnCEoS4WCS536oOz0zyF8IX
wgceeRxIC11XV8Qsje+Q60KZSZkeH5lYpak7d3pol7tXdhQDZ4jMCtXuwnXI9MJW38F2OHM7Slek
hOaXdmMM8IDj2kzOYvFPFlhB7YLDVeDs65WIyVahEwVTHjAxXErr64DA296uFR0tF8bD2EwEuQoi
v4LGa6ULMt++c9Bg+QDyajf5d7ugLAirXqK8ZlFfGw6CNKYeLrY6buYGuhjQ9AT6BPz3PRZSFF4/
+kY3t1U4chPQjDYT0CVTEIA/lm5sQG+Wg+m/Ztux+icbavEUFcqoS2CqY0s27xH1rDsiZqPmbN8h
ZQw1kx9RRXTss3Aht6eHZ4gmYq8evbWf/bw0ZNb7Ulz81JSGhLIdnOQtxoIYTlSIIqmvC9p5RuVn
JBrapC5mHcpAAmZLYHcdV0Bzo6SZwmGA2Fen0PEoyvVEcfI2Rtga0I1P3Fbjaz7dVpzyhaAr87Em
kxow6UBKV9pG0iGs/VL9OUeBoKfbOfIXw6SfgOxFzPQjL38jo1X8Gq7T0T1PM8Toiba6NUbBKiMu
/Y5lJnlcgAkCkISv1lffPTrEaD4t2ptqbLgqRa788MpnceR/HkHCTH3/zWX0IUrsr8BXdVhWcfRW
MmEvBZk9tefoaf8D75hOTkoPIWCL2HLHwNFlza6XngUZotKC3nc/0Hr2vK6RF9nFH3NrqIMEFEHw
2wQ3A0aPEGeg5pCw/YJMSDsrKRJJwJLGNdLrE6Fo7NEJC0T8pJuQ/K8kyg+1iqbOv9BKMlq7mL8Z
24eLTfdMV7ndTBpyWCiGs3El/nVWdJEW3jfrAVXEScvW2WIoIJwBG6yeLpuf53knNs9TN2lldY+d
F+SCm6AiOwlryJopkK86SnbuhbowywTs2w3iRuq3bhWlHZ6E+mj59r4vPJxdOWgawqaeK1sR9sFJ
QcZCEKH3cluiO+thgUfiY/lpOq/j+NU4BsDB1MT+mOKSkrdQFEEHNy+ZuszF7VLIERNk5kY161ZN
juu+l1K7J+E7DfHtiVZYzPkHDAHfVphICHC++90NEqukT42iJkffHKPgH7W87JQyWZarlYObpLYY
qpgcHkp9tY1xO91eEL/WQtO6XF6Mh11HcbChAMosfegYhdtPKYtSYDuNxkQh8Fmq3zATIcfa/RjS
t4bKdrcF2yO8tXhSaDTvieF/GwExC+zKDaRo9loBMx/zqx2tJ9ShWJCHDhiN6qI1VoIK+2j8Nds5
AYH/aFX9Zl82aq493pQUQhXlV+o4NaRufOQgSkW2pUCpXX2C5YRb8MKCLd8vAo44IGxsGh/sSqoc
/nUCXXqP9J0poDHC52t9MM4UO2pdkubB9KCc7gdBl/5BTxiCpU5RgBlMA6Zl/kHZPZxL5Mt18+Vs
w3Xu6Hz2Di3tEaYx8K23UsnMSnOip/TxdJ9Ws4rjlqR8eHQDV7iLe7BpAC58/v1Q9mPbgz9Pyz6c
yS2Ms7wcuusyJPWkFFHtk0LSqV7r61zXpK0seXudO4QOZL2w9EDHur6VyEzPRGPGD8R6hGcxizYM
SfoNyxZgn0e8wnor0k8XNIq/V6njKz+U8bGTPBviPhSzzz4ZPcNA8oAr/3lh6m50NeLqBEmwjMga
ufsQp6vVTWP2T6nkZsBji0dbh9Moi+t9JI0RkDZfgA5jDrMaD9D4888gncve1g8FfAmGlp4TCUm3
XLQ2dfAQrfr51mMPs3X7m+JbK4PjMJF3HCRpXvZe2awEPIZ1FYr6La8f/44UXtg+3VH+9bid5/3v
S2wLDRJ9lTOO2ZBa2Dk8pLI5DjLa9gzaonVAvLFqYtZZsK0gHCdN4NqCpTmJdBneoyznLqdh7Vmv
Nw7Tc6Ttk7Hri1W2ew1uoAaidvhpKq9/zrWFWZxuMhaxSK2P7fYPme/iIxYOqOPdG63dEGDJJCUn
W+oGa4FE09BTk9iDZcwj0++GdW7zV20FqPToAM+A1C1YdfBU3N7SPV/Pl+cZzfGkXgT+735VxkD0
3f9XBHm76m+XRKn1vFhxCdGAkAsTxRHAaVyaE4EsZx+O59D5L39QjJK418cFO9Gzx8xrWDxAWYEB
Wz/PCrhbI77Y6nJI8z5mC2NgEI1PnU5PHSl25vAWhFnaUcEbt40reAjl71DbXV6J2qbKvxqRRfKm
6r/VJWm4CijgxQWrn25k7EzqIdxVfolCarTY25yYmiG0pyrd617qymh4BCNdBXILVp4YmcIyWq9+
D99mUlLMahhLnriGjfZ5T+uo/b7GT9aAee61O1Ga2I47f+zPSzBVYXoCDTyMWWmOvdrC1Vk74f7V
m61DN8d3jGP0CdVGi4u0LELp5POmTLlujTL0yg40Aqy9G10Lw068pK/ucQXZ8Ngzuxaf8CMQJkNg
ITxIUeewYH2MfKz6vaWU7hsuicyp0kFXvCJW/f2mgfB0CV2BUgbtbwFYMnjzQRlNX5D7RhIsqUou
8CeEwgeeg5jrc5ivi7gXhDEx9hRIzaWY0EAllxAPm8W4VTl+ol5lmNrcNREzOrE4WPVosyMRVOxm
CqkpuwSAhOsWW3V6VYJTKCg7udtSPlUZ/YQkoLTR1F9vgxpRXTfaICNy11OeX3MNT7eSLg1+1Qsq
E1wbZ+6o+f6gpMU6NYGJDlDIysGOc97tcWYrOdiylRXI+BWHKTnoCoEodVzFk2DNKX7ibRVqpgdg
S7J1RDS1TCCbgyDGVlqT57oui9nmXM1u9xv84Itx3FjrA8rPPuixMuANTUf+5M3yW89BOfma16VL
FfomxgFhBd3ojeAPkCPWPQPYJwJ32lt0RcCYCCPdFqASNoGcM1Pr3jW0x2+B7x4sHTFNcsJBUINd
CXJnDItB0I+zj9mvJWfrEzm8s792gclvJhEFm20xyeabVGBYfxu2il+MgtITOaVG1BrYENHWa0q6
+HFy2wl9qukuGVCZ6aMGCjzHBWr3TUjm3j56VwqQbH1mV/FrSWonSI3OuFqjHNmjAUOcT4iCwjvy
wTgUs4+xdo3WPWysFu/iNuGibLkdPgmonRnPLeTW30a8UIC94F/a9s6GDMPy5J0qsdvmLcc6k7vR
iUPJWZreiJQIj9BKoGs/EBMh3gh7rLBInKqYCvB5vsSyUEyWBsD3v0h0G+nYadmOiVq2cfn16vU8
5INV9AoSdcV+o36NtwhQd/DsN4MmHDuSxW1k3cLUE+2tL+lK19G/UtQ7lOWtM7R+//mv3EB22jT0
QkOaPPmpBgLTsLvoWVqELBQfmguVh2IkzxXttE0bz0aX+Evfe1MvKW+sndBlGd6ag2qT0DiVSo8K
wvd1V9Z30FMuFvXV2Umq10zWOTP8OvJ1PW162hUYlgHeK4BRRdINSsrnwpUUBiJXy0T+058lQuIW
7a2gArQQhS/xKLaqFEkQnTAAo8lBNUVZ72jbZbLndeT64gsdbrMxHfHbH7NFqat2T2XtWKV7g5v7
jE6/BK9jAFPFeY1IneQFIWE1YZiSYQWaDYzhhyIRQj2AEjkEG5PD6xhphdbXXL+mAGPExTyV63ck
WOFJmSW8Cc3Op8LHMlm6J3zaACsre2ZTJ6MHjS0PuFdnOzJMHjgUEyGyEh7xQAwr907n4V3Bg0w8
vx9eqVtiRph3TkSg5vnP1c+tD7Q6vPzRboRYP8HNha1CsA7OVM8KRxT43RX5h+PNsZI8puIvk0dt
kQaz5IkHwKB2KTUfdBuLqWLVdM5BN9cI3o4r4gWeRQA4FcLCNVRxzMDRgz19yYxSUdyG5niiSSK+
AXHs3cM5wGhqSBhlakGxATHGvSdsAlCMb75pf6fhlYlwCl4qQ0a0HedcA46tOJsNyCmkOCqnJwoD
Emtp8kYJkEmixFygwhChWtIi0d+97ETI5UvJIRkmFlCrb6ppmKKgH6+ufHAYb0m2iLb2wnScBJ22
6iNyP5hbqZet0jpHaG9IYyHVp9HITkaPPFzoA8RDLH//0h+X+aODJzg0D9GUmPNl+g8c7Was4Gq1
3vtkaAOk9SwH5Iq694cqo9raFOk5w1VEKG1u0oGojqq16YRqzCId32ZXpvar+TUqx6NDl2KxB+Q4
omqGdT9JOeslA+FtJvDxwI9SECofmqlcVDT0dKzaFPubKVpoiFXba3RTojpurly9vHqjZDoj0znW
TXg3JTLP1NLosiymDwi/UbG4gBPDXZwEHVQiDy0xRn8TawkTIpESHUoCAuAHCZRKt+dGjDwwvp+Z
a2kaUOQlH4kLpIDPNVG8gd45r2Us5V7yBRA+gjR+FDSZCLOpMBkLrPFiM2udCaSWxIOFr5Au8FEL
ckiHauP/cOIOQbfPuKXL0b+rH/t7SenHKQQ/9sS3ySHDW1C/qJAQL0KKQxHLurkiyYHLq9HtBme0
H+3uXoD54DlR2eJG50u3ScAEoZOGctCQZGiz+xrIvAg1XKNGwaMliuOzdV2n7hX938RkUHo3k5Zn
Hq8vY3N3FLeoUD/L+1FjhBJusI47XqF9WdWP5wzRxTJJSf788qpc4B0ITHvGkPKCp9WpuiER8D/d
prJRqk8ufTp0hb3x/oa7Y392yeCyWBeZG78rBhsH3SGzFPghpdPIvfqFfHV6fzHH/gHY08ubk6eU
8a6JFbfST1aCaOFRftHOyeTOYexJaXUauwR8eiTsHnonzJjwhKSi/I9hx7vL8+3CbvLCW0OVf7De
DlgrXYmkJ2Eu3zVEtvdmpFI34B/tQDbLSNBHIKXQGxCV+H5uI48FObK+K58wO75OM9ZuClAyIx+w
xUz/CxFNdvIqiOmLroDVGIE2Vx+J91AStZH54iBJFhsqz2OXzs4MqCDgkmhqfa2YG+jGfynpcWLA
uYsqEjcxkxELRKcRuXiMuuAVwlICi6x/erEFiYPomHlxClQTHmof6/kNgDNb5DMYul2bkY328r3L
HDIGhRbQFf1UgtHfFdTL5MqZB8ly/KlIZm/0IErvAi74j7Gc+0eaDeLqFPjbgMZ+Tun6iDiwRpyw
PaohbVCJXl3lm2ag6fzZCYKTQ//bNGzt/WLuzaIcv5JkV3xN+O36qFp3cljG8FhxSN0tD2D7N+b/
LZjOTYwhHTJNIEfyzjN0UwI8db6hWoxvPNsGcXrWjBi1iSDveDzNAsYIEBZAGQhNBEz4Ic8gbV9D
e8GxJHsrxME3/CKt6O8L7HkbpRKF5F4XGDWCNGPL//haHv0JM6c85vLhKj/xwKDcQrsl5J8A1xsR
KDhKwCvv84tw+aYIcnt3y9RurdymBB4OziYtlXvN2BkNENG7vxsgMz2mHPxxObp8HYfGnj8CiZHO
U93xxYJMDyQv2Eo5NxvMzd24mf5XTkE4ZaWR+76ihi7nTpylLkznmOtTsmRlcjOCNz3VatgT6fMr
Z+lbx8PFNEOpX5ixiSVO/5b4vIte1f52of50wFBAjfuPjzDxY0Lw94w0TwHv/5mkLmSMIt4hiPd+
gkcNXLPLY6J6x/GTHjIcuxVXx9gcpN5EGH4Sb2WCfPikO0n76qtn0GSA6/EbeZ9ZOfx9rZWOsJCA
UcGM0wwPZJKqCTwZHHClHtnL23qZSzG7v+QAI5n+2kf/EAy0RC4senv+E+vdzjbwiHoFC3Ru/GV8
kkpunMcGXzhkSIaLATob/L02aItx8z3YCcw4n4ByWPtE7DMMSxkw4YCIyMOm7U7Bgzfbk3nRVDny
hrh+ptR0G5g2Rbq0vCv+4d803oVZs6N9ij7MvFAy1QRosDMlPaInI2alaT8BVLQ+oEgvA4tgQrNz
Ntmik1/rx8FqpCrdKjknm5xLV3uGGyGckmlOKNlbHVjaoAHZzFlLNwMDECr9fn9R/Ar+G0mcUmZW
hoz9wk6WqzJso7Z0iXi8LL2qJxkj3xBWJZQsyC5XeGjfprpMtiqe5KjxZYmLi/ko+0IAavhtQk6u
3DSjkK0G3XnjeFvIM+tta+LILPLLrmCsMUAVu4jz5/1RfLVi9Bm9aGz4PYooXEt+OUSTmYLr1n8r
3BpgNPB5nNIjAP2qlrKDycyUiMS2rGfGKWoin19xsO2lgyXXgL7V3KiJJu/6DXI4Hh5SRNACn8xu
KyXe3s3yhGOzQCd0Tp3hWpYYkL2BGzmneyl/ToVphBJrqzf733t94YRsLpKd9KDsNAwibMMRHSWF
JfQ2vSJjtpVqF+kayaQqOyRTYtsrzU/ZeJ3v1e9PFrukfzSBEfDFY3NT9FSeEaOkgIYzWfY0vOEa
jKkH3o7Leh8DGmyq+gkNsUJZq9Mvzkb7fQ4LreUwRhWoQYdmofBUQP9FFqu5al6RwjWAFUa4YBKy
STE/qniipiFyxNmi5TdKHvjIZe174JiLWG1XkNeH9304PuFTeoSZo19Dj1UpzgjkZEUiz1Ej9Nck
xHQA97+osbI9soAPkgaYjH4RpTGmXiBnowoGX3Z4M0goyHQYnwahcQiCXEfLpmdN7ZcUtKSI19nX
1Z7giAVuBYVjhpqRLC4vHnLTIvqjP/ejMrXLB+rbCrpW8vpV+Ds+bY5D1GfTNmBc+tVdrhQD0Lna
POkR6YcVVOXhLj9h+crBX8L7a1N/hhgwaWbidwTZSC7RgB77yejyyFhYL8xxELQmTh/XxZSnkxlE
HCjorqrVbdtmRgiUvMGDJD7E1+0Y5F7+eC5HQmSrtQ2NeNRr2vwPFIsekM5smNKSWEHEtVkp4WHK
Rwb04cQHFDhvIfX4ZmAQOOI45LENQnVWuZHOS1LlmF5okJJBlfbBqxeVxJK61rMLYPab7rfGu0hU
/83Zxam4tzU/87ihxBDEJydrcHwR9LDsFmx3p/j1ZoxFX3+8eKV/tKzlKHBi0ML7AFdnBVz8F1oH
9npoVN36ao+3ubfdXnoJ+ptJgpQ36POKnLCnloTdkyAHPnW9sNpBfsJbhyIReRNBV37EdnpXuhsW
WyPPHFm7ufuv1TID7XE+9c+nzhABqii2ETLrFlFlGCfAm5AVyz6g46psH2CSiOVIo46cLMfYgYeE
ctBnNQgwdxj30TfRjLSD2UxyDLPcBO82zHzVFN19Zb0DSpJlpczb4HO4TK7cDkDtygehWGJnM/S6
pm9vxMN4u64UpfUDAb6Byp8lW3X8glWMTzWXVBdheJ0x/TEKuHdF8LXM/j/aCtc98NPZ5JYlpyGn
cKDjV3mopLaWWgca0OSw/3bBYJdGmYKDcbPcKtVgIVxG4BAi0+Lj1xIVK8LjDJUvtnwaTJno/+kv
ywH4A+oJKwk67v2ztzx2T6T9cmBCKIGTA84ZXC/SR6dUqr5k4z4+iy2LcXVIHTHq+U7mU/SrPHTt
ynRwevQJUzG6gv1qNRx0mjAjJHbdpNlO4HtnOuK6PCbFvLOFW/V4b4YQC+5Smffzn6EzwP70MTM9
alIYYTqSUSKtP0/83FFwe1CpkiQ8PNnqMmGv/4WUhoJmp67mhylVmhZvbQogNHEq4dd4RPaMUjyy
MjFAonAW8qyKPOZJrHKoHdzcB1+UnzFZFyhIhthplY3ZDqfqtH5Or7m8F/1r71yVOTzsYE1pXngX
uJrWU9f2XfaFpBD9pdoO7ecd8oGugPskChFXcTYXBDuvv95LcXIoCAHjhn5Ttbata27kGtu7UHrw
lK3fewc03ISi2ePrMfKVd0+/q7Cms4SoGADGmRrJefnVKTtFLK1VjhaK535+zxUve9MA7B7Etp/5
dX4yv5oOf3Vjb4YTj2cJgs1qr+YsAW80YPWZYxkJ9uG3PM43Uc29KVlVvVv3IztbkxJfAXb0QMiy
js2prce82pONkzh3AjPa5obLLsBO93iusuFoD+3Il7sKD1C1BIGRg/9lbVMSy0MXkjezZuM9UtG2
xCfWTct3WkoZRQHvXwOEtXunryKW/S+9xjRCM5AhWbIGwxb1oxzExnIicIIZk7OurDpB732VttNO
HCQhiheIkUV37AkBr3O/UxHfJApafJzgXFNYhAowQAqMbWn/4VeH8h1MHEZgvaLALhEi0ZlnAQf+
iKdpsZ2wssDr4yiNc860Wv2nIuq3iKwu7XDWQFxvCMsyqCShvbra+RNvx/cnmYGDu5lIuC1wn8Xc
5VsKOZ5MbQPplPUiIZngmDLFnv8pEBJL3a6wozkhLIGiKh0DQ3aTbi4Jk3YJ+cMSLn1d9g3NkOMx
LuRNd89H/aZ4aZ4wQHj1L8RXtDGRbkYyDAediFBhKbLqIWLb88uKRK79EzZULMF/O2zRD6dtE8oe
x59Nr95/ifMfKXsVdi0s6BeGNoqs0WpjzRLMuRALV5e+FnMfO8VMTS9igBunLILV/YDuVuZeNPAT
zUMl4Ce982UrMNZCV7HEibR9usVX/GZhGRqJfbE4BZU28OMXKqT+Hu79PI3Ad1gj6JvnHjGoXeKt
P9vEvDfS1Zo9aZnEBnpZnOAzbWBSwyvh6S8MIH6FumZOdrcPKM4gGME9gfG54Pv5EpRowRq8rPlw
P1NyVflLalr6HR6wEHioMYwHlvIzQ3ZrtYpgQWVtwDN1bdczyRhg4Lbvi+/dJsg1FhbwtmFX2qbu
eI4TeXQtotsfGFGr4Usce+T3owDk1uaVDTOD3x3xXiCm2jIab5Cv/yyUj7IRK3FiW6PvL9S7CszJ
t6kH5hLuQe/4U90N4EBlluhWSw0aE/vrxFu6sNbM4bfAByjsbtVak8efa7uD0ng5hMVoY/rSY9y4
ceAxGeZj9Okq29rDcNyJ9/Vvn87F+uOUJ8zQH8MSfHbg7R6hzaELUJWyqXlRO1COEQKBLRcCwxGr
2c2pzz8kn07vYfRCQiwY2P+pCQwhL/M8viR+nZ4bc3zMSL0aRmdsC5yKfH0FVeR5z+5u24244uqY
+gzQYA637XHW+/beLfUYF5/QzZQo4X4C68lD9bPoni9O2DnI3MBxmBtMhr/6FiWuWlDNFbYuKGrG
vKt+QVRfgtbX/fTdU6m5QyUyeSms0P5BNiQ8kx6OkExQyOTiE7NJxD4B31kMeRQtcLF2a0kvNTvt
CDMUL19uLsNFlF58F4shsk5yL1XcSFHgszciJrLd/Gl13CwYNysT5uZXZEeXAWCeKk36AIYFPhB3
SbFkPYeiCU3XzBxsMGsKSd1jnrIiIJg/W7aBI/oetwQJa7+0Mkvw87nvCZdFDAgGsP+HhqyyhUF9
7iMBQQRr0HctY0G4v+45AfSfahpIt9Dk62IXMptHfMwMsnIGQntegAhK3UaYyHNhK5ItwLkc8gWx
34fyfcDMmXXFD9V19n02CU7YvmDzWaTzHPF8WhuJtykPqP/xtbueh6OG7LtkzMSiT0xxNOhXISAz
VAQ3P5KLHnOw7rfcRR+3rQxCFDue5kw7mUh37h3anqNQcD/LQpLXxpKGRSTS+uXbFAyGoHFH3c2G
GfjJBM0V27TMZw/VhOXjucXaCZi6T2bQUpmtQgSilOX54hN0fXD83y3cAu6/69aJA/3bZaF6vPQD
nzaA7ko3em+QNrvvS6+1xToi2+sjEhMC/FPrYMtTZJ/uwBnESV9EMXbxgv5p6a9DuYnnBb61Bt5K
68+Zj4HKNPiOl+fmR8ljttKKQ8gBmypzpn8rjQxhTUBvI4toWp3GJe/JZA6WVsGngCbo2Ho5YmWu
deb4FyscyeDPn4BOSP9lGjwgSLT3h7d6sOIrz8tzNhP6BQH9VEjBPpUWYjEDMdAANFu36t50i6Jw
narPquyksO3+tPtq0QD2vJil/tycoK1cPE97nPxC+N8gswzuO//3js2oNxCCPOiTdbiHYgXsLq94
zIWIMRiHjZfaUOheRN3DNvKH9b3auIEynOBVM3WiP0uuy5S/4eEYARwQ2lc4d11YIiGff1nFpUQ5
8TPwCWKaipBY24j8XFYRn7xuN106vbBsy5i7tJ/6NIUHO7WFSMrJtLUPZY3s3Mg8lPVuWJ/5wnWZ
inzOcPZzvMOPDK2Ntn2dPTfrL0vpadwteq6r2C9GZldeaqyX1FaXZ0LlNW2Se6yoVfhj/uJcmcoK
On8YZOays14NzsA8qsS7dxTDByrcsuAdRPMltqjzgUMV07jNoXeRPdmrJwz7LT+s3uVkMa3F8xC6
NJoqdAo9hVHvEABh26H+vWl7yUuGOzGYE7gyX5kTtfTVFAVbClHIsAsdxeh9NLHXk4sCDmaLQonB
oZbN+9S+Zi4Yxb2Vun32J+GC/X/qNl6u0d92ALURnNMl9tC0KQarYgogiWTXp2jLYzBXxI5JHGRf
UZGi3cfl1gY4TwLgax70u+HHeiv2Xckg3+OwwgO2GbH2AKyrffq6CZWmjMNtDvSyJz2nzq8e5SGC
t+hCmfX9J/bR+/Ei/oK0Bbr7tCkeF1O2gJfo2qZrmkTg8BUPo9WAXrRh9oYrRE1z1iiAdQ5yZc6y
ySE5nexXMEah40BJyTAcWzFOONQ/HFzB5faNMRwBfRYCkCyVCJu74iieuqsSA0EH7iAJcLnnuMRp
IaCnrbigWaVdm55u5IDZ4wvNKhFI6s8A2AEM7zXMGnhUEDvGG8MlueTPp8R2nSapZl/VkTl5GhY7
YsscgpQMhMNEORAkpIV+jmsI4Qxa2YCgiw8teTXzejtNYZbMn0Y+jonXE3XNUKjsr5PGZ1BQX75w
eowOxl1kWbw9mVA4hBEX1OYSuzqYPTnFLafaObI1SiTxIHK00hjcoUEF7WwEh3B4yIUNMnKgDxTr
GhTonOgTHS+Ju0pOC+GpsK4NBNnxUwKLu1fPm106MN+te5AGzfx66hVOUuQU7Fezr43CHZqMPxML
YqZKmbH3XUJzjrnWguccvhwwG0uMurcrUgT21+NOSLDZyW7XM74vW30TAAltoDmZ+DXHIb/+JRxB
jqSrJGMqZjLxWMHd9n+SgFGTZyNhlHAyVpCo3ZmufCr6aHLN24qeFWltt+CRFoy3c9hvvM+tmPiR
KDFaIdIcvSbJyO6VPQUS8r0Z8G+fdK0eXlsm21c8BicztmpHEDymly1jODqhZuGLZnkh9euffKGo
CuW/HBSIYSAn+1wKOS/p7LJexN7IZq4l9xo9JtU1POnrCAPFjcV+l+nSWf1U+aCxTliv8qrT9h34
mQGyXgUoktWl+mN9B+RwU4k2UVnHZf2Y+x94uLa9RT14M8xzJCp4zNSCIr+R74vy+EoToY5yzUsh
+8I40vTZhLe1g2/ffAW1MCGXTZXHrbSbwLC6FHZmyqWQIRNCkxhH7emg+zPSLBSyG1qVeDhEuO4t
fDfUA4PFTOjJE24af0o8sSNg8Nusu5cQPxg9JMtvZ65GTXXvfg735gW0FDQOv719zCKsDAaafK+I
iHRpWgbi/LQCyuFQkeaZPFLRVaZt1qHm1XlrKRpX+siNeT9vQMfnbYCLDQu+m+Xw3RqV6uhyQI38
fTfnRgHt1DK70qLQos6r5rFDGDUYrgHjhXkMno8uV2Gv9zZwH3pmZq4JXOUDg9ixcziD71ftULPY
ythYHfpQ8dy9LBEWzep6BVyW28ofOQETUsFcHoYi+l8iMnZeiSq9raJP/dd7PEOtagE78qdOvt+J
boPNUCPxuHGRGYT7dhWyiK5MGKE0DMS/dcfrA+x1S8CPRLaRm2RcQ+CP9qX1P7GN2L+BPhlqeffh
KnT9ZeQoS+z97j/BGc57cQ16zlZORbEiGjYplR7kYTlvigVNsT5IkUjcK7h1c0/2UQgLcfYuCewF
QCy1aAjePPi8jKsm9DaVWy2k5Trqvbf1fbhSGkV43rB0cFOo9+npAXNNrjkTse3d5pF9vxU1/7YH
2CUgmybHo0gkFTqLwDVbWwOCD7PHX2NtxqclegAOgfPYuyrhBMqbhQTqK3EtNSvX+82L5aVYEPqO
yXmhdSnjmjSch5k4TNXc+N3bD5efUIG/lHtUhjTMPJEFN0EJgR9mCMy2YKKQZ3gsVgkOffZH6lhl
IY4pNUiGvZ7oIKSdxLSJU1rZeZaW1sfIdGfLuuZ51x6qTRfqNlllvL9cDgun42ezTEFbdZsSHiZl
LaF1ryEek6Na+gHjYH8LfBNRLDLz8KqLQ6cS77ZGkxCm1jZlKkdtUpEEmBsKrb3DpAeuebNi+z7a
8qQ1q4oj1b15xya3XyGP9eBSO581LLTwQF3q4T64weaBihA32dlgyA5gp7C1mfjQmL//OnwFO0UF
tbkPmcFKavZzr3ZPe+zKs5rKcrsTE8MSk0OxhTItQuZNr5Rp2BavUbnOLvxmd+oBl8jBHB4+trKW
F/gS/i013BPNgLZHWP1E7iISuDkpzF3W11CdVpsFx5AH6DBIDeNCfVVh/sH4dxYzf/JsC4GxEBi4
3z6PjuiJ2ZSm9VhnWbIcQ863yBrxXgUok3px28/1hXgw5seubzXVOL5wyHxHgGsHG/rZCyab5RAl
ZYY6cDJHDHYoxuZCuBBaLl2yUQpaZCAKrNVSa/ZC2LiBgyWKhq1jPMpFIjT3fP9EAR0y0v6XGq2B
+bcnG1rP2IyjCpwwaYYxHLObmxVtd50v3jA5YgL+C5MfjjW1N3t2dUU193dxeOfotz80iFYeybWe
Cyiv4Kjxb4fwnFrJEFTbhgeQzkgy+US6jNDqyHiFouh+ed9BZTakJtL1nuoK+lGaV7GFQeujSOan
2NX6ky1QfiHXAsfGZZMrpwGJxp3/ZMY+z1UBHwNUO3+4a1FTKr5gAYTKgU3uRCSlpTQhKv9SePTl
Vqt/DXRSpdw6ICfS4XZYlRdCT7yZ6wOYmSYE/q3RnVZXBRtu4ZZN2+Tz1xZRNNZZaJbkcDgm5Li7
woDRAQXcK/1CL+XBkcp7J4NMX5PDCHF4ZyIsMw0JRGY7n9J5My4geRUQDoSkbibgxQcGVipayxtA
SpMSxP/nwzvgU4gF80poTN7Qv73iiYsd7N1d8ZPYUMkoIAGbUSR2/8gojabQEdBRjtGGIqYAyDJ6
7/xALm00qDvfAV5mcTbpHaxkQXMENAtyZ2gYrzkfcfA9igy6dWIyUoCKnHbAyJ8E3bKRCbM+Ar34
uoEd+e3v/jmg0XftNCLuLsJbThurbfcUqts037NvSf2bEk9Tuq+l+946pC2xoPfVk7EW5EO0w8ia
GVYszY28rH0jp0PHr6tZja5iWMbF9mPScKh3pMJr3/NAX1j+F84jVYS4oivWDUTMLeyCyvVd4Al4
xSfoNIM41+Lq/rj8rTDxR9hqDPp8eokALGkgOy6GUqPxg2TCkzCMpTrQe3upBs5zaBr+c8izwAQA
zxRr6rpH29NG6Yucggp2Rzn2q6GOYt87daCocjv6PQjQX568IF815P6MTrbTnKaUK0qrbTfLKiHU
3ReeDKMVJZ9U6iKQ5ahFetznDO3tOAKWjvvzHzuE8xpD4uQkmWzDdpB3hS8QfSSO+Iw+ayTA/hBO
OZmiiN41M/PzV2DIgCrXrpsss0rbkaYu0D8Jx9f25utKQqr0RikHbriloOA1/1s9nQ+DZ/dwnWBD
f+IAyAZCBgE2cAt9MCHOYG5ooIqb7TkaVHVfdf+FonaDPe6meOhHwXpPjo6orcfxOR80SySExAg4
Q0ch6XvLNrlZ+v92lA2qP/b05C5+Xs2QdT/fFUfYPAV5Oxjx3lXDdVqvSeBsoLiieAmRf4e7ZLgd
BBAC/U2DAmLVYDIffF6m8vDMhP5bbccDfH/89IS2TSCTnHtyfPSTTmqKvlONfe3/qQYA/I4Ybm1c
6C3XBfDoCVrdNYv2xgGxe8ZpjEvxC49ULz87Na/UC5zQCmtBbC/aNbwzUv2KHYeTo0LJAD9ou1Bx
Q569lsP2Ikoz+1NHXnKkvfVWYxWNM3yZp2wQvdTDPEmPfnvB+VrHNRiHQYb1f2gPWE4QCnzrirem
FmL5YeJY8jARbth+Nk4kbS7idw+czMf3NZQNpFVZw322SHFuQ6LwjhF89D1d+yyMwAEIdOpnQr8Y
Ka9Hy2KHqUArLCMFrUNPefPlvn1oN1GSP9384CzLR/7wbBf8MmJTALrWub542nz6+m/X7aJBnyFh
R1ipeZBFF7xQanY7dLu7EUdEamQncJei3Wp2beY6J6Lukgdxwv3is5RMCrofl5xew4vqdM6RHsAb
qml1KP8H6oVRXjFUF8WOpAVxawko7tnCBL0clE7oUIt4KRn55trfWbIXxNQVlOz5cxqkEX59W6FI
2YMzFeF+vqxFhaw7R3WJNctIsSncMknPu0QJdvzUi1MgOu9H4O7W14it8DUAWa0Y418r08qxlvkd
10udViluxlohYMV4dUp48LezUoqxA8APDwiVv6r5/kkyc+7Rgf04toGP3ZqYKFsD1KndXsJEy/9Q
9G0xc3CR7r4umBURJQNnDZouMSTuVCX5+2Jie13Vq9+Ios6+sj17tpCSKyh+IYD0LVSTU1SCVxDx
ZyBtLotZXwSzQairKWU8ym7BoMECW/1c5b3I/XoyE50c2UsxJ/uCCQE6JfbcmICC2DCa1vxZI6VJ
d2osxadJffg0EpI30texiAhpM0mHVrXyACk4VA5cx3K23KtShFsFW/mbinpf8nrA43iDFgkixBPz
jWKWVKjND5yeM3aY4KPP20sm3p7fECmrILLIrKYqtz9f8aCOVG7R7Pk9bn8G4beGMKuo4R7CZBly
vGS+k60BgPK+ZSF+34ASyYXWkbRZHZ887PE1MSaa0LSFDDJSSbB6HziMfeYkYnnVTZhXSvmuW+vl
wpsmuGiuNvjXLm8FjaIzYv/o3ncozEecOd9YXRnKA5R3WSYGCh4HMhDmCwEBWphe6wcarfkUuAgT
WNTC10Pk/9pCSjqQGIzc3f8QhRBZu4TOMiUoG3KVUOYu6MUujI6tS2EVvF1hRfCy+TCSfX/NwnhJ
yFlpxAyHh5VpZf1eo3fVT8dIv7XSX8GXkHfD+0zPec4zK7+aVQMNWM6oaugBHryjr+v7mGbobuYz
VbfwEdiB7xpuG4AWIepoYhjlmgdCYW0+497ReH1jWyS+nm0I/SlNCe1kByxihdizcuIO7dCxS6Gn
oMSV+LjfHlyL16/eY/jau7woALyG2HAMUqg7t0oG/xLQhaBoMeu11JKqj1dGGDyYKKF6/zgolgUp
1gWQC4JX+m3eEL642D7WbPyO2m8NOuQYq1MX3gAKn8SlIWpUHdpGgwMNbgDm0frRJPNHrJLMwdFo
dZQ5lNOjTS29fpY0negpl5xhZePU/s86sRkHoK2PwuAAgU+am4I+anoasP9gTkq1o2+4nNjVJQpA
Ea9vHgpnIknAHRjI9Ozan4pHEnETv1L2f3eoAOlWOFBInxZ3YOQ8tUTX+EHwv1UApwMBO5Xk9H6k
RsfexdVlPOe2/D7UtQyCu8TCdiNR19eh26oOePVLq23NchQoIk3WdN/tpQICtGma+SXMxJgdPZas
41Yiv5G8BDGunfFLhY5ChYQK3TMO36zRhM/0SmtOTyJ6OLlRNOEdX8Nc434q8Vk8OSnf0ZeiMkBY
AI2XwhuI6gWNw/wr3k1TXUggSqhiDv+HikR5pOOJ2Kq2naW6/dwC8j3h3RdfuzMUxLgeoiHY3uBY
J286wdJjzn9JrqUm1a/I/UXI9JeGgtY/I47uwpMvaplEbiIzbz3DQBZRNDB7073acro7S7QSebmW
iPDlEedNJfJ7BndK0A5RhG4pnVwhppJEJRlWuiuvamky+raZ9b8LdgByqcnFW5Ax0uFTUGpR4hAq
AamepxaEpk1ptGeaC5cSyFQfbqPLJ+n5iPCHP3rMySb/ORREMSk2gyQe+tnr3jVKggjaAc/X4lOW
2HpHUGXZSc3P4fzMI+pBVVjbROHP2xpmqX2VshK/rIUUTT3KeQpVixKsUSkEyINayVatTq/3SQyB
vqYfdEuyTq1V7plGLPRqug/4kRB5KUxRjV48mAKouMJh83W/my7pTCi3Whc1Xmx1sG53PH14RIh1
IjziZOu2BFpOUEGeSvgLe0MUZq6bMXAkx8O1uJBv+f12bv7zKkWEMsIpRhVClK/Ccy3prgnntz1A
/F89nzuDwsf8NRh0PXIasQag7VY3LfrWWjMdpT32Iuu5mwlgXc4AN3CGBK1Pm9XC5I0ja9878/9L
89M5/Xl5Cvmv0zBmS516kjMcReTtgaHgXXtIIycwtYZ4Am/Vuio70NOH16vb3NZlZkdK+WuvNwPm
TO5XLGD5g9ao3FMObD+h5FJEUUX26ApiD+iSzKev4QZcZM0GgBZ2XwgFauDC15t1w0fL4wze6PCx
6xVxa6UFQso3dzpeLYBT0goYawSQNRsQepfCsL2y/8GHkCfqaNJ6HzfmZHyHOEQj5HIjbVK0JAn6
qZGtKndLFC3Mc01An96SDU9/Ryn0fXMJKxWizRmbaTMolqqgsGZj1YkLB3a2U54o1tqEU+aG2TmD
uqCpZLl/mQWO+5AgLQnFakIfnlAL/5g8oSOhrxlsVh7FOvN2KPfgfj/JDdeCSowrWXnDmf1cZRIz
dJou6n5h1X+dFOh2jaKLnVZf7h368ZzxmXaQ0mLwze3SM2DFqPYQh3G/X1qdZE5VHkkP0GHnC4BR
TzIB/T0nwTrxViRqg+0j4VWaUPRypFUjkyjMPFV5bT6MWldVuJn5d0p6tzHZ4sWuTo6OwkjFYSeL
aCmDtreTERWRQgRTlWmxh1kxRHzXZNF8zC/Xkvf8rx1nscgHrVz67e6Lkho7qY+LcXdE6MK3mWft
jc1MH/kN84eQEQuOxxFpopfob1nFOvc6j0k42RVEtR64FqfVmjrkEywui2vC3OdbvnI8Czn7BWV5
IVcCl3TFuTtxdICz1pJWHLnaMEx1WX9Wfu/M99ga0bqTZk3LKkBEHaLuhHW867z/AwJgmm5QqFFK
/xqCa9LWmzC8RYcN0fGrV9SF3lzmtwno5WAqQMV9aks+5xD5BusG02m1UXtIpCifPhyLlxCrI7Zw
e/hyCscRM2kMYDoUCq8ShnpqbMfmfQH1KXm1EuWLnWlwkg+JgTo65IP6llOhYQKVfCJjoJoKYyGr
Erq3hDqkyVMoBf82+ztXTAr+nP68KSK4tON2an5f+570BftZ3YulHGeyUknSflZ7E03w/+J9FkNB
M6ubyF7tcqc9TgB2O4oGtg3KnMkPfhZhGYlb/LjQM6FOs6uIkU21winiTmT1A6w8g54jbPaqOI5t
XT75byJpdke/lTCOZhOG70g68uMvI+xxS4Oe2KA6WkzLa0E8aOV3stb3M6GAhOdUJlwIrp8yqv8M
2jjjt+yeNchWg/BOfsASu7F4Oo/oIdozW4EaZ1OYtxpMt4aaEA+3im6UD7MAWp+SjdEeFm+vnh7O
0fiKwh3vVNneTRqxRC3lwBRp4NpD0odLUTfSoaXxzOz+842ON3T+tmUIqJXWObYbqac57BQOr+q6
8fID2waCJHsWoRInhNPuwpamksAAZk2p70YxrCw7DCZ6ou/nCYiHlz0ti+a0hTS8w1wu81gg82XB
qz33lt4voxBZIsuc5Z7xeb535JBdeK75KELJQINpbXo4IDrAgybdCEd09yTn2z2yDSEkBXhpcBaH
Kj16wORsX2n8+VPqLd6jkyWS0abrikDVIaxiGnd9wN0Km17vVg72Zz9KW5Ci56gmYV4g694xCF5S
I5SixLSH1xQ5LxQvqS+EEMObErtnqf9XcHHlxdAVZnkYJ/OBQh07CJ2VwD9UoLfkiZAUGCdkRtev
/PRQpw69Q41SiscVLPvBacemk+p7df4K3wdadkxfNVtLcKExReoxhazI3X5w2MFe/l4JbYoQFsSy
pt0LeadzHQrtUThBTOt+H0hCHDryuAi9WT6coUInjDnn7xBur/UZEUSdTW+E6PHf69k6FiM3FqUj
XSPtyUsBFrA65z7xFUzt7moyPo5SRcIYcO6ypwukedfqdfffJtLZIv9Of7pQrxgI4iJrOCXNux8h
ZG+QDy6Bey7zWYd2DSVI0KXvTOG6MqfyevdtuGDTMYiIz+jsM7lVruk8yGhPMU9a1h4hkpFNqmGe
vtAM7GFTJr4iR6zyBFwyBXar5v4qK2WrmO9ypXiO6MRvXCybhgjn+I9zMoaP7+oGtIwh0bDJr8L/
VnQGwbQtBa42WV+FSNk5S3ANPehOv9FAHwHEJ3qYBRgkA1+Ygw3+/929vgoRZ2r3BjRDpzP00RL2
qkmyt2OEz4InE6rjNESrXLaVsfzet0JFaLx2pC9VQJKf+sw4AmoxXBJjWfvZtfDroHu5PDRjaw4Y
qFbVidkb1PGWNZC4h7HB5shP8o5C+xk3gxIOkr3hTQWZf9eHzZWnQV8K6E4ZG7WQ0QYbaBVpnHjw
3Hm1xgtGQFMcdxFpqcF9NwJ3GRnWsnv8hwjZze7X/eijif24b6rOzBrCpEmKSX5jEGY1LXa0PItJ
LWJaxMTK/mC9yJi970pc85we/T3N5gdG8YNreEkzJvzQAPZo2sSed04q5o/1/WVLBwoZz/uBwONT
Cc1KLRRdsTGruLvKENx9bX+4s4u+xgyu6tAfJif7yKE4mxA2Bb9kd9zqzLJeSpnqxKyW5sz+nMDP
1fPGg5Z7P8WLrPdAkVIeja41gob9yX0Pda+IAz4vnzMHOILiyuFQbJUAjxT9HP0U3zwR1iumS7Gg
QfuUKDRjaM8V9W6RQBkbxhDVXHgiM3V9UoR5BGlLxONO8SpmxS2LfuY6Q1YZjNVlUr5p+HiW14oU
EmIaNnSmwZds0YcdGdFnArNPd0s4415CMGU9MlwfXRwXm0Hrvzlhj5izBFfcXTHxVM3Yv35uwu2H
p+WvZoxKFq47EIrdJICGlqp4eddqw0DmqiLzgWBVYC5iQxRbp4Bg9Ai1HZvQtVrqeRAxqqJ5Ucpu
nTKj60l3DismTHnNhIzyS8tpxeYTBg2IPc75OwR5fm/kKUU29OrTFjzvx2S15zcJCLvP9qoNd7wd
Mo1Bi4X3lzqVzfGGO1v/1nU3tZTzjwPaKkBN5qO242Bhqic8TgLhwXYHvneMoq9oUWJm1Gl2w9J+
ktE42pNdsZcRA/PQnOd8XVmq/X1fBcCdweJr3Ho7AfBUhqnT+v2JMuoVMhxsyVYQP9xVUmS/FXL+
Kmsh3Oa+FYK7uo3CGM4HVL+qqawZDIHTGvCP0/YJIiqaFOMfZOdp7XjHTW43/396MHm/M717kt+a
6maygS6FM3qCfV1h9J/8lh8AKhbXqNzCaIVELiKWuWBGnJ6O2R+ve5Eh1WDxwLEDAzfqQBwsH3vI
hPp/xRhffSdYTKX0GyzzeQ+plucnJj+fYTPamQKm5jIzV4vqhH4TAJIFExqbzM/mkpOwiOqgeEQy
eQ0PywT8YLmuV6JG0joLubzCgVeiZqZ1bvrfIKy+jfLcC5bg/RDxHqIoa9kkT6AzGC2CckpAcTTY
i2JIBoQupqaecDd9Y1pDB1VW+Xp0V7H05Xpk6c44NGeqlZ94CXSseLmTBw6OrKmtA4a6HGhMHKTc
P2qZ/7ptwECJ28aY7WMEwQgQHOsBngNARV0M9EyvywBLyiC8nm0BgjB1C1UlUrhkMHRLegYD16yL
1FRkvEFzZpTj4Q1Xt6/ELV9eHOISoljPdf53akq7xNVz2YWbROlCmo/th6YIPszZBZL7A7s90UgN
z9862imJeQRxdLNForUelTD2hqQBPdPHuEudG4xTHko69qXiFCF10MOrolvRgN7ybQu9uxbD6/AP
wqai2adCqx+8/xc8gFvUuTwdqJvhuUCYcPXfNFWqfR5mo9fnyq7rkQ30Vn/14OZCFedm00sScjfa
WC6ERI6JNvqbbgq57xAmJtoTNNoZhJX00ltsdV8sv8kLqFeCqMykfRSNN1u8ZpXcK0sp9VU7TYxV
SvpLhNGhZi8W97pui7GZ6Cz6HBnaas71IitgBn5fnwVqmvds6OZ5Rbrc1PTKq20pCa1KQWolA7xl
Cr1MWHcsNRU2ozYUnGE96+yav4py8UmXNTC7lRwSl/gWt/AaMN285VBd8D5mIrNV7nGG8YPidYc1
f6hmcarGfZoecM9xq7Bl6hHGY6aS3NennAXodH41PnDf0gkj2dk1xGbXQbrkKLiW6zyfuvKAzJFn
jL+tN7bTild3P5SwTLo5DQfM52Z4NBsjuxiQWLO3uYULUH8Bsh2d5kf0xszgdard4dJrO+jcT9v0
kviwa2T3+7l/FTL0031ccwzqhpW/7dkMUHezP/EVzGkKDx85+kSfOvs+C/DOcQluRAcF1zQaTLbM
xBdRXonfZ3y/m0bIVNO54z/HrH7FkFSwlz3FQ5fFzPcjTEslcIp40y4O5DrydmolYZhA352WIf2Z
HvybDY+pkprHDUJFh5ej+1yrGffRm0Bh277SLlSSQGEVjrHE/pYK6fuTsfR4otRTEmxMHmxFjH2A
du9RsgMkMmY7eFYZVsFFl/uiQxkM5vkdrX3OBDaETQcZYmnHIl2wFtDfjDflgULTcbA+fsRvTKE1
hy6tR9g4bLVbAClzSFI44NJ8byTgsm+do36+A6UMQBGQ+eHIdt4fBlM12zSA/D3jcIxh2G0DUG3G
BuPbcARdVAVKK3Vw3kpL7jKlfIrhAtoTWYLXTqg6egFHeCxwuU8SFUFEeMMXw+6QoEO8ykiaCWaP
bXIRME8dyrI9c2y+9pwX+QUkw0H7gm540GjH4RTdu1Iiq+qrj7SHdigb1WzNSzVEpGInBfahjkcf
pYpXgF2dAbkSxSkH7AkWJKssmSdCQIxCFiMaC0HocqBirWqtOTiKDnQnDmrzl+Wx8Y67WGySQyDt
UbqA+O9BRT0VtNWoOzegDfMG4JfrmODVlh1WiTcU/joiyBQFm3Urc4yU8EUqM+RGeey+K0679JRK
ZQK3UMQq3wJO8Qj2K+SlvNny9C0uWyEfFFnGeoMrQoniNf3Lt7GnL260fQIUa6FK0E67GQfspLw/
Wy0qNwzMOihsjE4ekOmMOHCn2+8e2z8F5CTkntfBjuwLjY2+EZ8E1dB/dWuRFqJgrM7xj4ipMAPO
N0yALytfKMRAlUkipQcOUjFAOBDipvHGqmtZ0gMRQ7o5mwzusDWhoJCnKY3z2GOs2TDFQz/hZdZn
rna2uNU628ZtmjgYDW2Mq48cQt55Zqg6kn1CIv2tS0NFFsl/j12OI9IxBq7BjKGOJ7R6wtSjTDlb
oRQd0lAjNBE+r2juMmvMWMjLTY/147E3i2CjMvc7c4zY43NSVM8e/2UINfj8LhEgLLgKdlAaZnSD
mTTcDy6UdMPAuXKMfYSBqXJew/bIEcBip3pdmqVEiBgFej8+eHFJeEpSVlXl6YkMjiLpVSD8Dap8
drDd7RbzZGGFXzHyGjWfn8j4m0LGakyLVOc0Tp3YM9mnPY+34K82G2oCnH62mj12xNqnoT1rSsfd
chbDxDFZ05oDYazCpMORfQGbQ/wOhlAV2LnkmBffafuQr16OLVrH6h4Lxo4CnQ2zsvN3VxzufdQz
gpGaXY91UeLIK2Zjc9ltRttEZ+u+Bu0Luc+Ot081DDhg2lARK+HPkzxZwXZPDuO4DnRNYr2HoPNH
rkO0fAFR/UXx9jyJT8yxeINOqzLRqarRdg+FAchVmVzmRvT/ocYFtRCDc1MFY80GlMLY1lpdZAW0
RbxDRnG+TEaeiCUZAfhwMFwjcEDfQMioT0l58qvWw/r+ZuOep/qJOdWUz3ZSuZ+rDnWZ27b9KYEK
TM1/T29l8NLqEq+KaKX8w3J7uEeA1jYvb7BkihGvDRcIfRpErKdr7jHjjXy+WGzM9wUrJLZBnSx9
+LIQ1lw18vgSWTS3OtDWJAk07q2sPQ5zKAcSWZn5NGSTi5vslkJCj/dT1UdsfLebWr1gD7aBHvz2
ZReiFIkNUO0qRfvDQJx8FHYNnrA2zx5729ujTBsE3EEDRUEmMVRm3C8UeByzz1wqCQ8kip6X8nHq
o6Oq+0B1FqK24HSyKt/Cb5cQYvb1WOVkfoGk7STD0XBzwHApU05rsY5pB3Y6KYgCsgagVz305QiJ
3xushSykIYNWcaJjTMApRgln21TJSHU1PFcfJ/sCdXtWk1PvYwIG66L7kZGmysM5F3Q6ukTZmRkS
VnxIklCy5VQeLvTP5l87HtI9tTFGek5Hmd+rIl4aFezBuG+ASF0a9j1NYjRY2WEysUxAs4CZqA/R
FFRuudYjSXT28LydSXsW9pfZ8Jpj15GZyuxtdt96NX+3LEC0JygLxKyTxZuQr9fDez++9ydE7SOA
zuzrVVqatTW789glZ4x5PK/fC1t4Z1M5vI/3rXwJVQ9qjgoQzqbV2CUuRP5Lvg4JlqVFhz8kCOGb
YZzOSNUqAcX3tJD/AMmNTXOwqbg+/N0P+dlkqz1KMmCQRzcbMSE1SFJ7LtbA58sOxWqhHsZA4sa3
kOSwZRIEuCRePwKxaI6iYLx4yn2WZvI1j2pd3TA1fMv17U2j0M3PId8BzsNrKm9VP/AGMRAhSkFg
FdSKsfNdYgouFudcpAFhyFc1I4d2kGJwPCyhbNhkbeOQAE3IBVWEEiOH+O85dCNFMzujjGHGcpat
dYCD4MftK9JelLKxtQQ+maasTQxyJLQx5rNAetJHrqq6xaaabGTxd8flM1E8keD0FOqk4I/CGffO
cciBxYP6imVfR0xngkn1cGAxrh1foNF1u4vvEQXp29EHXSg9/DokO5QmMFWsthI26cRH0lhPuXx+
JjIZOBUN/kXxawd8X4FIoJfxXqsD9Npw4f+83J3WwmtTFlKNH5s5ickqI96mLEI2gJMSZo+R+9wv
rYa4ykHXEnRdlD9c+jKhRa4m4wzRlNSDRFNuOc/f1UKWywSlz95OQlDC+MirJXkYVAyzg+FbIBvD
91J8GoOnQql5FkYAfTRnroPQQCgVhF+w+Ywo9a1aZ18C4M6KEAdXoTjit5oUY4f0EWetCwcgnyMj
4dJB+TOT6G0oquoD4C+2TNj/crxSufsmllJsFuNo6hPSGJy+ZzS2Tp3q+2pPqFsxAHq2xQjpR8Zh
8QDv76Pu00da4cefsfmta5huL5Pb6tWWVGXgwMnjhUPDhpklzMOtJsG+bzUYhYkzTuu65gDPKm7k
oemFFZyBtmtu1IqrJNdRRspHufF6WXDADdtE8a6oZrHD/wRn+SG1twtKKQ0j3pS0yfDDwWk9Qfui
ZmYvOpjhGQ9/gKnxA/y2fz9lKW1XnHQdVodN4cqqf5f+Gb2aibySA8BJ49YOecn6iOAQb+IhOtZ5
xr6XP6e0SiCuKZt0LJTJ4vTabUISaqjQhsVZmw/9nQiBlirblHKAEBmIj5bf5KK3aXf58krjTS25
y2cDg8HeFm3ahQXQPir7lWOFG6aNrUCsVCTrBxYiLHd5aCqzncXgjDnKnANNc9/DuifNu0Nnt4Yb
zvFGEA3V40CWrEtv3CiUJnKT4EtgywYLJkBwMvmLfKJG/7ej30Cqo4Yk82zGSf/iGBcetI/l3Mw6
3z0R1JjpQtaik/0qPvgFNTQO9K+/uwRrbmvX/B74uDyquQOjyV+5LS1Xf5/T4XEAdLuEzm5NLTHJ
HFmT185+b1Icue3rsz9dg9VXq7cic6+XHYAnSfCuAldtK+lp+RJo2NJg83Gk2zzCOrKC1xRcIZnn
Pfst+qL7zobALgym6nJcOz6vVgtorzbC2pGDr9CEvYN98hy5p1OQoJSzXu4hq/jmDrI1sFFtPHpO
e11sYC4EsUuAg0igT5MzHUgVHtCF2wp3FGv7yYyeQEoFsz2/mvBLEc4ol0R9NNpXysFT8TtWluvE
CaXvUMCZoqKGFmL3u8Zelhgrir4JHt4jac8dRVzRnEMztOQ0RdhD7VRDUCi2qd2qk/u6vmDCJarv
j9QlxvqYx0vJvEEZ3ju3rHOT2K3qHCtuA7bWmGJJooMzFEdg+k5t3u+umnC5il1BDYXcUKSJoOwC
lNKmIYPk0hkBi/HQgZ5CnsU8ZtcssP8b25RLiopMqYOTW4QRkG63HpM6DJJd9vLbyyd77C1zb68P
WQBn+QHy3aAyVr9e9kqltLKkR0/RhEU1pNjzc5FC39GoKXxcmps0loaT5Kq+ovMGRQytd4wQenJL
gDJpPu9sea9fx3y+QQuckQ5OYEXmtQE9DPQZVCTTyUGpkMffJMKilln7SF/RdbBdRFAZbVT+8th5
KJL6tL29y18ddixmn9alo2xZ4CTXVDHkO5/lkIXBHcihQ3EBvAdTo6mxJO4OeXYXUmOB3YEqSJcW
hrvax9uPTyKB9aj6P1WgyNe5DtGluHGm0iEbWuvM16VFyksypusjB1StMVEzrl7C81Op2Jd54prx
98t7IowBfz/OklgihB4tV0IBmwoQFeQiXTxRx8PkUayGGJTQXzmwZCCkhnoFgoTiSnd1syfKlnuk
6oR4tV0iA8bGd8a0dIhrYAmib/UahSMOX/Np7d9NUoKT25c2+Rrt35yVZvpvDIGXEtiSYnScK/t1
fnca5xg9x7kaPxFsI6c+FNJNuKwOMIVBwE6SFT+pCKK86c3PofZyBDWI7Jkuook6C3lQqk7vhDFg
VAps7bPdT2ko2hNtu1kjZq/9ekREoLPXNgM7H+nYpefp3vmxkffdvUPPdJGTKv0c0GBmpQHt+KLo
7rPMnpx6Rplt6Cp+KonOqoz5MSg0OMzBuriLU+b76uhnoqzlRJwlO+QgY/pw4QldvIz2MxsT/xj+
mq6qqzjaCsglwyBistIaJni4sJtr8pWOXee73iozgC2LcSHbpyvWwjy7euPWqboD2DM/2Dko6b1a
qPXzNfa9DM2otJIXYGbUhg7r2NER/33JD0yY8wu22yvXpq8eHjeiBk4GNm4r5A9CgS6VPFgrA7qi
D1UgD/bmGF9hOmFPuOZuLqBOp4zauZ/95Yrz/GBIdefTlnyLfa+DihzMHtOGAqlbmc4mejTUrejn
dZuDxewcKbm+aEaOyohacrQpqqtnQW9/dFaNNnzomjEgD+2XyavLhe3iq2lpZ7z/GIkS0fW5Fw2A
rHIDB1kH/OM9pChOspvQCQCvKXpH+UASTNXKGjSoR22bCpIVoRCQRJrAl0U3LIlR996xksBd/2dT
ha+Tx1smQ8Dm7ix8bNuzjromY0x8pNE1iq2raKKnoC7w0/3j/p7PxNX2P4LcxsxZ+ToOYv7eOoty
ICnwxxYMYjaaa176EhsimVjxEjWzlJop8uRmmJ5tt6iyUUyUbdDlgQpg1bNUNioGdz5zidbcOBFG
3GYANrz6b2qAZiZ7ChiZ+Rw6hMOp6Cf+3/gDWOtYi2pXD4ZsCAeGW2EWBcntjcFNikFWGnz/yG+h
IIb0Y0gQqw/Cuab+aCmUTY9d3nOPlFkKlZgzKMn+LZTfAwBawFhQt2e4o7SivUapBSEuzJFr5dGJ
sLBWCV3miP/uVeIqz7V7BRhp7ZsK38p8MSDoaHaGFVpElsRwOilynGeWmSf1rEjdxoQHIxMhSIGH
u68UOrQc9RW3+mkMzxJYTUGGXfBZY7RgdRIiyyr/VhoPjFD6A8IbFKiB0oudTO1Uzro2AhPWbgoO
cYg8Ttv8dEHCTzG48nouyhN1Q3pOLFRQJFQMj+XlXOONWfQ0yQDl4nSAO5YRJ4AzO/gHFObfIU/r
VxvoqcxHklfq3HPT6vtsuUnANF60zJLY5r53WJ1OLC9NdzW/U6pkX6/el/5JaWkxMXMQy4b+FMs3
18cGWnsxJmsk2YGFqcACyZA85KO8d7RfWTDbVxk4olqFEvCHRCCYp66/XzyR3OnfitRYeMMH8AVr
OwXQUgymwnyRsJgILumnx9SY0yAG/DSPtwcy15zFCmOS0P608PKhA8CR5GrTyeFN6/cCJxMhsi35
cdWJQIDrgsNYd56kLmMnLpcYTN6p5R3xS/12zbf2zh1ek38fSMasLTczTT9oUBgVbByV835omH88
otvjKE0jdZecsfu/+DqYSV3PijNtm4HCsik5zgJmXgTPVBzZk3BGNEzk0K349F1EOFOg6Zyy4hRL
RXlcpPXWFe+fBWCNeqPfty31tlHT+w85i62u/NniUWphhYCBLqKfKvMtrq4PG9GKlkvq0yLPJ5oJ
qL0P3teWpg9kW5J0j3aJgylijRBCx6CwtUrSKmJEsYon3A+0NRvNLCnuBFiIcpdvM9JdtYEAT5wE
HiInkmwI6Xldv2/7WYvbMNu73OE5QDdYQJi13SKvMlhdxPUeTjDj4OQ8irQeQEIUoHrCia9w5oYZ
PhXkAXHWCRe6O9MQ9lXH76+SNYf+bOxRU6UAPeNl+aUimseBCBsWh8nBk6ENqYJkdM2a4+OfaRCj
+QE+ByA6tHKBaXOyyzZZPvI6NVKorw08wGmiwzC7uMnHGnZP9UMZbCKUMha4zmN/z1kQeO5mNVbH
fAR4xARD6MWIPO7oNvE9YFCsfuRFUK3e8+wGh7M8MlBxoRiIY89OZC23ITCcdcu2PF5xfZoSlvUV
LiThIZXhL/HT1rDFihWU9Q5qW0Ps6Lnrg2d2kT/nZRJ7Ux4VKUPVM+11C8MZvIxJmDlwyhN7P2Js
WocnZ4QQD4/BN0r4w3f6iK1LV8LMjc4HQ+YpLr83d7VW77h2usP0VyL8Zu0heHyc5U0m2ZVfbhSP
N809E4ZUHNyUkeq/4eiPubwsr5qrPw3ofnnT2YMB2eLtNEy9q7ZZGFupbQkYxpQ/ybVUc15ym36T
shXrYXyC8GoRchInUjnxhIP7qSH1IUNnFStAVf8YtIxpx/BzCi8+UJt23Ns9BhhWnz8QNNYUte1B
bsVC1uwsfzEKSaIpy3mFwgzkqTTyLBIbQp8L/dxoYUrobUmxRwyr6bYLezo0yFKGRkNsP52r9VQp
8h0co/EUvd209h5PGXvuLMAPR8V5vlH0y4PCSYYDwwuazJs7jqcehIwbj2Vq/6JbXwofCSpA9y+y
fCUjtD5mdzJ3Lh89RtViIgMv+w96f1AdQKjWe/W5eCjm1JNwlHVQopimF2am+AIXBcF7csyFPvaQ
n2uYA64sPa1D4MlN5gL4WpTv8B0CxM+ksc+6HeeuLLj0rkiM4F4QKizsHgEC2KN7CO0SqoHtYo2h
NBLUCsFpxikc01/Ndaa05luE7hJISlrX3evPuLjCmakSrXjCcwMjVY5R/2NDhDylg/uB9cLjUNaG
/is2exphw93RukOxb7TBwQsfvR08bfsiJnK6KPIgQLaLxn8ryBlxC2REw+dNiAu3b/GANS967Yu9
AarvLMg4NMcU6jOmHzP36/6WBOWo6TNpxB76OfQxWIbji3Ui3GqlYdUUiU0aq6nZbOzsblE25Vcs
ECiF/Z1drXctD+vsSg08ow/gy82oXtJ+TVNygeMJ00ssyagUHuMDGYMWLawBhrN/IuROmEdEX7J4
2dsLMpGK84ECWUnTgHLeDKcvAy8p7wE7bEMxsW/rWDRrQ8t691HAxwjH4XLq55rY1Ae0zCHFnzb4
cVke6OS620CY5jpm5ari/UOVgpRgWc2NbIMaq6Ydg+jOrgPKl4ralugUwUxzDQKISOSSzwroTwTw
qTMwEnnRXqJUhmLGfcZf2ZwoBaXD3FneopF+RqbyUYSmWaIFkIpFbS1ocDCccq1Uw/ychOHNODSB
2qJs9L7FmDD1zag4l3NY8586Rzy52eHSw1mse7APxDSOouyWXVQj+8ZFd1mc3unHbzZUTtXZySZN
SN+mKRz9KFBLi/6nkOr2hUmLtDG1gZ2mcw3l7FwzcBEpRpyMd4XJYT/UBjRmptL8luXPNP1DIEVj
Ey55aGToBRVtOPJpOrbU/RjMKgfTpCwfzk/y5j9udQX/eeK0+exOHny0R6x783lQ8+Uvd5C4YpPv
bBOd9/SaRBi0YNTP3seEzxrlRMemoi3PVNq1ORUB7NlMvG1SGr/KxLecKrLD3GlQz42IEXS/1CDc
WN2sAG86dhH+hwadMx3wIpbMSTpWdN5poPulwn0RJENBxJtxbr7D7Jm0RuezEtSHD1CY2o13PCQk
A/ApEHsApW/fX2kIMP0sPUOUPGNgbApepeFkv+qiKwLv6Ou/DCSQk389ejO/fMoHfEyXtfuzvBR5
QqdfUdkpEEM3TFQh/qkPg9zYOUytMWge7X1NIJzzTrbXqmy0LIOVY0wO2lAgdjrZcPbxcKlYtnVK
VPFxUoIr8yja+3WbZzhZB1ye7TPaxM2exNuoblV6xoYXheNArCTfH3grWWNFgXkffQMVdHYcNuh5
9IXzht/lJLQXZlPfs99NWNlzB1EehXGQqiDT5FATZNBJzDByuh72pF+cKI8h8FYbH9g116/+uh0X
wCFNANHbFRnCq127bEdUz9u+mbu9Ns9r9tqptVDg7WzuvajqIvmCvwOLir5Agehw26GJBOpW+jKC
lfDpiPcXm7hqJSJSIbUqVJsugRqyfn9dOrBlh+V5mpc085mHKHk2bKJFuDB9gPgrUajZy+LNNqIa
kFSJ0bZ4s39mp0k3Sb4TQh0EhOgdBiud5HJcglnh+n1roJIV0gtDqeAPZvihTG1dhyehaoKtseMm
xBB0sosgdRK0PSckXGSwxEKeYZgmv7v/fumlLvbPJBegzh80vpjUuWiLAojeOXBdIU3FhqIoOnfh
8YbD+fgt/AaXZmdJbeGhMHm5IIe1oAm/sv29rVOTvyKr/pAIR0uO9fbfhyFKr+nswO4plzlbgjM7
Vd1Emi2KL4FKZXcfMPuydDNW8ZZ4SYlHkxERwKrbPNdVN5Y5hcVTPh2Rm7YoGT7wx0Qh7Wtd9vW+
b0liI7BFcicHp3mBP5wDM4QqMLLgpqjc246QJOLKiYrALMjnMEilN+Y603+lnDGCmA+jRwnwmeNZ
wA6Lw7rgEKx+rtzRppMz9wyqn4TLceCRNfpy6Jge5fP096+oHLEFh0u90E/MeIExCc6W7lkrPC7z
bPA4HfzyaH/tK2RFq3jcqKeLmRqOQUdFFEkKsUPnNg0oT7xbCZuqcI6uyygTl8kFeysU6IfwsK2e
r26OIkocmnGr+WvqLT8WYCSDnMuEANVed87pAD/FnndP3WjXfYwSWAdZpR+TycyHd4T6jT8HDnZS
3BKGocphWp2njXjQVUJMFUDV39Cge/nBPn1G/ikoRcaTGYyyvbzmkruG3vHLYd7+B7o0Tw1/241k
mAYxuo2JaKoMyneGY4Vsx1e4wFOXRXzMK3jyGgloUx8hQA9S96pDWaQ7nIWqalOJ7WgwKQsrFHzf
eHScq4J8GfggY3goqaJKUWvF3NBVJGhMkBm6KSleloMvhB0hhjWE/tAVaL/91JuDRFkjYSUzmVZc
SX1V2YlZ6ngdMpEG+7c7uvzoUOWAyNYTpmyivM8ojDHrik/FoOft5EP/nJY5ByZTVxJbmGF1xtFX
5Yadj7bp9/RAPAXmWMj/LA7hJ9bA7HNE4hJ/FxWCv2cx3tD974jKINDJw9CHMNyg8mJZXxNIg3ei
lj39rvreUU9QFYYvKXZhgxcUV6QQ1Gyo+wTTpj1LE3+S3ManGOBt0ok2T8NSB5LV0YSNC219yquZ
+SJsIOBmy3SY+YpHJNfMthdExQIFxI0Aniltx10cwStEO87J5dBiF5vQWNnWNDxeU3yQ6v85MWsk
CvBKS1xu3/E1/z2NWB8jBJhoVYZXHBiPRCyohdx7SEz5WjoZRnR95fZHj9/1wvvgWkvjKi66YjMk
9nvWk8Af4QKucUtZX2cHBmsfgjfNeTQAtVyEpSUVUd73g6loldxqzyVXBffVWGTF7kpB8DcGQ4Nx
S/sUXmRZlwj50ZV8OejhotzRmF8MzpLbPrsfi7bwINAB5Nb7dKUFhCbF18zEixwG+YmnBFjR9r+5
B7rAKGGPbH6b3BAWCJeqasX7PLxmtIGPlvfXsth1XsiQQ6zAvusIRFw4irENzyNIJlHE7UEZnvvT
piGPXpKacBFsgM3QKLwLlD5iLyvcPFicvFVzaH0/5MEs90rpJyjqEwGAXGUFs9doYSGQvurLH+e+
J7S7Fexvhwmfef8+fTTrw/0vCe7OPiGuFYFMv4p2vwXYbT3EIoM5hcFe9bRjYSWHkfJK/OD12bff
LqLc9tT0V6kZ0uIbxwcchydV+U3+28pzZLou6qOlxHLxfL9RYHCSf2dBmglMrUutnXqxVHarMRr5
fBalK0Z7MJCtvMLhx8O7fr/702mzaEGHd6YKnMzKhY1htKkXwCUJJgXKbdcKZ6UjJ67bLtel/Qhl
Mn8hllvO6Daqutfe3RajGtvrr2ivCEyI4HjRboMZe40sfUG064BiVufojntZokWFcXst0+w1H+SK
B1XmbBsHXxYznHWPqOppPshk65N+F1q29fwiuU3jXa1KB4LSRB+fJiDZ7wKK3c8u2A5eEDK1S0jV
WQkpc0qbBL1xvsobFxuCEQEhNM8XKexbM4UMnnPyMTsiKh3yDiTa11VouecF6DzKq79jGd7XQWcM
ETbUgMqtTYQJ8GRe53Meu4Drhp7T33/Nw+XvnSir3m+emM0fVCuSZg89DBwo1gJWii9M2OWx5+gA
5HhaLhL0VwWicAG1HGM/R6/hme26PzF6p1sqAf/6cwh7TzAfGRMev00CJAcYWe3sGFW5F4jVy8U/
5QVd83Oxe3SUuBTzzorXKFQi+Xkwm6toJozlbuSn6opUb6HM2mz1BKnXzcilbHebrQtwhXTHbgtQ
jWHvMKmaZplc6rPo8sRKQrY9Nj0txUfC0TXADgcPktO9KXvoHtvHykjMXhSp5Xzld6ktxPfO2ugn
QG2mnY9hbq7WRopexID44iwh/QZPv+CoflmXmNAQrf22H8daSVs7PquNkyfsP8yMZtI1ouzQ7rqI
40R8I4hZi2b3tzaYZ2DXGvgLxYw4oLmQZSBdmzHzya9xb08usV3dCILBytvnCPJ0CyvvzdbfqTZJ
6LFxgj6Ry0cCwHjAjU61muIEOio6CF1QclCa+DN1JncU5OgQMrsJdddS4PriclpQJsmJc/4zjcoC
S5SFHsNPE42/AtERmtdvBDIMVL7wxO5AEpilFOBb6lTolxtq3zHyqte6Luxvt2UC2YzV75dWXpcv
HE7RRHcgkK70AcijA0R7sMyHwi0OhbgjfH7FNL3o8fqX/AxqD50BUxlju47sSKaRHqWvLkvjqbQ6
Tukc9fPiXS7R2Xin2MITmKKw+WPawCImVy3iyBEAreH3jnbuLe3A9MIhRx67/IBXL7xc7FzWhE4/
EqvTkBT6WHQJTzNj4KhlyLACYdv6Vbo+7pweCvR3DxLtIk7nKapyb7uzElB26nua0wGJT/eYtGWf
9kKGyiLok1alf0RFv4OEcXalvCAhiPt1Kfbh8MWzkpdtXYRrfdYCViJAyqJQ+Mi9ox481G0bscvK
AqRCFLKZcDsMUUApds4T2341SdPyYv20zUOssogu3ghNaoq51OqbvmroGmx5ERKNtxfHaSK7/bnH
U3TMBl5pEGNbbvn0mtIPuswQfTQ7vdZWw8Y7s2g19yJ0BhedDcfhVvMJRHdVht5H6LchdsHNmVNY
PIaehjbd2ZeYIeACOeTIeALD6tI7gyX5W5P3HD8DHASl4nPKiBPKmBiFjOOtNKdWLNogYtVdaJaH
7a+uEq/YbR04Jo7RPndEEne/upVAW64QwC25eoqK13kWG7KRPXtsUP2N579r/A9clSzkGLYuLIru
lrgzXBCnMrMHYd6f+oCi0F4Y156pH1OtVwxzda66+XYkp6HC/2whZaZCnmjD7igc211mi+Xr9X6T
qxq9K/NQPNZRAE12vNyJl6JEN5k/+t7oyzzsQC5nGzjv3H4ArXE3cKiJoViFjt24NfZSV+E2qOuA
c0+J46UHC71wiDF+rn0fP7oF9nYBTVE/38i9gjZ1ZpzqqIdWXOLeqVCZWrFOg095j2KJHQvCl5V/
HxizzFZD0h9zk1gt9UTeVI03cs6rucJyRFtBcwZ2ktuGv1oLWTmtLzUy6GdD/iELauGg2/LTybcW
JIwxTuHBp8vAffC6PmvYn2cdVC+WLQQpjta/OYi1Hg5K+pL0/Niz2AHKqD16XUsre9/WHL6kECD3
4qnvS852hX0VGh3HBKNtlgOmKvG879zPy1lVC6I1vNAS4AKEaS8f2ztFerdmwpxNLTDTJ7rsUVfs
PSUnXzM+9yhu26vBUw4IrBkla/zIiaPTWadGMuWgeTh2FuqH5mVpNgJWdDbDCqP1YPUFeMloF5ed
McomKP9CYsqrLJxpi64/XEq+2aC7FRbWeOXAwS/wOET6t12RT67Ll7gtMg1zj8hsjq2Jr1bzypFq
PjTNyFaZdX6WG8oVX39sXrWS+ve9vw0ik3BWcLbHj3UYp4NRwTUbKeVAi9WLy8B85TUMy/NVSaWp
utRnQwjU0vWC0SY0uBe5BirAQL8e1isMgkTJ8qwr455Ro36/Acydlnj6prFyfzwQ7XsfJsb8uDpq
yfYiaohe+K0U6YjUmuqFOiQdghbTbP4nD0WYHiCh+nl4S+l8qCeaLD4EMLvnsRL5aCQr7shXZzZl
nVx7P6XxM5pQ1LGzT/dmKtbut0JrsgUQyCrX2CVlcOIFxQ99eAi9fJmTv782yDn7K0mKfi+y0r4z
Rt3q5TBuSfXjC76oETHFpvfQFZKcGlPMCpv7h2odx+xsrEFZ7H0ckHENxnAGGmtY1QQMUOkc71U/
9dE/ccb6RtOgvZHKFv6uFLXnYIgeUOpwHZRy0pMMCcLws0bGgKxtgNJf89fztNNISwJU9QsXpp41
KLSDGd9/Mh58TGz8Nl/7m5NAImhcC5XYAEYySoe5pi4oRB7n5EEsVWQqroFMMSqOI21HTqkhoLzn
bv/CYadejQVlwpF5xYZXoR21wceYW+Kh7FL/2R3hSo808WA5B0CZjvS9eYVtUrLKibC70fUbCsJq
Bf6po2+SMF22rKvr54a7M8ig17mj7r1yfgQaWSCVdXnisQ0mkO41muW/HGiHfSQo5fVxIZ1GssVq
JLMRowphsaiBMblWrQS9F/Ul8493nx9RttDvS33d9IY7dc3wwKQvjFSgfAyx38n/q9wtAZhI6s0h
2zaXNY9KH0Ye4z//JhOR441M/hxiNa71LAzaMXl5V6Q0X03LoMCsNjU13TFdUililyzFAyy86NnZ
zP1UGyRrGD0yjShsOns7iG3z7+Kg6VKKF6q03XkPh3ikJwYwvR20hYXaKmIlU8rWVwEzMZtGyRAi
aPeTRVi5wLPkgdRgvdcAGwFrEXModxzvdO9XCSVO5mPqmBAJYRbOi800X87R6jG9W69wp7kOVMwg
y88Y6q/9PautpcJROW7B07GwGGgc8InFOI8u6wV36/4+WBTCy1XgwXuQVBTztqc5P6ldHqPJja9e
KFCo2gc+iVbA5ee8QTmugEAGqQaL9Lf36U26NrNR57vxagMf2x6DuUgLl+4YJvpFkbLuuhcPIqw9
1dnZqFiyTnCcp8HQI0Ws7r2UzURpxgQNWBZyZNQ02CRbqp3qDV2fEmcZtwchZg6baQE/XDvyGS4w
eTjDXRJepWZsW5rvo4UuDAHlaYM/43297gXraDSOJ2se074aPgD1ynHVOeOIAF8UmJRSHi/Hp1gP
QHnMg7T7GRV6/cnHKLaQnV+lfZfVwT1C8r3rnTHuNuUt0RQnqZuEYscL062YDRYbOSTyvN0OBr9s
loeQ7/Y51bOPejy8IfZAP62yg/GFHh6MIl+tXOvFkUpRzZEqaXVHp7ch0ZAs9EtELDPwlpM/a49I
fKSEpmwfj6UliuxvUpDVjj5p2McacIkO3HZ7tBCyuvP+vf4Lceh5hdA5u3JUmyhcAFf4ONZOfU+g
Gh2Mkl5/bf0QwMjJZPldE/gztZRCgWyt/qOEa4rOfxthI8+5KO7d3rdMV2PdNnuRVpQ+S9J1dumx
q2tbQ4W8yPk3sdcvjxcpEU5gaVTb1/tHPC6+89kVIuLbb9htIX6iY3pewhoqc/947i3grN7DRPrr
lKtcOzao2NW9RJuGsXzPnvoqy23D26zwwv9OyA8KA+HTdCPJtH7lRRyE6Ck9JpWt5Sz2Dnkht6A4
TiXg0C2i2kNnjBtmpQmDFTYYSHmDE7HAm1rXYTyC5o6qVK/eRFGNg0Zhy31uo2OtpwphGKioiZ86
7UJEGEZx0nMs3Jl7Jvjc0dpsMl5v3tbvWJscnJGZo3uT9eDOfTfLOxosHiocB/eDcR7qNhgWsueM
8OE+kSET++fcMZ00IxHTehqDfyFTBUEirocROUwaPBo7YXFcsr6GuakGInU4h53Dsd/Gbm9UR4Pz
aH34exq17pSmykO6c8/l5cQLgdHowhiG140m1YObwgwb3PQeN6c4kLRKHeSoReRGtJIQrNG8c/Zp
QgeOzADHf3ir2CIOuMsWiZXKQesCznX4sRaQV1vZFFvjCSTCRp+LylbLuXomAeKx7b+k/N58YpLL
ShOk/tiiksSNG+7a3B0ylDW3b9XsgD1AzWrDKAYMT3Qro0cTv0A/MQ7nTi05B444GacqFeedGQtB
pSaf5MeJcCyTSMRQLDfVpLZvVduJDbk5308xUAl9vDI2uV0h1zo8YdBtbn8FuuDYcxf2qHAvETgf
N3tPlLuiM87lr79sAZzEjYuIzYvA1uUT55eysK1NgTGL0f7qQxnu+W24K9S6+2t1/2szVUeqDm+d
EjMmy1GswYPnc/nxBYvNutTgzHgxbAuTq6svopAIc9WGrD+/kgl1O2fe+JqMshdty4dlsKYSG+E8
DG1EP+lo/hRQLV9tv0vvTRlLDeWAP2J5bs+f2Sa1pg6S6wrlBNQ83RMB0TsE+e24SK8h+EVT9nR8
2Ogf086rLqAFPyDJb/xY6pOgw8uvbB29/lY7fXpQFcZb1elvAP/zaem/5wia/KFJK5+kOXMMtj25
+KpYfzjmH8LHMmJwMGOKBVqWIUmUbzs/3VfKjk5XqFlSYZD9y7yWXhF/rk4ZZJesvtDk5vzT3uWB
G9xFFxU7psT0RapE4eeYbzUyzqEFx5h0FKWDWUPqC/qWPahE6QYnKtY3DRaYgi+m3l35X3w+sFVN
PAYCmUkxyab0yvhjt3weln0hrY2lEDL91SOeKIi9C4Xf6CfDYE9BcJPMvF62PYctSD/1XCz0Vv3N
dCT2aK9/o5rEK/s4qCZx9y4BeWQmY5WDF6CPwyuaa1+Y/cQgFkw65GZxTnHNSc6zB2sNWYTOPInE
lMHyjU7EBDB+cQwm9rYGtTzEjNG3AYtIqwgSf+bnYTddfR0Ecms8Xl3fN441x5bX2qdy26aAcks6
QCDXIyw4lIGDILvlShWOnWYUQyn6wG2JxHTo2tc0jQudv92zUFluTFO+3KThi7xFY7Hny8oJBwor
TveWn/2KEy3qa4Xabic1ict/m+NDZRXHq1u6/tjiOovK8q7G1s+jmYDuK92jrj45PfMJGd9wPHZO
yBfe0pjk5u5/u/PBZxu4RM7B4IpW9k+p+YVpggoirIRw7ZtiAhDOj6p01DlIvNgkC9Kj14C78ETn
VwjvHF4w85/0qsWZJlISWFS6nbAIKl2GZ3YKnbWQ7P8oXjThGnns+akqpfhHoTxMQJ9qUPPLD5x8
4WcA5O5yuCyRtyIA2tl70AZV6yfYDDsXPOIxRgJyY6UM6XWY17FwZO/Oo+JVm5x8NVCWFd2hSxsU
A1/J11T02pu2KyPVYf8aUwHYxvWlUG36MLqUSXZ9HQbCETyT1D39xKx7JE8YnuZ8zSecYB49KAlr
nCyIQVYXt3skmXFVe+rjvbczG2A72ZfV2t7gpql1ZoUetwU/tM6CA1WXKkZlQlztHyqOdTVSyPCR
AmrJ5xTVypiSWdDkhVGWr59UbRVfqiA8J4GcHqgxZ3TOP+AtX5+4W0n8rabyGkbu3zalSG4ARKqg
iouDPlRSxNyWKD5W8UtHKqN1XcfN0gpVDlqa75rd4RvHCeMhEyhR/9YQMJkoifE41+i1m/BRwxSX
MBNkXeSUV9ju1D5klGjP32qIHkPQ9yMmVHUjP/wSJqoXZM2AtNm6OtOfnYufH4xH9gjVibyJvl4+
Aua1fGm2xwlWSMc0F2NwHId49ZRhsKixfOrvSz1zSNMgS44sgyLbWxRD8ViJdKNzmlMCVHqOgF0X
JcRAadU75PEtln+k3FJC1BYVQ8MQvMHScGaehxghDL4x4i/QqSB4T+JYXBOjxGzU1U2sWdId713j
faz0XzyFJFmzRk8/f1unuaqaCixrfo7ocw+K/D0/DdsSfAguUsXD2/AvtBrmUZcPFtxxb6/gQo3e
aSR21zDOR+JrmIIV2PwSV0qpGWLKc1DaKGxMGO1sZ76FwxuoHm/9H9HH6SIA95R+XJ16AaM0kiIS
h3VCvbyNWEZTvqmPClJCCkAbMQwBayAc1SfInJzf+LQI/cA51a/M9I0v2NcF/iVLhHaZmqp511g1
7+moNTwTHZ/XF/rqxOym9C1Hdgo1EYCf7PyYruSXc05c8AY80cLF+X4d82ByXPNRaapnB97ENCz7
MCxt2tGtW8tdfOl3nbxDmqHy+ioHrY0Fspsn5hU1NZKaNKRePP/n5t3gjL5Y2iB7BuHo3Yh8n3O0
zQWzeZZ1Kug1W3Fd1HKMEEmswyjry6UW4x1uEG90H27Z4x8n5LKQr7UxUEwmCZ3SU+FUNxF9YGQ4
u+ndcbNQP9QBC1jSsYBKy2MExgS1oKY6WedGUA4fWEpsYkSW7/QXepJkAZP4voMiiwlzkZu/4FCp
lSWg6suJ9Txmh3yWksieG9jDoqZeTV8nRJGVZERpMDv1eYjMdsREusA4zi1j+RBnKXlfsFOWY0pz
kIlJIcELllHhUmJGG/Tf5bX45AR59l1Wh/dRxmArgWB/ZxjZsLtjUw9XcoRkLe9vGqwaKsiUPAMJ
OumI6KbCsnqDP9Y64w8eKdW/Z0mlmgrGQ4nm1Ov+2Ti1GorItYMl6mT8PhBi/xMBVoWSxkkKBfyW
12r1ZkE+wZi0f6pmxIaEHMdzPmCARkn9bj1j3FxHHF5PL/iGGnKsyfsoOXZTGySX6+0I27HMHLI2
Eyr4crgcZFPX08XW3t/tz5O8cw7ENTPwtS5pQfhDRvtsiWiqMW6iVjh2bDeRd+TC6JDGHvXpnWBK
rP9UPQGERvJfjlG8DbWGMJyzGfIwuSuODmqmMY4G8F59WfLBiQ/FvMXn/Da8Lz7HGcKG21Jd//gl
8sIX9YKp1rUtDx8eEnIO3KTo8I8rR5AJ/GhRp2ibSsSr2nbwpBlQmLLnEhj5Osmr9OCiqveKZpIe
hm3THz4yLHE77+U40Cuz/g2A2M6dsr2ePusAEgZTwHrMC6/8kS3EeQi8Xyvh54ElW/qmS6495KfC
s/70+qoANT6aWMG/relzY8ynOUv2r4jPur/eMYY+p6hcn1GECxPnVy2rPzAR1NXlAKJHZGeXp/w1
SyQqnCTMRbGKJreu17R7DD/KvOpQ3ALrpx4YhvSJ0oMadESMIhsT46ceq7tjZ81O7ufps00KmB89
TMA1cwfMTiBVSzOLVz7Ia46t6gSI+JfF4ux1NEa8HrOVRitvnMaT5dO+Q43ZkX2KRySd+DvJ6FyG
h/SoS1BicHSU1d4XZrnb0qtQGnbwqOLTUoiWR+CtZEQ4/6W7sth3b572SSCnlg14jiJquoWtvfhN
3WTki+jcVhBtm4U0ucrvmZYcVRbs3MbkI1FdS9n4sINEQ+MfzvKByt6KSdegUo7spEgOS5pk16qK
pnqcAQ6oh179BkxNYrV+hQ2BtAP6FBRHAaUHrxXCCmOqlRfl4Hj52aeEGegJWdvp3Hjv67VWEkBt
8rPh4VA0FmV8VTbivMllDa+XEJ6RhBQdba3zu5uPJN7BRniRQLlwzn089hsOjhcwHbvWDyIwAyxa
K98HzlGSgwXQivRoi7ISHVdQsx9/J60W2zlWfq4eDKbuwMBz/Pg8udGS+O+CrbIRFn0scNm4ZgIp
5u63s85R9mjMeulclT6Z7QapJSJ9KdyeKRZJov3cAbabIupB7O+skcXHavyT7upVDObw6KQJKK/0
TBg5NdllnVlmc7zvZV/gFI0hDpTFq65lPwtSZjI/iyWDv1Cy+Okw5Tw5YHnF37ujm2jxLDgJaHiK
YgafohrM4bbPUvApX2OO+C4lE2g5qQPy+y0xMD1d4pIryEn7ndYiil0SI7HM2R52YZZPcUiOEWIJ
aBZ1fpDIuxbOmX/JjD2lWJXqiSvwaojRT+zeXBtSWVPinKOjujNSCqBxR4aFooysWV/5l7D8KWh9
FaDV6W+c45H1CF5Msj17KUcvURynTV53TwqGjuAYJnDjhkjv+j0PsbgtxuOps81TZARP4gXjUtkU
O1tLH9hr11vIUabCzMACpmuEn8OmIzWgDGp5nTqg/7nDTbwBoHpUI2yBbyI4UT8h3PxSmhwk4O9u
hMZYwHyW/hRuy6/aq3TgFvdB7/85qzXT54onWgTWizProkt5wOCHn6regJHuk/j8OKBJJJjDs24K
PHgXcD98mprW+35X43bpI+ft/ELhYRyCdbCNBle42lrwLTAqEGu0D8dZ4TTUrraUrNa+GWuVO+e+
XKZUYg0VkBKwEaYOFbmaKRgf+ABjysknAxC4ClhT+KvxxFaxiyu4+6lkSdxCTzaQklVyFhQvvClV
dr557C7gbato3UEyIG++H8KAVXfm4MDMTMiSBpe79MPEIpMcAvZYpAMNhVdYySNFT+VUC50IBXez
KLkcUDsLtDO0t3DXpfgTdtsYwt/SCdavvheBSg0vd6BbPcKs15orB7/h/Tu7hfFSxkHI2xdu/Yhg
YeBaiDtnFjy3Tw8u6P9srpPcFUJ0G7IYv4OzKYuIhelCkJeIbDwiaqwOrWzOdUnTIL8s+buxvKRo
s84t9tvX0H74dw0k7yNVe6hDuTGCpmzCSWELIni96tcYL3cJ3ixpA7IFv0jO0f/ipHyOd2yTdQ+b
PK/1A7k48F3j5MCiIjT/+dDnJCtSiGcSZe10wx7Ia86dPg1qv2WQFuPqtvJbplE+osqIo5AUAP9o
Pi+YwKVXj55aXTEi5iFXtCenV/G5umHQkvTNpPt1GbwsooZE41wtWheqCr7w49sAIyK2+TMKC03A
5jddQW7YV+qyeJJd5TMAhL18M2HJQGmX+u/s+lgFIg7k72Rg2mjtWmW9lKK787XYPCPaBi1h0spC
hRluvjGkbJfbRhV0RJ2mIppDwjQUwGP1pck4D0QuClBLF8FWnb+AkuHmS8JWszsWFIbFRVBE4lZp
mThUBxTOYfUUIkQcRb+33gR4Mo5YGeRrAGChZKzHZ+gj51Cxao8PV8cDAsfY6nseBBq4GN+GfsyF
XU9XS925oU0Ji/SzgmVAaSdV2m0jqlry4gvcOml/Eh0Dwm2GRzguMAOkLH1DAk7p4wmsmqt1VhD7
RAqoCtuB8clAuYAbAE0nGaArF8GgosX3Aj9Isdh4omtIQS+VoK76KurPJ1GNmKwcHDHogRw+RHxa
ZHiDWbOuPfITHfohGU0lCeSRDq+/rOOybt7tITbbA1JwSQHsTv3bcXeLoJERoD4Pgdc6XSPckSx6
MWICg+31kSpLXE6raDx/zWu9kIySrxX9A/epmGeErPawZ9W4PSN4dBS90tmvvBLbO//Te/7gqOez
1aVyN5t1ItafgiNOKlId4XGFlX8Syum2NY35CDLbRX4fcYFxE4gCPmdH/HC0Ozxk+tHFqD5q35vr
t8KKFYMR/uQ7u9b5M/Am22aScsQo6L94G7IjmrieHZs4xDqCrNj6W8hEbi63ayt7FHQj6rdqjAHx
ZUoJxTW5nqshU1CPDz+qvJWQwhH1BNDcR5kJ0SkQdzFs07hs/9+4Fai4NDQBbet+nXp4pl+p/qbI
GZLVBFiob79q1Q5d2BioknC2JZhIvPQFz9r/E5HSKmUiW9FOrwJ6RRDbaRp9BoUpb7WZCQ5vdEh7
rJk1x3lO8555TaV47CHX4pv0o7pjc236tm/q/G08rNw6R0+0lFG42ja3z/M7w1iULd2k9iDwGAuE
bN1H7wjKicUwpO8aJJZm1eHUnvQUoWyP59GKkjXEz06Hu5fUPMGE7zJai4h5ZVpmc8GdC/Tr5UQS
hsA0eSEnwaUbJieK0db/SwoVCcqRt/QaD3N9VNGMUdOhsasD4sD3eciptTv2hvV+ipP8t49v1CuT
opZ48oxUr35oQ9CgY9/ahQYBilH1zV8zglQNvuEASFV/PbxJkMnO4CjNbSYN2RlVcV+/olkRgTLo
PvfN9IZWXKDd+UabP1AoviLk0sjVLg4ybmamz5CdZxZXnjc2wWRAEoSffKreqLL9bD6or4R48BT/
PRvo2FPRB6EkMbwZzeU6s0Yc9IDLMN3ez1yja5mmBgERDAmuoQS4tn5pK52OeXV7Sr69Gi7UVSF4
oetQ4YKxM+Naqd5kgMn0MzCpiEV+10gmYrqXT8nzbVpVcQnZ5f3TUZGmu9u1UUw4ZFx1Tt/aSWF1
XQXtHBA/fBdOYiOTaKw6WyR2Wdidg6TA8Yta7MkTulWFq5ijAmWB7ZI2Ir8YQMKiSDQkArd9Yfq8
lhHFg86MAjs8cuJR74pVt21S+V9A5cJUZnKJ3U1rHsVXYw6M/lZuGK5R3rGZ9R74PpTyeG1TRxjX
7kU1JtGsAVWyV2sgbotE7ZWO2vx9w93aBTsbHwkm7EP0OdE8GSMm3464ZMKP4MHP1/ZCJogzHiAu
UMY+rix/49TLzfSDE2mh/gN47RJ+8fDSgKHvc1QRHCP0m+QWMl6wrAg0ZlO0bpTHBC4ibFE8ML4F
cKyv5At9NDhu89uBpSNx5Zmws97VLp+dFSF/MGkomdjce6Mx9hBz91U66d1aXt68kk64cYIw5nao
99n90k1K6UqZ5To13HHcgalgzHDepRNTZyc0b2sX0bYcxsP7jxiBEM3v75EVY8QkrFA8LRBNTeO3
IAtwrTG/mVs1LIZ/DaMqzXPJWkC4GPml1Gtv3BL+e4KJgxMZkHF+BNZhoA1BkzZEyGVC+y0VamPe
X+wrMTp0BVjazuE/6RjARuNUwAmoq24cBwOU+r69LuwyeRfkFJAXGgYy3TGGmGhGgwR7V1/z82pD
sN7HfdRAjwPQnegjnqI0g5FiUlO98Z3APE+pncM7ejDQgLZfrXY9cS6H9h8x3UQRN8b35Jr9XnI3
rdIG8jI5MQkstlLQgfkzrbzxUJAVcjezoiFuy8TB9H62OCkfNaLu3ESsVt+5/Ge8R3zpNl3AxsmZ
aMmDFzUaJkRslK3hRpkeCw9e7clqgD9TKBlvwihnj+N2p47EYAvs0LwDMfxK4j2TnLuEMFhyppa8
57KedOAA44U8ovO+R0apdMabUVeW+raZIC6IztJPGz/bvtmP4CjjhMGIFK4pIEtSt5PCQwLfGl0/
Yy++RR6QSY5a8c5LoqiL2Rr2VSCDnLXfR4s58gpblBBeNsAR59emIo2wTnPbzAzyUKasc4CemXWU
NU0rLKc6I5FkUSXVilrZSJ9DrqNdshKx0NUlA8znDxgtDtCVJ9O2XjtHfDOftqVUw1CYG1NJU9/l
aTvQgZ3fbGhijsRXGaEXgGSuOgnkM6sVlUc7l8e2usWG5k+XWqOYgEa+exfmqfV6Cc++v/Aesp2J
COmq6sCt9uKLWPKvcrlSJuIoKuEGdyc5oWESSXjUS1T0kd9jvypK9wbPcYQ3gw6doLP5Ff0dUwgj
DfnvEusxhfv7pZ6DkuLzifSx1JzZCWEXCmxiR8N/m2W01013gQDnqLcyLygT9HE9AnMChTC0tdH4
jWb0KrB0qoPSrlpGShe5v6UaEhbj8FNQ17ntoQm3cb7F0yrJEKQrcOGpRji//7XHyQqu9ysw3Mx0
Zdj7yP5DM67ozSmvlq1D3fdIfgRIiyqtWn2jcAi+QLsKzN9kq4JIevVB57eyKWv7OogkPunr9qsU
TYXIz3G3pvlqxPmtTxSlhC/NrfYucGYipwP3DiBqAOR34f6ev0lJtSebhigufM7yOesJcnLuVCfh
p7e7+sq7GfCCjArKWQWS08+pgLludszIV/josgdtdssndCMoWRAWKX1Z0OEsKf6KAMTsIaj4np5F
fQroxQut4ipW5y3SMQE7K+Xpv9DA+Im90ubm2/8DKT15zaON3QcqIEdA3xwp1mrZCJM03W2O/rq4
19fsDZ/ksW05sxUm5WPaH4Y5Ztygvm7ru9Fb+D4W1sMfCHv+mBPvIc9blvCY56fOMGYQHVeQj1gs
Ja7OsRv/D+dyysZ3X0L0cwJiy+wTaF/ktBYbPSdzKKYq5Y0rcpPgyjuHa7V8nhBkRnjKD/v8WL+Y
cq62x2HXPEHIrQUdoY9VlncQ9hFOSwCP4F3/GRM4ayXisWhJ9Y5cXgwcZXwkrL9piTxkc0VPkH6C
dzube8necUjmXzfXVf7R84dkCHJWlD2EsS41pC4BVXjt8/ivXqQb3cYI11cMVBwbbPdDRIrWyYpy
EWYEc3gqzzceOTR6ltMSozQ1tJI/XMCTqR6iuZ4Ae1wWe2oszFS3f2520tZRLyVhyObIXTth6Y+z
Y2TLUMcIMReY7mAebAK2F78gwV3y6D/EyI4F0YFFaupGc7EGQkg0As5qKb3hDcn4WjiW1sSKywnT
9dbVZQhrweq+XrALvUEob4mX4vkk0XU9UZk6T7M8IbkWvMXRW4t3dFPQV2a9MFW9Ips5ov5tjIER
wf1jho9W3aiQuo4UM00joLNjKz/aO5m8GV1Kd0ASsn6f++Ge+mnC2Jse77fnLwSxD1kKVShcZGD2
S1uZ06K15WZNCC6w0AWWVcMme7bLzSrMPHG7DSH4XogddSvy+phJbC4sHe+RB447bP30iF5zFtaJ
PihRqhzmrNkVWm6YQ/pz2uIekJ7JZKTdnd7Y/2mOdVeBkMCWTve0HeSo5DT4rnzqZQM2xW6Pf2r4
YxEPJG7H7mO9hw8OKYlXJIn8Y+jfkhgTQQMD8/IGmiG6Isub/TiYrrw9w5ncVU5OWto3Xm93nQCL
nJKkHWlkUg3aKaAMUhFH+qYKh9LOzfebUZKq7GwMs/Lidecbe0mWlG2qNDME2fzVeU9v15daH0Qe
dROriJWtkqQlPt8SbIj+6/hfHLBsnGa218YPKbQSks7GHIoGdbC/NQhhp397uz/pkLtPbeidmc/i
HDu1XRjCfRyDX2hqRIPpsZzmBl4hKTzS3wfhFFs6C48QIMFbfcCR2EUxDpTB1Gka23pr/S/U7wys
H7d46CbQtM353m2ujUYHJbkJj9LC3VyUqlqs5w3ejKIQpGIeEQavp+56NXNIl5lDdOk5/v9zyOP2
PONgR5xzNRAdgkG2hIzlyy22UX5M3tCsanP/i8Ti4AKJE2KkpnZ+Dv9Ma5N1wxmhjTos1TFKw/rP
d85Bc+8Kc8IYQBdEIiuZI6vkZIl5+PyZwC/KendIZzp8z+n6UtSENpcM14/hChJTlLHr1Q9quKWZ
FAOEvr7AEZgbJ8tjSgPCxxXS7xEoZOxLNeNrJyE1Qb46LVM0rrJZJ6RxHTiozCdL4aDKqLKt+1jb
nqLwPtcjyMLCVMxuB0Oc42zAPg8PvBLcUGx5CkrOccWxS8cDFo+Hw7W1oTDmDZJjSyPgo2Q5F5WB
McMA4KC2A5JJqDMrsc9xhfQtYmCGkiHMbUsKzMKZLqwhhgaa928LC7Kgv9pJaKQOQdGLVMskt6E0
9g6aS1uCfTC6sBDXO8cr//T6cuIPQCb17TR/rIYpq9VYDcWNQzl7pZDhiIxujpJs94ew0cD6th9h
Na0jWL96aiLS9kNQAxv/VFGsjuUeo3fNZQDY1Az0EKVbOP5z+o2vJT1T5ws08WYlqoHRMdnpT+OG
j6dESmk5Wx6dI1vfuG9XinilSYYzJdGIHfMUUUNPgGCYrLErKGKQUJ9igw7r1Dq118zu9SgpdZsr
MmDUMNw7h97WHUcqdpu786C378NHfmwPrdw4BLW6G6EfpeeK2sDKXsFScJvjFqznefmZzaWYUX3F
E63h4uESSX+LBtQwZ66Mv2WJIxeT9o+FEAQauk+1iKGWx4Ey0kspgc4nkFW36EYDoWDP399qUIyP
yjHSQWyZ2Rfir1aT3jRW0JOQBVi/jHUKIGlS7TsNYKz0iAeKdysZF2M5XKjOsZCDWMwGMvZfoXYJ
jS7MPvi3VMRz7gfBOgOXwXK0J6AFDHaFqV3Vl/p1DU3ny+HlWYxl6e3Y4o/LJZ+yKK+iEUxf+dKf
D2N4f1m8crD9GK6FOl0mkS0OlRlzJdjLos4nPGZtodNk9VWwH/jHYL79WPX1zTBheKDWpLGNsGxd
6AI+FpPQ99Zq8kj6nN1aYxDprqnfWB5u9TGF3OgajZjWx7GHgcloXE6bgBSIQ9EYZr4/NnADbHQ5
1PsQU1UMJS9FTQ2ueZPDPnXbpIgkzOm6OYQMNdawtK9whFjq/WYQGaWUjsqM+EkrWX6CxuVQqX0N
wXBUQ/5aLvlRhU1FgMPhmRn+qEyyKFfjjqZguQVaYrX7ZIqLHbQJbzfkqHoqb8VofC8ha/r3pl/J
knUip0oda3JZpkTa5tPmwyDJuz7CHH7C1Dkx98J7PWcInTJas0T07exUTaFR9U8NVFDaze+cvKil
8gn78h9nF++DmOm5tSoWPx2z2zvoqvNMxubo5I/Dgz/NmCsl4TM3CeFAaN76bhGGdgCxAPN6qbLn
C23fHajRcua7nALhYNlOVipdAAshZGBa0okLSKSbGIF2ZPqPxYcW1I6ObZnYocJz0JfaXChdd/LM
1xB/HbR6kGrc2I4z31cCPQFh6jjPzIKkifEt5aD1SFb8LwcyE5FzSJ+4lA5dPg2N29yQvEF5SJ5q
fmQ06pWKpQBfVurHg8UaaD47XxQ6/Crq/39+HaHxvjismofBQbJZEDHXtBVqR24Vl2dP+YWUzx1g
GX45wPtnq8QbzrNfALs28Zv/0NhxxzNLKQsuGonqH+Vng/bpRKFGTg0OtWdv7MYXDqjiuR3/ttDL
q7xBTcrwkq+QP76bDz+2VHdcH56Zh3GjlbZa4oVtrBzQFnG5vxK7lTpZfp482ObWEDtg8d88kg3q
w18H2AGK0QF1V+rxmK+bki+84qC16FgIXUoZ9oD7m2kcNwNtjp2OvCh29Q3aLcuF8G8A/tzVRJ5C
DhYOLxp/CRqg54dHpK5pVP1RH6t0MIaqQsvDGYT5R/jOsJnlw3DHt67C4tgkqqZKXYOD5KQ64G+j
JnFLvkfPIBfpDkYzQUOv3dozVi9xjQIlONQBp1nhNN8yrtgr2sX2n700ZDvFTZBIUAQ/651w0km9
sbw/j38vH48P3lNNs+tNXcZBZSFVzO0LjVh6OlW6ep88jqzUk+PYF3PAoxFCzNQaz0CcLcVya566
eqJdIAMbWTjFajJT0dbiHy6sz8atwlNhiP4bDYrB+kZM6gyqD9rhyJUetD2q/56XoxI/KFPwsR25
gi7JUx8PaddiHUpEoPBDf6eLWoAZWj0CocjtUYKWWCCycEAWUgo3DmvHbYAgxGQQiWBwt+ZvOiQ/
FIpskPBXJaMswPR2pUenY6NMfEy+HXITxJK7hMM1t62E3rGtbSnCojGaiG0dkGt46LDLtbsCEKJp
F+1GfraoHr+AyZM0ctajy7uKC/dqcr2IAGZRcyf9qNbt/ytmHm7MrgajAclSIStL95NgILIkpEcs
kjuy/Tp3Cj0QYcA1g9TKODx2fJUnUKIX2Ikaq+QQjL4vQRWqDMchGRbpl7OHbYtAcV3qTQQoqhB3
DcAc5a/ZdzkX3OQoF8/VwBCMqntg1DzGMH+W8kU1SjkblA+Ow7fhu/YDZO9jMuX7bY+4hXpJBj8y
tyrgYi3/g3DN1RDxzv+1MRTJlwBOtybFGCm4gN87GT+UYMDQMbt9Z6Ee5Sawp6DFNIn/8qg1UG79
CDFzGojzKlTwBauZKP0tBQMXog/bia4K/eXayInklXm+9hfnLNVKT+hMA1YUJwkW6/xT7gvI0r7C
JlkcfJVhwjfXLSM87ruINwKtcZhRGnkop7h8qNoi0Z6EWQsKHXCZRuSdsfnUN4gQFJvrnH0wuSTT
D8lN4WYsIS1Mc4D9NOeId7ZdqJpgwXJsdck7kDiRonmtbqLiOuvpIzWiEFQERxJfrQZ53U82Cy/4
vFtI96b/z05jg3D7Ewqu8krLW0DkN3+vy+6IACRztTOX1QrBNS67HveZGyd+IwDM3S8/5Gft7clC
QsFnYMqsZpqvhxzUAQw3rS5UQqRYWm39OwGAewaXvLKA/cP51PzZiAyxM8NErCH4efgEU4q07amP
XM39qJZgDbZEDGk6YX/2tgUdXBxU2MmxfB05mIWmA6W39crARQoMH54kLxlSj982gRFVjbeXLdpn
sBN2+YchsY+RRsTH07UerFdzsoCZpOFveYSzbiBcBeYi38oVLUtOv13OoH/05cHiup9QMcvog/1c
EkS+50NlG2ImARyPiopgegEU6LFmMthXYOq+YaAFfuupr3KRcbT5/jwu0jtBf6FOM7+t5llV0JVS
48X2sle2sDJPAPMFCmu6kMUR4vB3nkJKyVR3GRxLsr6Zq+dP4vXib8aLXTmXCOYeaCeA70J7QSRh
9uqNl3vWiPash14OqtqEE+GydyG5TlnCDth3wgnhFtQLe0bIPygMRKvcK0baagfIBODaTBh3ijUz
h96J+tHgeWdPpDKHqo7pYyZ0+rFqn+tVwXK1lW1PbU2BAvtntA8UXXNON2lJpn9S6hXu29pcsRzk
96OrkO7F7h03Xqel26/joGWlWzK4WcaVCrRPT9zwSg/gbPYNKdCuoRdumJvHL1KzLF1RhYzVEPb5
FGwvJ2IrMz7L+gLKyoknoIXDM+N25r4cN4uvDFbJfsuv5umqpg0lrAnajeoE9po+ugPYe0qoPL2x
BQiWhClO7IPjrACh36IB5rigUmMXRaRkNksT0C1sIanC/wnwdbr+7kZPyaaQF3C6Knjb2407zH7L
2yaXTWmUB3OiYiW09NhjntYaw9Rj/MvBJfjB0Z0BN6D3Wpa6iZw4h/D40GAEQYUThXtU9oNmZo00
+tRKph2aEDRcchkShPFBOsCuzGljxAQnLw7pUimqCZDhrA+EhKYZMU6XR7zcmNawN+edjoIuK4nG
SW9eu28B2OciqNfxnerTb3f4aY3Hla7DkQwE7Ii0JmAOyPpgQ/8kohNEtLK89HvQy6zA/aFfPtTs
MByQocwTihTQ0+dCbat2G/C+unheQ9oH6nTYC9blmzx38LUUMUcuuM9/cE61mYicnoxqRwI9hDkm
v6dKytGqGQAcqvEfjacYJ/xuqyODTFzX3Mr9iy98Z3Za3yo9FAjA4zZgzEbgxToV9mYLGCzrdRK5
i2QU4vT/BU4Vbl+Xv0PD8EXpEZZvfwpkAyvHO73WKYlC9wj6VDP8XOggh2SI+Reisftq44UVw18e
KIV6qUgZHEWwHybuFqSUhvFmUpA5+D5xAk6qB4zuJfGdjcyE/FcEnl01T+oaemP0GJ+Kj50GpOid
arwtS56I3KbOAfv+o3Tnbs1Iy9WlbFCICNnYMzRMQqajccDPnfWgjUp9VhAmAWfB9RaEUb1psX58
hjxdK37x52H7EPv7JLTJCZYumDFKgxH9KxSMgaYaoAx9ia3IUiLDeDid6tt4RT8LFZvAmvJ09Mo/
nvKIFgARiAnVRecPfDFtCNj+7pZsvPH3B8GI+X5JA9TOtEEM1FsTp8ohwMMFcMHTLK4X5ZZ6Ht56
3HZA3Hz6ciajKqr5aQKgpPWuph7j52QfEAI0yNj87trlSf7CUrkiTvhQPBeUr7GYuJKus2T4v87C
RypzqM4KVjrZDWpL78jzd6oUq/+g+E1v/zhuIlUUlaf2hGvMxDKHtCkO/sFpL6wRIUHuiK9Ugm31
JpgKXaOuhQ39/AK+sHJbSyvRsQuttYCyj4ab3eHfripVRDnRZsJpnsU/SOnsNELmURy4MfzpxN+e
eHw90p9VsG85V4za5tikrIL9Z2sL517mpUST1j6LdJ6atYkmqOEk8Krd/HEaf7XE7Jny586vr4f2
csWzm3GMdCicymMCOh14R/SqL8Ca0gUfANAXwMdsloNUgO0DsHF/Vh0bru8ZppMKb/eQi4xGA4qq
O6iiXi7kzPykitEhTPq2pcdMsv5iAGIdtddJVr00fwE8GvYoXef02BBIYHzyQn8xAK6JFUoaMro0
qIhFN72SX2f/6M7PmAVoOhYyGUHFetmmVrj5HpestUaXPGiI+Yg1AeR+xSL8QbY7luwv48kI+Cpf
472f8yZXtOc1gki+tS9XJ6m1nbYlojgeg6KkY5jr/iPVEDUgpv8NPqdZmdVUnzu6dIWys2qDv8MM
oBHiQ82kgarcrxWlKM6z6ZDqDuW7l4l/NborocdLRzGNOJ5gn+MIMtsE3GARILicKDQInps11W+g
2GniG/SvV2rMnZNM+RfLNW2k/SBwoJ72uRauMvSco2kTSpPy9G0znGNsKlhQvKcZhCK9Vj6O2isG
t77mJrESulvGtpMHxUISrZhcdzXTMwrjujl2dqdlVnAbnhAbgNZomG0lGX4m+Jb02KjeyYbK4uBs
GQV0mjK1u3G/pLsX5IAajk/k2lwsN+IiemAJwFSNZtPjVVYst/DH87m0wXylCZbvoThbr32nmcPL
1Jq8RRUZ8VOyWp5Scc1mXDP086WHLRLz8RqJWM/vTuKFOMG3zciuRYnh49nPFoKMKXhU38JY0mKa
s2Tov9MKVuYtirphMPyWF6vEzFQU89ddegjCIJ7H3cu7BoayLAOmc6a39c/Zzs9YuNCwQHp1phZN
DXfokA4wNmBncclySSP3ku1NOcPn+3jYre5sE0x7l83D6MGYmb+pEgoCJNI1TPQtmcDDxFYzEBy0
WGXo4yHOjMq78kw1dqTUumgWm+5pxZTlSlk6rKNqjmcOL/w+vcjs6xs5TuZqO1T0+YK2IPUfqFOx
arx8P/JaUba6cZ/SKm7bN34ky/Cw/DGKeijkdxP51w6aDLkCrsq8r0DdA4xR9T9P38Q9bhbTSeDk
GNsVJQeLg6djdrbiglfeFwEe+PIMWcy2KgeJ4d3U1p22TfxQXuURS2yeKKBsNUWZSYAZdDQKn2BP
lkeE7xAdDKDeOzbmfCWZySjEj4cDwBk6hfKJcIY6tboWndvtFqPh+ZMJzKgfaHooknqGSda7rYG9
iGOZ9LFg4YjKxQTZr+vb/y5+XApkNC+StDOb1TVL4ip4n1mWswmtEsyOqL8z9QCLzfHI/4OVYl2t
1GF/uPfExZ0w5zqbYdNSPKQyn9uP+4iNsoVs1G8CdSNA4Go7fdhPK6je+B5S+P9zoOEdmcfMjf88
2o6cWHKX793juqTwEamk6Sg8JWnMU5wL1/6RNKTNx7aKfjb/VzInjv3FZpEhSS8caDIN5NKkcyAy
BL13oOPQ1D2I1z/qAzotbOmDdwCKTXZPdo7exytgbhut3N2XtjlO55WXnxKrM3Jw0mFQewOQ6ftY
egT68xmaHzr79XgfH0Wq97buD3DQRHUn5QaPW7V/FYHuNVGVquerSiWqmWttPpcFBRiLOd+4grpX
ej0RXXeo1YQ8QzyPjufkMXwop4/mw1v/wJzKF9Y2D8I8l7CRUHMSGFoY0LWP3kI776WtxZE8DchW
iDwFhU/AGb0QBu0o0ctiurdtLT8/ryn/Jq3Odirl4BHXal48qMT+Zkv+c6vqnEG7GijHyJn5yHfI
XZGmhzeJeXShe9FwV2wd//erGUIrevXz149e7ntGlpSOGS21KTTtzUoMuKVnrX5OjnZTWKiamKxx
Ii6luQ1hw8isZrM7tjdZ6jKJNdMNIyFMUf8R92PHfbJzFLs448LfOAv7E5laspUWo6fs5M2HnbJ2
J7Rx5lACywWuq8xTDHXGjyRDSndeYYK0/kmI52IyVhx7gcmthYV2CRQINY8stxZZVxN5yXObMNrg
wGd7aBLHOBGs7v9xzxlwzYwCPgj6Pedd7mRjjJ/Yo8hJG94oPACPvMpORLoqHbFGXCAxa1h+CMXf
cXW9xzQ4OglZ2I31EFICDN5TUAl1kIg5xzLl42d6M1vXhBY0bVSC6pV4nNW+5XwW5qDogFK0Cujh
1wtrG/NJ0CwZJ4MxwmWHNfj1Gu6SOmlH+eWBb7993yxHF/anC9lgnj15dRtG7uufTUsJ0tkENt9W
8N0IYokx8Ci9v8hWAYjZjlyRBsiH6D/vDz7fDV5DAy7iQXhBDy5MdgmeM1viQy9YdXylYFBq7kEM
/jSQ14yFKCOlO92FLgGVdQndGtg3l0KV+143TgPvrKyPd0vLg20ss+nf9ESCh9+QvAv/ocmmIEeB
h3lwTaD94pcoX+FIurxJ3VnwpWMZwkm9BXRk01b8ZOKrhcFVMLsOQbd1wpY1lCnN4IwMHdZjzwoN
uW5/iLd332NikH2/jx81OAX3QWvI5/sL5Kq6rxHgAcjSELd+9YT+uJiTpOjJt8ngKIgc85ecgJCg
4+Twl8A79cxSEgGtdYIgt8uPjdaTIVm0+Dw/+UyVitVu5nZsCGfxExiSQFkbbuba7+9BNcOumE+J
ttdpX5SRBgmQSnBYtxTptDoUrcrdDcsbzQiuNS+RFJLVucikga1N9S5GXmznS67ZfiDfDgXr8CPH
c32BA5aBkpnOivzxydg0I/zOFqAuSE74VGfAw+szNWtXR6+MU2GfGLBSwztXPnLVrvlijKARUP6D
biMsMp/aDhQ3c+B1Jd8xvVrqygQApmsKwtAHpwmdVZEXy1ihCOMjzvhIGDDiMTVq23Fty0o+mYzn
mD1vUfyXp+XxcRLkcNpgtllbIDgQbp7gxF9rKGTswZKl1niaswJ3pqmOyIo9xFoAXDn5+4l1/2kE
YqCEBuurHrCjJuiHBxAmpMUCKJGL8iTnfpTQ2O6vu2Ez96ty+kHykoJ0/72imqkXIWYIpftfW8Cp
jx5Zf1MvqeL6HMDj8TKcnWjjmWUOG7U3NcphZ3mwpgO1GyzJr2Fn9KJGtEPuXqDGjzHvZXXSGiUU
n3YGrNM/ZwHlczoQXcT4/Ne0d75cXpwUBIMhMSwh8OV2U+JiVLym2J/ZzLiUO7zuW0FiAeuja2+o
ffrjy3p9Ait4UqpREFt7tIXIoy7gkBCofaO3epSsMGAVsE7AydrcGoiBuslT5qj3rOJmS3Y/XLY6
avFzDNoWEu1tlKIC3L3mCR86O2mp8mOWLY/BElAXe0aavuQp+S6ohh7eFxrtz9L6gpbb1ADQZDYc
5Dwqr0T9vlhVZEMWhDvb2YArch9b9WAgyYQc0vaBWXSME2IT6JS7nRrmymFjSOre+JbwzU9Vpy7Z
mkLRk558ormd6dth8UJIW1mJXTqnwMIi5f3LagiyWyDAH/vNrH9+LKXy8QsnDb/2b3Omw+zKtZcq
CL42RfdEqjuqzz02FO+V01QXeoj3QbZBhh1PT2NZlC7OYWDTPY36uMLu+KOZNbOCHZ7lLRAxxBzL
BOhiHfKjhvLSyMOwoVqJ8NeLhSGjHqt05ZHecfnPHk0FTZdg7CFqnWv6dgipvxUxLYPbZ2N0Qpf1
klIlx8eVThfGLwyW14WhifcttYel+QHM3nVYxhYu0y8cmV2io5O+msyxOg3cHLK1BljJ9kCVYdya
NGWEXZm8R9jfa7EWY5+kbb44sZwly06GaMty4bNNBBQCaUjyfEvv53lGzEiTEWxQyU9UNWLsxXAk
xcaYLM33Hni2xQ0wtA8NH8aczJdI78BjqoSPGyz/KxqsJG2XXy2xo9PTXRgrUXjDHlvfRPwuMPXh
ucW6u07X86Atmce+guLQs1+Qh+R7U3hkP6392c/OZhWwxgwGt760IVRAxoFumelNoxR7ltP19VZ/
Mkr60S/D3/KRi3HJ1wpNx0pKQaH7lFjjvOpHJ0GZ+Kt8rpwzZWatjZGOWvJ7A9I46/Sxxa1eX5Lt
XYlL2r/jIBbVGbfSfpdE7OsBACmfjJ50XbhhtgtGa2K9LcpT4mEr/8OgUAlWjO1owWYPXYzc80yk
hGjeDgr8+XavJkbEoUYbvfV/qTMH/kyAxyd+/HDs2hi1BN+4jLO1ZDzmKRNbZjTtyODZOX5sVlAc
ZY9DA9vdN4oapq6jzBOrCKqvc7s5BpJm2lWQo/1kk5KFHMr4aqp+I47ByG+/FSlWis9jZU0j9AdQ
FaoxfI8XCTCQtReE201FVK0MA2yKRJks6efGiv759Pd6MJexiDg+QCpErGxG5YOu6+WKhFBhqBss
jC/fi6n+/OwovWVz2UTWWaE+Bq56FJb1rDpFo7MfBxUOY2RtyrVDWlozV3ZXfOAmPWwSCV5xguN4
kd2uZOi9UvXpYh8C+zFSzVVFbpSzA3FUh0H3kfda9AJD7vSlK9ihNfHxYTCmdtK7+xNFwU0AuaB6
uH/h/cPpxmMZXZfNeDPR1uxmYQMYq6gOzrqFRZh84aZVDyuqRXWi6vDteakWYwquqWsI7YKkiDaz
n8z1G+m+gMrJazDYrvWhU1WVtnloqqDwsytcmrOAgm/HPNSa+oTxZeecqagi8fvgMvXx3pgh9IlN
Xk5SQDiVoVKjoyscOMXBBfH0pt4i3DiXxP8wSNFux0krWm3awhx4GXS22hlswS0ups1IJ5wK8ttA
jF7aiUYmNJFqmJFJDCDKKxZz+4BBtia/ZuMvOFB8OhURkFRteHnedo+C+4kLp4peX4JYLL4OtgTW
d6c1eho3n85y6lBUqAgBgtds5Yz27Y+DBSVkJOFL4KOVouwgXv6frCQhZJR+5Frfk2g9ZXIP4MZS
KafO6ZK1JGSrHSiMyH6HcDhgaAMEN+nG+lnvk2vQtFho/EjOHgCfanXutUKX3pSrM/6VLru5a2X7
XYPKM88zXVAWQK8YXAYdWqhxw94Wd7XzVGL8p2OQ9LPt3K5LJOEzrahVAEprFNZrUQrkx0gsoKCU
xeis9fOqqnMO3482G92rO4JYbwGAfsTJ8Th8CxJS0x4PwfYh/JBOyPr5ex6U0PFwfWoO02jRhYqx
IlJyjoV+QeV8X3e9hWoD6p2/F832oDa/aHus7GSvW3pt1LYFUqa1PAmQTAXQqa5L9F0BjpJeQvB3
NAgalYHwvgI/urTqE9I8ag0AR00lhj35DhjfNJxISZPBG/Szas9DorX1gVQWG/V9fMbxGAKopf0l
y4EAKNYfQth/ULSWWX2gq2FFSBmT9ehgMf1vH2khLOJmlu5fxpx4iwnHT/LA7cDI/bKuNm2Z1omV
TBjlS8LESEWSATH+GVNUbAPxwo+2kJ4umKd09wuY67T+Y5NdNUeh+/hSz3kMdzBRwa8q4tCwd6C7
0QH6fZKmOPY9RqTaAgN3LWYNdzFbzeXlPQ0b/8C1VUnonJBDFCp9OqW9dcCZZMeMZ8MCNXUvUF5v
crzsewMsPIznLxVBV62RDOL7v36mCvkG7NTKzR75Hb2dVod72k/R6JMI2FpBgjUfP3QESzQyJMFS
oZ+ke7s6ZjImPs/v5lOSwFz/TCvpeJs1PzT4GuXwmqKHKNcxEJTvaE9LEOvsW/gQH75K9U3t0K07
YjFYmtETJXpmYmPzF5A0wUHLPox8lz5IHEY/vuiL6eiGQvW8XS1kjhwNZ7a08H9iDf56IAB8iE9N
jgtEJHxFasuZDMctV02FMXwAVThsUVwA3Am1T7pWEIi8qZDSkVfVAgaVjFHOqgtUGpRV6182FE9o
D0B3iBkeZSXvutT/xDVTtHfSEKRcfUfk/hAJBfw4JP4gVYb1OdohKiocUG6PLqyehNVqBGlKCOUU
XDeaMRkY4gFyRHJ1ccSSiEgdOwTIfmle+L0bqQare0uqGjZv0XNVon882ZCw4CqTls7ntK/3vx2N
mQwVwhKw4C3z9hcy2FeA9CwRQ1pUCF4LpxoRcv2i2ONv+rEkZpQFzCN/hZmGcNJh82v/NIHNOQdK
Ws/mMK8s/EVksfP4iZYQ4zd3Ce5WyEePqcLTaFiFdNYcAIV6hKC3v+IuJNkpbdIV6QlVjO88MiDx
C2iU48/Ui/7rLU18AcFHiUNzMxXZpbFen1vdj7ovWeBxPfyoY9KJV/2SxXNOnFCcgV2dncXekLqC
DpfPKig/2WT/BoV9UqhcLK9rEDyHtr/zdIr3K893TpEqWj0Zz48RQc2uV3vTcQ+43PcY6Aluuygu
3ErNJIra9Jd5nB4c0ySRf2TEVEYv3o585OMy9lE/d5Pgg273Byr/Zq2W8LxB/RSFRMotcGHIxWS8
RqBtlh/ZW/qQOGit9BEak3RDHYIeSZipFMV579Pikt23rF16/heqKrycbQtMGdfwVvmwIORCeQYE
DnHjctTImQDZu+3xI9aXk99B18+S1q5xlfpWsk+N0+TIJMjecf+qOvi/IFwpjv3VObgGDryhXRT+
g+8XWBvw+3tuMVlYvsJ6JgOfmYiHofSFZAIm/+yNZtUsJGBJV93ik3x5guIxvysAoTnkaC7hFLww
64TyVRwkwC+ea+cXVOJoZgvH22Ku0Vi8InPuJaBSOrjgy+ah79vYQSGUGNs2dv5ytG6B23BErGVg
7FBT4w1aXky7JN3cu4cqvdmWaTPPpaOY1RThNRv+uxPS5pcNAMeeARP0DPEheMmdJ6Qq13xMWizy
Sl51MsfEpjSdleF4YmtyY1IKTYylnB/lZh49wA5NL0uke7mtwS9ag8XflBwoFTDCSmyQakLLNQUT
T1zVGy+KqI7uT+D0S9LcXGCCp0BM1b79SeR3CMQ1XC30mbyymvaHQXm918zwa2u81fbfKN/IP2VC
N+Wdy32PVRWcrty5Q9n8kmLVY2q+6TRgV8Yg8wuWXO84klqqJznYANa7itUMb8mOFQo2kPuK9rX9
V6l3ZobJcTJPH1D4GKfFu9AYFIMGVnNMoxQMysO6fjSybVeM3vHCTIWVUIQgnA/xglQLg7dIZixr
yurHahcTi6y1P3G1BLkReP/OMLuF6xSkhfzG5nMIa/EqjXJ0bs+6bJqR8PvjmqX55ZIFbk4/TFh/
LjgIQfx4V3l9ia2xRFsDx2A4MM8enGQBvTo60ZhGpqiQxi86FsWZ/EWajnkFOd8DRhETwAl/FedO
Ae6dGuN/CnZczJ4s3Gx2jbKlxHJpJqH8zDO1wBdy232NBHP07NRvERBm3XHPzNfLGAeG8P4H5Ifk
3Q7zMfNqKSRnxnsUdMEmDMXoL8TGTRDFeqDnR6KDt0JJvtsDW4DcXj+nLtsUnC/FIgfzJiHNZwoR
gD7r5aTzxXT6LtIRSVNYwL4fLEIoIGcc0jfxG4pQmNA8tvzi7EdnAAvp6DfijbvAT0xPO+HXuYbf
dSM0egqHcdylb3N+GZQJ7871WNeOI3HPGcbJlLD0p84Bfzjx+Ecd3MTNwIDsBQyONb+MarvcKUT4
6g2Q58FjgnOjHyj+EuGcItyxgDJvdbp9OrH5WOnQEDc9xAwpIt9014PZZnLxpQgWVHOQevjx8sdQ
WtdVHh6LtITz9cnvmAE3rgIHqW64cSWd2H5kL3n6deAHV8gQplU4PzzLAF2qs78o5u53fci/uCXc
Vt8RmTa4dWIGI2/dk1w8TLI2amrXCy/q0divn1Tzshal7REyqjZN0aFxRwGnoGYGWjeaqH5vI75e
rhOQz0QcKZH6NAY5VXi2M61riL4Q7hC+Ogc4aqco9krxTPGu5m7cSeVL+MOuMIRgEfUhXYheakzq
yPZHwvcMQs6F/KZiKitm+e1oAKRiGckxJkxL38eLmqXqriND1FjULgEzqrQ5ZqAjmcXOVr7vn/+B
8dHigXd8qnauuqLuqGPNw98Q/SQgJLAhLPIOelOtRxL8B712V7C4lapv230JmrAayhrE8F0aZY7U
HeSxJ+ELSrjzKEXChNqMAYeLs7yUMR0AjaHNayA5g8D4kyHZSJ8r1VJOelR9AQTzbWDBe9w3dMmu
apdqfqlLBDQ2U1AVXB3gE6NehUV+YfrRq2KFIF0EXbTH12m73+VZ4GXJmlXKM7prlX4T+L4krog7
aAMi3+PCX4EQ4Ic8Ci8NBuQtl871YmIwBcebK13rYkht9l7k4+JuZTVpLZJCIVlso5ig8Zi+JIwL
DrdJZBUxAYtFPpyCh9F4xiQnd1nDKurVRDozuCHW07unRyn9FuYMkFWmMykk+EZyvQnTNZVeksmK
GXckFaEUMVnuY4K9BvDXU8E0yHry1HRzruLViiJx1XqruKk9CpXCImewTWp/U+rYl9DhgsNGCJY0
he7ivHwO/3PbgHbNveSuZFPDVi13NpFQbgqGTQIlkBY/T9xfY94KnQ8K/n/YSf1+Z6I+B/9W8kcQ
PRgfvJYsAABYEdzpkvs4fXGT3HciBNM27+ZcpWHJeHXJ5hnlKAW0LBfAM/t6BjFIWaOkY9/8yCID
NncLyQzwLELHY5oO6zYZRkbxSw6a1SJAJeGW0CN5kYMJ+2rLvw5tP5v/buXDquE29ISI8jWSBavj
Zerdqeh04kduHTAqjnN/955l8XAbI7CmnIrjrZQtRbqdgZNPAFA60Y1z28JEeIqi7dmnteJ5lmTr
+eIKM8NKXhJ/43l6z7j/M8q1jqMLhex+rFCQjSpFyqIuJ3fJT/GO0w3sNw2eN7QK25XCzGpM7uVJ
itrSCOtWnf4zFrO7lOSqytqnAKbEHzdAdXqN3eNLsY3N1vzHUS+Cnhh9gjoPo/9NELUwMTw4SDuc
boKtx/9ZbryUTGPEQ1Tw8Psw3FhFRrw50N8UjlB4rhmKWrEue5LU69BZknVsiLKvfWXpyfCj+eA0
OGXdMJvmh72mOr8rBk374UI0Q1l2CX8AbV3jxSrbt+C+TD+gVs/AHPjOaT6zlwIgusDoR5Yl9+SP
ZQ7L4NdPtvZAVtju+/EzkvyiAnJlISV/qDn0VzbBgSr3h1KmYdWVo1a0sV2JO/KXWOHyimXf2MD6
o9BUIs918O6DDnrvWhLUB4UUa8nIrq+unn8gzP9Tc7lXY2qNTgVXHpviAXFs3KJZarzQLjgOVOgH
VMdBIiMWoNsBksMRtlU9suAYBOxfpChDyl46EOILauMRG0TaDIupRD1yyAW9a1+BszowCPHGlL0t
/ccUT9hu/6W22n0mimRUpJvKlT6sFbvMxIRnJXsL4G8VPV/u+imPJYt2Uvi10Lq/2+H2SkklXaKW
8gCnT8lCImF/zB+srnt6YavGEJBcLa5mdocc12CnC9OB0Wd1czGTr5GarToEmqojMWzr+9PFfB3i
gcACVZlfh0DSpwSO/rOogICuLyEhzq6tUdND3o5I9VtMDO94j3Mv7e2UQ2MytCvZsKhfCUXzD0X5
l/HXbBN8SFXKLeaOt7/laVf3rM125wYRJL1YGRKaGrMwq+3vHM6HJ+qkNlNUDnaiEq5U7hWUbDSW
tQ0mN7FBuQQasAwQVWAKTEH0dNFRhmSogffK9mHx8u9gRXggUoHZ0cMNZvuJKhJG5zr3koxjUKUr
YGvQKLn5DuBroXiVJyAd3XJeVQGt1G0qbXrdNByVnqWuqFIOwTLYhEIx/DEDBpZJ6HZD8tfSc+e2
9P93xdSrjSXr5YP36N+5n2K5d47Sw0esZmkoqYifVVPzibZ/sEQQ0LkuNe+n3LWHUmOvTE6K5VSB
OfAQyIjBJxp6uAb9Yggm5NC1EE0FAH64bMLTJP6+aDyZwhyvaKi6r5DEcU+hGQtbYfbRyuZjaaim
phQ+CJvgigozG3Cjzmm1C11cAhjeo3+qpru5ZbgBArN77zmfnkcgc6qHKwRGuV1eHz101cZ8rlZj
Uj9vwi0JIjk/h+b8IKi9GBMkVQRYrrhHKPIyghc5ilG9FElLQ/EWtlrg3jIg3IKad92jJXCFLau1
TehB3LeKO3NZS+reRuWjQVGys97KprPU7ONv0DFAwTmXM5Q2NhbQ87ajLdBChWOh4fkoLHPJaXcT
w8HnCAE9TK+GJqpGmYLhMuDlrwhif7a9fjYThQMDEUFnFrytebG8hF6Nkqnk7O+sghvkZwdagYX0
TVcNZmq5xPzUPohizO1Zzde+780CYj8QSsNWTC9CjodttShDbC9gYCKKVwwu31a4qLgD4pS/U0um
MPqxdDHnrdLleqfhnfKXRX27se5AH6a5qSPKmor0H+PzBLm++VxIavdl5RFpIblAfjYAvNXIitMl
nKKA0KUD8n1TTmzNzuFlPRgsHt3vQnTorNx2t0DtOMMhfgd4OmdrvdeI15bbQy8aUWJYdpXSS9Vd
/8bRMqC2lik6ydJLRtymFUwd5zxkj3AAE6yheoLz4iKiIgCA7eDIT8R9sH6ToAs+VCAfiWSZtYtX
u5Jw2+9n6VCznSamJPV7m3fmtMXz2wVpPLhiz0+QH9PbGTTanACCwBANUWyTKvV69vZt1YWcHB4W
fqIf4RJa/JkZDQtVJP8ozRuM73K0UkzUkz+L4yyXRpaPfTzxrc0bIEKk5IwMPEOkvNrqSXLX0iWf
UlP9cOgWiCFmnLgE0dl1D0dQiu/PqwIQ5DnVjyJzJm7pS1JeA6NIhfNjVTPCUXQ8uVRHXpefgc7J
UU/CUkmCYAFWbHrDij4tvT9W58x4Y69F8zvwYLX7Y7l0Osj6qjNEIYLOkKrIUj7r9W303+parNIn
Y1zab3PpBg64VMx+qWgVgt9Gdv6bnq2XKn5XDjZKGOUgwnmpgDAaItkA6vIeSt0dVVOy8lmRh4Da
CMVpsIpKZvx5x7UQ2TiMm+lZ3J7bhwZPv9dPy8S+iNRGLa4zBCicFfiHh6Z5ZWB+zFtyipriypkE
g9p4w6p5/bHiQ7lOlesDSLJHmNSUWR3WZDkJLgiPaqVw25NFvKWau5YE0yBLCRdiewnfto7e1biX
fwUZ6JLSmoTJ5E8vKpSK+b0c7UxbpfxlhfNgwbRSLzlcjgpgCiKMsb4/WNWfFA2u2xKug6dyjnfh
5ddpphmrVJsYNNwAxgOu862E1kFFCYI3X0aqRROSLw7G6FWze3Ov7kN4HO6I7WNitEjLPNQOAHfS
ByItEMXc5rRsbftm2+T8u/uYSDiudKCGFQNqq9l3jOdrkyVIqWsQnFPzPbPRSDkyEP/0VZRfkrbs
mHvj2ZLp1r/WFvzFimRWRrAYAEdBWkDZRPa4qQYqyC19uxP3UKNQ5qaVeO+S4+Wk9MEihv7CLI8J
5a1iE+mvjYJrtMmKkdg8BHn+VTDvJXfVf+Dmi0cQU/a3qLdgQ+gi4Xlu5i0ZHLUoDkSGelyX/C4Y
AmMhFdQwXtjBQmgexVKYKzIfbwQZ+vN+RxT07wqAPIyElSN0rP4X/UPe0dghfWpJ/0MxQANdP09n
Y4Fhl0sPKPewoG7HbK0hRjZaIZ3QUf4ceB/6m9MPUZhfoS4po+SGYIhLLA6JDPXPwc32ypoGNCQz
IhA2C0VJWgL0ArDcybvbT6Fdwjw09EFLbO8foMMKZtJXXTWSNtHNVACJUkzkh6lUDKLffAHt0oz4
G2VNcQajYp9WMrYZ2x+uLlEj7JzjkvTL1+2QNxgxy6fjqo8nXiNZancjkXmM2IefW1IPBKQcc7gJ
tOsoRHqpj36N9drb0napH8PNFM6Puw3rwek9qI+p78LPOiMmXwjkvNS79HSCqLBW+VFBV8yt61LS
R7Qlc+YxvEEaYQL3jC60Yq+SubuTggZ/8eMHsSbeG91sJmUv3K6TvUKkOmUI9YlzF6I+jOgFjVNj
n1e71sPIRwSRMR4YYCFaBRl/A/1Ko09FUzpeCpemxvvlbdT5HGUrfbWWGf9ZS+gCLzNiNuGfAz9P
tn6upmwr7QOf7qAlm8+ft72lfhpN2SI9F9POtDBebpBz7vdaU1gixM8Y5avBcbQf1Cr0tR2vjOj9
wAAR2Im5dD3fWeCjdNmbEL8ozAWSHy76i9GMhxg6TT3JNTxg2OuFMkcN9EvuPRxqRZU4H3nkj8TD
vbJjcbixxm4IYE01yax+BKo/hYFkZqDcZF3/a9PqtzU2VCf8WgcQmRDEZARSrQus6iGp9HCXKBDD
6aEJu5QPFMd10inXUnvYiMgZHHI3783zJqkczB+lscabINCYrTt48CLySss45ultbau26kQx5+w7
eiNQpMZYxE8rOvXfTIPFKKOeVGVD8AnGVczrDrb/jlDJ3cLqOE0KTDA88X5Z1gUYxKvHfb42ZUZs
hTjqbBoIK5nByC6gRBjDVa38tXeAKDu/z/zJEMiok2mbeDuRBgbuUndew5yULfU55ni00L8QOXEH
5sKIDJp2Yb88meE4EjsYnj0/XSzmMpgG0EBiIeAXQSMjRE/jJkB+2Q2sJo9w+mqsATjM2dYJhD63
0WXPDwVWzbYstmkRj9FY5SAFWEIccBEIx9QE3ho4vwOqY8M/VOAqO80E3nQhN9u/RdWlQGaQDBXx
1e+stcfgC09q9Mj3U1QD2u/1fHLv30wVZpPulXTzgiZJUQb5ap6abR45/+vvq0eqWBle6P/SWCgf
aFEEYOg4mtEdeTcngs7fV2knPVdtJ0bMv4bUVsam9mhAnm312jBNaZ7uimKqvnTiZqiqyPIH93i+
QUwTOqwyIc8FgV2LMAUT1y+K7N2SPp8kGAeMv73+7+eVXJHFzvfz5pl5UlJmirO/K7CJuOtXvXVe
eO/kjBzd34YOXd4HZ+d/WQeRCvkGTqbNQQGyDDDvG69SUKg7pWJuJcIw/Xcgic/8hFmuEvMa1EP9
ld3IcSY8Np4TlI3GU3SclxTgkA6kch7pH8JHzsEF/Syz9hGQkND23HhOmG+3KxDaJxWQYTggcadq
PzwMcZUjo7YNpQXc9Tok0KdXO/PArmfBUGGuB5pWmXX6Cwt7cG50UiSNArg2nMVeHFOHcoOeX+ya
boxXcmAAtvGFVtm+u74M+A5WXNYzOU9USAr1mT0hxG0iKVymWvBZkaLHro4zFZJyZJE2JYgN/eAK
bcr1aX8CtWY8eSR/zh7aypmeqBBa3K+HsZGfj3MDLlRxJ32Z2n+vmpbO+7tKvOTtW95yKRTalmlm
FOgux+fOE8SbNoyixN2Ma+WvJXR1FOJQyW0R0S98MOY2b69b6LesLFfj9yBfY/jlfUXMUaenA4tU
BWimXWZ9oBFL5OTmDsds+eWW/sDUyrJTGEgV8asAbqiwBH2q8SJnFeJuPoj02B4p1QI2xxfRzpry
uFGuPs5T2jEiKbcvzF1RekPHwkebRW3ZgFKO1DQfCmkw4EnjaqNYed4U8S6Zse7CHCJTXTHT2gpz
ekrXBgf2mRyYj/xJ5w07aEO3Evk1BwOvfUt1ZNMU5qWUTP/1PgJkrDMZ8TkGaW8C172wpPe/+aYe
WqRpAiQlgRI7mzaCu8ORZZJAEVn5KljPbmT0Dz7+MCipf6q83xXVioH+7wklHvZGh+GS59R1lqhz
J7FN25cKfX8kMF/gDfm1zjxFsaat96L5K8yL5VKOut3nYhUVNc36+glQ9RnwNRvKoJmKP9KvtnQu
9MpoADZxEV4Zp1Bb3QZfAz+iglMVeMmcLz6ncvrGQjUe6h2wsWPBC6MfnOWxHYZhpuEf4cgWDvn7
nPLPdbHOxfUaj7soUDpYdJ6+QpTaboCSyos2nwiOEwV6UPJywisYVZAG6iZammgAvn03QSqBh4O0
uN3ytB9us/A898HtOJpazNaufc8sjHVyMyDO5qCCkICDHClOxhdv73eeWR1OJXzWDH3qSSTsalQi
TiXxP7chLcL8OzAkQMKRbezBIUbaPfGT2pJ0Bi9gWTzPLzTazbcDdsjdgqCyN8wE4sUNQMnu42hC
BJuhQp6Vvmo7l92pEyyzF0la3fKigZmIPUYNmP2erRZx6qVljdBt/wNrwKqgbPhmIdCXoBMxZT/8
oDlm5YPlRhFvVGauPhIT3Mbkozs2VzgIfvb7fA5Bi343r8ZPsohPxx8qkSgQ4NH0C2FqNPUZDfuc
KfI0tVzt0aYXHaX/BRFu4pNRceWR29TvMrMA0j7JuxHtz3ObZpPNGrgQGS5CZoL0TRUJBfWQkjhy
RqjwnuFObkA8hMhfi6fOwOsyWr1NcFndmylafrVOpFU5PJ4jsWgoJqHiSPQidscz5UPdm6VH7qPy
TmBYOkVYN/e4cfcIiZAdDlCDZ9+UhXoKsMl3eWTelz+wh+3+e4wnvF1E7nowofopsh84THdpEiZP
5DtbcY+AEZ7WXKF48l5VyfodlgvmdMyPQ4neNpCdXSVySBCFdOmydHNUx80E6hVqFoeneEOR4rFs
ihjuVQZjfQQg4RJTgg1xL5DT2y+0sX7Fjvo8IPwbbNrTEIEOAacBHwAbxN/Yos3hwPWO6DzH0rXE
TuEata2qx3Q489GXmV9jNgJkQXy+09mRWMaV5lR4Eu+AI5ZJHjUzJ97WhtYtW1czJk2vqkNKj3yh
HBJJ1pFvCvyVAy1Owehzj/5ARJM7MD6wb7+S7uX5iUQU4AX71x9BVK0Ejthdsq4at0FcpEm1rqBH
JSVXxY9wkkfVUx+U4+9u2rx+5aNYE3wMRqIdb2sdbGJs60Xn++XKWtqOHm9JF3zeTaKkpWLNqc4T
RAXuXoz0CpFi4Lc8JWr7aXqioeGAYsQzv46WddZDSHfOctYAtl+RmEvSvOV0xDBBdDgXR0t3dhR0
GNYIgbIwjfPej4MAERqNk5xsZ6bFQPmbnPCD25dKmVcd+pYQC0Ru4IxYfztFl9Fb9bNt7kPUvLht
W20eFAhEsr6bdpkMS6e5qdDkg2Ouy5KS/2QZIsTVsFR9xxhvtQ4dHjEWDKFwc6rhMErN2z//SoKb
oS5EyyyVXxZJjDUTxXxwwDxYTccaA25mqmdPN+7w1Bsx4GtFiGWouM3u7dCrq/Smted5L+FHK1sj
NKiGKXWofgzU4f4kqK1Lq+fJbMgbWL/up7R9keBTYUOy3pV/w41gTsYogM48NJ0NHOiSPmvjXaIu
3g9aUmwDvGQR3+gb7TP1FsRD+v/IKNm8oZxs5GcPFQAFyUYO7e7kt2PqkOv3mofPWBqyD5pBTRep
OLBdMu1oZ7VIi8xowmAOEa9QdSKwBKJRnj2vGCDR2b1XXYdP0rrsO212eXZF0qdT5mRs7xUAr8Rf
nYvJCiTSd7UPj44sHMTUCs0XDCIvSFNKxhOvM0D8O3/GBoVSTs8zSwwT34WbVo9dGKJKTGqFA//h
6H0ZeYfCWvqgTcdfxjWfiXsagL1UPPJp8TOEVsIIOr3cMYzCiLm45SZGaHpT5ZnjRPWI8jFfAO5R
d3FRm9IRYy+JSvYPwM8bPOySzw50DEzyFQUOtBKk/Hweaf1yYcj4jYEqtiY+qeAz7O/LeGEUNTqY
/8qd96FPQvN70XVaa7dWu8CkvcSllJ2WYUL7lDLBFWGchQ8OMp0+gWKWAb9lO+L1i/tM+MH6XFP2
L+TbOTLbAhc9im+oj/uChnX7WPtgx0kLT1aP9htmt3FOTfADEge9fEE3MURnHBSn3B0Y2r0mzLuf
/xBVuTQTaIQZ7QyYmTkZjpBLBTpPu7FDKXolEeujnuWMwvcfxU/2BXRoZLYmQH67Dl2BCQnOaGnV
g1L99wYASX/DA1oq/v90y0mt4tHYoBMqwCx/rbdj3l/lLB26JdHAxdf3db2WpVkqW+wxcdGqNxMZ
fWBDrDLVD+rE4DqBW1YPr/XjIVGF0Nz7GifUzVEKKvHqVUbzBMQ4GO80Y36fqIWyT7vTcUi4K6Ha
Bydxavok2WMo9tUoUVaWstrqgNqzM+neOXAcn1engn04cxP0muG06/utONMTwZUDpv9QN/6bwVs4
KDFnEf21sjfznTfv44ngFvzhmXrmYJQUObORoH3w7Gi1qOAw3k4oexNNuH/94hx36uOaebprT7St
xUSV36UG0rVlw2RSLv7GWzEYELz2zFV2ohYm6YjMV06d/ihJ7to46tn9sM0SpYM1hxdjAVY8p5TS
pCVDCmvi4BRiW2OG2QykcEem07cjqBSviXtAwjsTiHWE+4eIx0naw/h+VTmnkpcqOH8O3/wI2guX
YW5ei2y6Thjiuxv8WAmHDeogGmPq+0mVyCet8qwHjsbc3uEHFbZjNkTNNFgKAKAVdgULcA9yt+lP
5+Z0Z8qV58WvhmNvxEnB2hJ9fBhX+FuClP1QWNvnsX1yS5X3P/hq3Ete3tkPaZQwJuFw1VBjNpq3
TYhXwXt2jnws2mUGs49+OyfPtHK/vhvr4rxcuJVmSPeuXSKMcLT/2GaP1IWuhUiRJFTlAm7cE61p
l79bNs2lBUzWgQTJls3GrO0po6UCLO4Pg8O3/5Xq4eoXRHZ0kov1v3OqR/FzQkeyrC8e4qGC3i1K
v98/NJawdh1AQmYT3xUwXfCLKolWVrhxhMS/otQpqHMAEmuE5Z4NFfNM5whnndOa61oEEO/F6/b/
1U9W5eC+aQwdsUdIpFi+4sIdygZbnlcHDPy7SchZKeBIdshfZw3K37WJ3vMbRnq7Ildm3a3+7MJN
NJ+9y881hKTf7e5rs+HoJB5UKrohSEenqwtBQU+WNpl7XtHey9ciO9n0JtM4KJBEz5u1MFIKPXr7
FQw1zmBsSVxlEZvLIBrmnarhbkaxOaxxVoRAV8qzbMjllHmE5HTrU0SKfKsBTgdyo3m7dSsQYAqS
wqQHXKyPhk4ztx5FTk/+cdvQT/0Ub76Jpxx/bVtWMNj9+MsuV9cEgRz/05rQXfGjrCsc3xKfYGnT
aZEJ3QLZAR3jEandDtcnkiJ4BP/1kBonD6pNEx3Isp1UOf/932LtXvmZeET7dN4hph8SYFHcoolE
AhUhCCvEC9DZZD4xqWp2Gh3HbQhNinmYtsoti/w587OMTx6fJFkoIsl2+/Qo14RQ7Bm13yfimdZN
PEUPi+fgwabBNIajomSoWCJX7k/kHlTXIQpLHiQgHGBpvs8pWFWH4+Fez/HPfOwyPFzA0DOUMZ49
bs9+M7lvNJjO8ujIbWPoFDNRQv1nJJHra/3HXnJXMQgUh1zR1ZsrpNpWMFAcSbb2Ru9PUstyVczC
pSylUkvP83JvnsZjaczWmJh6FvtryyvshBGayc5XTxBymjQ2RQrA8Xfh2fqp/ndshg9VlCpgKk4I
BMY/ojr7hpAlrQUcXUocsiVuq+QMQ7Dx+Lptd0qp0Mf+/asZ6hJ9P730zucostzgxw0ORfWMmR0m
uQDjCC2geGqxOYepp+4wpUeCeRbxjHJ/sCq11lTomfyrqgabjzte2D4ExEI/WzoTqoR0DYnTZZeE
PYYzCCAMZXAlriZByZ1TNeoRevXwVI3QvJQsf79c9zSccKP/o3M+LF4Ygd22XYnpUCq4EbUd4DGy
OQliboYsLJZUYlu7+qDssgDuCgBFkWKusBzPxpiYZzQsNj00e/Bp23MP1ddaw6P9ggQMqQgiwfrt
UbyoaVzD8I/s6IXQNXIPpcF/y5l/RSXjebV5SkQG0OswIsFbm6koDRua4EXlqmU/VLDxuTKKA4U4
Vx2ZgsnYWCWasvKU0uDtB8QiWZ1QaCQF9CAwkCW46+Zga7MUtqQ9wxc08C5OKZalgjY4BbnbdLhS
xPzxrxDGVN5jq4ZDjaqINWv+amZfHB7ePOLeK/2DQsivr18Tehs4LU2w8RtOHXOsbn9IkWdc+RTA
4m5QNuSXprTWHHSZYfBeyla/EPp+KEHAgEd5zzZigOS09Alx1sLuH8w1kO1KU34Zx5QGomk5Asyn
rxawnDzAZcqeHCM1ATlywnZFuqb2XNoRuYByehdif/G7aFoUycJV7VW8v523lo9bvH+1JoGpHFh0
4bIibLCRZwxROKUzqC09Zfio/QSD0hoAsngL4dDyXWYcqMCnSke8HJV6T+M3P/qNoJH53KiTBzTr
/7ZwPYCHoUDRjUupiROYqFVZERRXZJhJ+PBptvQMv3QT8Rw7dddYbS5aRy2NRlISRNXMDbscTGLu
hRHaFeyllctRUkJ2ciRcThBqhEWTwzXq4FLJM3LNCYLLXFuqzkGL26qcgCnAXpg7YMMe1lPhN6yt
i6+ahuQZfM6g1A4RWLKn9DIuWofqW2nVh51bCmSv8w7xOKhDpZb+0CvYCrSBoGbBs7BcFJ0m4Nus
LnpUWYxEE1DL4dyDRJFyiIqIGkm6mukYLvJSs5WVoilUhbjp8f0b3KtQ86XJXOZFFpfXE4VWo5a5
59PnUWDyOm2s3F2snQbOeesHmbnGHc7rQLivw6yjNLQ0YlnKDzvG1F7VxfbNUvyOWwFD04KyCz1g
W2QzcuHgoKDXOXkA0I1fdnLbw25En1fZLvdjw1OkPawO8Y6c6neKEXvGKtx49ngMx5XApstw6sHU
jYEOAkzLqAvAo+8oO+32UlyptKjmkogmk6qYwkNq6KZyAH3v4jISt+C3Ly0ae2gUgvKusNPRy6PN
CXKcQGhnMBeCvQY0nLqJerM6BWmst/yjh8dLU4lW82+s2agqQLZgBGdCCXbD/n8lGWI4jqiI4Q7s
wuK8Z6h87lYnXAaShAeFxAM2OPEwPzU33aoMYJ8mTcTXZeupnWxt9wCvxjRl10t6vLFW4xso9l4v
Sb1DbOQ2pI/JBQMHDp+oHVZabE3+nKOI4aihhzyNxldKxrLNFNmXefFRsRA/smo9JqlGHuAN0njL
mLZRtEql8GGj+tXWlXHtX7P4Y3K0cfbhjON106CHIbPHm8l99gHPIUpvYEIWe14/QdmwJKbYvoFl
5BkqY7ucZdACGp7rGlmFwKzc8xvJh4vPlS5vrUyc5CcdpHisDTO0KhztjR9HncvD2Os96C8DmJbG
7Kf1l3LkreB+n9qnf1xwA7nPU2Nohy8Y9Z5hitTJKK8Vfx2Huq9eG0qe2G+pTDmHhLeiu/0xq+Mm
gBFLgYDJXC8CS1u/0ZYcD8hgf6WAssTP8SDMXWEDtDa73M68j+nOri8H/EHc4cGlKk42Dsy9cuVX
1t0FwcPwroeAEL5IdRUN7PN9MEquWsJphxXE/wv5tb7wheSjqTVMxWg6emqQYDp6wgmkw92v5V2t
W4cFmH3Y+LC2xE6LQDfi4EOkUjsb/rN1tie7lmS8uz9IcD10uqrJwGbqWfmrxg9bRcC0gaOjNMF9
W2xpskQEPvlLFkh8XE8suBc27kHZ5+4i3Ok8dxt0ZGiblmXBc4UYMGR2pw4JKLCv3XX+M02Ds/kg
YsIZK9vraC+uw8zdXkcOWTdE99fDGip7A6GeIt4JMwhyZqCgL8uKi7q8je4ZPt2xvgIv/pOo4Vfc
Fm+uQHVAVvxdXBNxQWoNc3Eh+fP0WmHoVai68t5lMGgU8r4p+18fYdiONwJfJfoQHJUola44faLP
w0NgEaxaqYB1b2Sw83T+yRQoO98ceYe3TaZSCYgY6IWfUCjAnT/iDx4TVnhXjTrXaXzRwdfXPXjA
Q1AJ/MVONVei3CchNs2Ykbin6k9VpZuTdZGVUIbAxQ0SzKqs3Qu4CI4jsgpiu+UtwzuOjzv36ycZ
lUzDyJF1OeKyYguuE72HdEPZPZaRUf7LzTGIRuz1l8/tA+JSFRUJ72L/X6w7YN3U3H2T2GcL6G/8
aHpjtIWUDHLlMYvqr/abbV1Iad1npr2hmdd2xlRx0C104lyCmaAwZ8bb8nmb2tM1O8qERNUpFGSt
k4Qxw474fOAlJ+zAUueF4M2OtSCiaCt+GlXHTNFftVOAXg2VB5/5pYoYSlSF6qKSJ6Ei1XNjIP8A
xEdEjLueJajqdVSXohrFMVYllX6lrLGTyTVsnUaGhdjlOLDl7Z8ydaT2xXb8D28ZkCUu0KgaJfbg
UxDFt8cUBP+nuxQz6gGHHfEMWE7ToHf8AXk4oZYm5SWaZm7L5+1KfTtMJrLFoZ2Ifd6iZ6rOQuzw
9n6yXYfxQdagyPUhCSSte33wVvH2igCaD/Sa5vnI5IKTLPZaPo2v2P1N6IasLJkr+S5gnV125wRY
8Hdv2GjY3kJo4/i/q/5mtiJaFQv0pxD/yQi5o+AnwuWXZOtkbuqcKf0Pir7Vpck3kFOktx5VJf4q
esfWnmns8z63vVSDwKt16uaN2qLcpwi+PNa4DYZfo8x9JG+EPy0AxqxPJdD6HDJEz08ltNoQixn1
ZAmjdDwUiYuKGGQsIZMhPfkX1xaH50BBvde7nQSvlLSz9yc3sE39R5TccGhPMxrBK9BJ+UboCbxk
iohYCyfq1OSSJbLoB11TlS7QeW09hVs8PVN5IMaSCJkw5EYTd0ke/MmzBaLHjWexii83lm5Dinha
9ZkzU3DnBLB2IJ4tsMhlqpy2oIxeCBFpeehq1D0XdlQJfj93s+DV8UTdSO1PV1EN/ATbswcne03+
+wlKZIccEZxiqVbl4mFfa6WaTnntf8QStkG3ivWxuG7NoRwD52uayhMC+F0y8rnyTDdqjbpjYnVR
115gclisw6Uw0DZxx6Jm2FQZsNeYJXc2b/owrAA2rNcH7KOnESeIHqGpwIV/rFR3CusaJQd0klbW
E5egc+0uHQIfVSPOvvo3PwzGDZlVi45HW3LOs2ByuU+/H/cnZUMEr87KHm1pko2sVJrErKYBUTQV
DIDEpylqXB2wAkkSFMrUEheIr8oy5qnBPOt5mSitMJpxBcvtl+BKrLsmlLC5yw5od7q2JPm0TOLz
ptMmbxnp3ZPHRGG38eTkZ3BO3cbyXDVa0L4I8nfIRMoPi2ky3fsnwJ212hfJThbEpQUPR/vNhL2e
+qvtSmJL6c30uis2GhM1O99J1SNiUAS5hGPonFEZE+C2JwipMcZv5fIGb9mzT76uSmqgbdXLgQ/H
aDqwFz4nv26aUjG/Ey/6wJdPqA7xAOgH46k2FamMwyisVwyxq0C9zOffartuqALqm2JhITbo/RrF
JAkoXLuFOBB9WpqWyIyWOswUFc5DPhgOevnCKa8Xje9GtutcbpCdFJFgnStDKfkSOWLjP91jpeAN
vMsgxUS9uVB8f+tCDHJOD8NJcIYuyEmoBL3eYuq8qiR2nSt60SzlNoyPqjRSUKQ3FIVIpzxmRTbU
5GJtpevZ+iA0QEKHYU2FJJaVukvzPfFhA8Vnt+cO73dtRMruHkhM05eTG0KvmbyCYeXAYi/VNqdi
MTd5wDAgpegC98qIeGAe8Fei3k/sZwrYUSghW35lX1Ufd56pq7Ii6VgdPhh/cYDHltj6HVCqjEE+
Octsi0lZBbA8yeyVUQR0lZ2rzBYnjQ/pKNRDUqMCAykF76W615U3vRejNzTr3ZcHmkW5h3CBJ2KK
UCeH57y3/v7eqykg2x+dFfaslfoXtC6SQZu5Q6FSdsrTzcUv4UlqkrdZzYTe9GOZV4ZtwA0cBw/A
ymEpdhlymCW6SX+P0H1T3Do5QopW4JvDkPiAmLJipQx1k7MpSkMAYv6727mLYJ4EuyzXIG6ZJeF4
LfUGf9V7AJ0LdKbGaayDQy+s96wTc9/0R5n/IZEg4LnVh0pMUIDDhXj9wwJS3VlfxJB/f7diIh16
dZegp+Q0YJlUy738HuNHJN5viH8PuOAIrr23VWBIO+WIxTzpJT2TSKQIWEkKywkUTaFtiiRnov85
+yYJu7I9T3d85QO5yfKYnkfU0nu6LxSPRJBG3TzRYrDmjew77poI06G4bLg3bAl6+0q9ybOqQsH7
o39l982bN2B6kvQHyVCbo6oXLX8nWklTfOB4fx4A37ueBmmgF2oSeFQX0CU18mYB3H0PU/vxBCvJ
Pgmq3ev3PUv9PX7z8lrRnaPk8gBQjhAFIIkN2cPc6qiqf8ldpmNHWOk+tlMQwWkRiidNpe+LUcbi
YDnSu4G3Blf4oiG+yWISsh4X/jxhbxW9UgnsawIWVIjtN4N2YJJrIAnpZ1JX0Xneso4MsIK/haqL
EcRsZ3GJbG4qK0fnm1MXeDixdyWqoYDc6fmLAvSfXJBt2zfIqzQlLokC0FjmOEtW52L1C+wswvWI
AnQLVHd8Xa+G85COqKJCxyf7fKAyras1HVAPgnWcNjweCdayBelWFi1HaoP7Mz7pIFIGd05qg3FN
xFEr21YsZT/3uUNYy3E2qlz/ugWCazLvJcy8N4H2sR/l2k8gX7IiKT8v+IVy0M0n36qJLDFTOyIS
y2jW4Ft3tjJ7PE42/UEeA/f6oSBrwb7iB8rQ8SbQbFqBgs4mGVjq3QklKEup2v+pJgYOY7ecjhCL
Oqsw+aNW82idgaKLBbNX1MhLL5cyI5oZ8My7RgloMNgun+2q9XyOPLaLqGM40O0o1i6ddJv45cln
Kv6bBuajTWdaLtjdF36PRS1dmN+lJe8kQbg0QKgYz7kI0bi/C1ozwlpilHVIv8of17Gw3wCgUskg
0G5+XAWXKDyLFxfSucdQycecOPKpGvrpGUp8EwfWyvm/JD921xb3NX8JZYTY7xhD/s1JZGCN6Ciu
VlYJZ8gb25UOPlxr191EixtXSA3Bfm1itTTM1DHG9PojpGNeoFDlX9o5DtdpbCUoE1q53slvVAfJ
nYWEZ/q3EiHm2ho1OIk1OLPXuFby/gVkr5MRVArak6/Epcqa1ECr6Pex7E/LJHwwdnNRUC1cnKwd
fy2EwgFPeCyAPFvEtpo8OmQraNeuPiP8oV4X0HcGqDiusulWWC2uXM+5l83jeelKbvSJd3COuhVt
pm86PnMyNRshrPebhHKFn9jocld9tklSJtBBIrS1/kyXAhp4t50rTGYcD2vkIt7xheKz4eFXGt2u
XJhGfwBMsKXuVe348IGlBpDApZ3QqL/edPPnQFXPrmeQGgIrtIe2ld6CfVvJwWpVBhKkkBmE9Xd6
pdjK7QYN0u6AOfs4csUt5tRUTbKOdzBpRuIc5iE2SD9CHoAxkXZ2jEqIN+ZXaMsBNCV+RZQrsja/
O09OhCHWyvhfTzle5U+Dt7uBrg8FYE1XO+mKwNY5+KbPAdQWTzjL0bESR4oicwoHvx+dxBfZk/rC
X5y04xx09BNNKxNYn5jUy6v04dkAIVb4tyJsieWv3OPoKlWzckn0y01ITwfR0O4zbq2Asxdw64KA
JJWN1fAU2uIJmOUEOiLYtyI0+P306cuAMMdA6dt/i5d0FRQCaakVbrH9CoTw/JdrOEeS90C4h7eg
DtBQ8PhRlagIg4372qgTxqbdYRj1QNKsYNPhJNXO8BSZyyOIQEeqqHMpuX+eHuTc0oRwikCAJoL6
wR2rOzSVmgcVkDk6//mTsRbJdhmOiRYIPLnd0M1IlJa6lFZpsfcx/7rdjsFXY9exs63c/tUZ934c
3zasWS42VddklhPAu/DDzEkhbY6N7VcFgcDFkVzPR3NtI/pWby8mmEom4I4P5ptx4z5ts54xp1hc
wSUFg543KmQ6K6WuU+3dztUkmMn9UVCWPQQwQT7AkjEoEyOWdgtkmjRcycBSFcHYKKZq2ytwhHDJ
G2OgIMxvmY10wkIT/r7tN+NHXyw1D1Z/4cKGWX+RSblIjqyb/WmVixeulVIpLD50FA2lD8w1khIw
fV+bZUQqTttgDa+dMY41to/2uCijAzFq2s2PWe/56LNJHgv11V2GT2YlxJzINzf+tUhgc3Lh/zxT
m89+vAVfWmBIGK41QRSfuQvq0OmJn3MCbtZGqx1J4L7gNGZM7rbUuks8oJ0HgsDgHdxzH3WFg1hJ
FYFqHrPmnhoWQqyuhtvdOdOCeeSehYaY40L8g7Dk5IwX7tbCQOnSJaDny6t8/DXo1+9jk/TILlQx
Xxm+vruAnsGGeQPLu7SDtOZ7hWuO3A4+MFA1/z4IcH636MA4HYTQEG9BO0Xai5UxwBVFf9IPxH52
iCPW7nShwa5zqSSFbF6kx0uT4i70wDgXmgKHtt1IzwU/KSgjml8pkaWXz14k9WvCi2oY2lQoS+l1
76mlr8tEoJMof8deqWHRSRbW8632Ug+OgvtXjxWXR/wYSsus3kLmms9cJpPDvwKnSSgNyJPTi62u
izKSpnWPIhxAoMDGGnBCcNlUkSuX+8XMWq4yjWTAPoJ7NF/JTlqMPVNuZf1j9kpR1d4dYjXKg0DR
rEdeGx3CQdPhdNoTq9YBuoKtXqegJWG71+DNWyayN6an7RXutNaTt/2jL8U3i/C5TPi2neJH8mVp
MPz62qMyoR05J/SkfJFsOUuxs5tpguAEfEa76FoVc1Ic+ZCzbW4flNbRz2iI7d5QRjJxWTHw+p8F
cDX7VaZ2AFG0hW6wVO9lnEWNwocIESpsT77q6vhmmjOzd8nzsNpKC1MIOIiAL1BWOLJS9RUrf7S3
hMygW2rWkXpTu+o3fE8vf7hN7e1nv4Buo5UlM0l70Kp2GlrlsXmr7XioDwzfUCq2I/PR72cBZvMF
EnGn6zfiuQEAXHHWF2pGL25gkyKC/zEa+lQ0uCDN0K6yytg7yiVoH+HC/LSqroWGWh3Agsl8Ymle
OWzbfzGfI5fNi5BMGXeE2flWKLZq0FjIljOtHfxQ1E3t05RVf2+LTXDauAYO6TUS4/bNUBetcCbB
mYQ/QUzUX5ObD/NyWX0R3p9J9HIkMmk8NmS+U5c53nSHVwdJyjYr6rIAfuh6mOht/kcWCr3f6TtO
W9jq5mZcsrRwhPMPiqHUuUEDAYfAPG1DXk0i2vdcycjG3qbtqRXYa7titCsxVEp7cW5E8czp/JGS
AxZi4luBnHVE+PlMLiXrhEK0udMIVmQh8CWS0cvaExXp6SqfZ507/444OemkovbjI0KuAJnxvZH2
3wA0xgWJ3m+xv71r8yNsvcse69OWJ8hosbgotUARJhYWTlNefdKkNoYsDoTyTbwUwqk0DNSqgRw6
4diHFX5aKyQi5p+faeor2TmX6UKNaTny4RWWFFdiwvjfPg/6UFgOwWSWJTaeaSmLS3Eos4LrJO8M
Zx0pVHIIfgCHEn2Ir9SZe0zMBwCNkY7YQJEx5crdxs7Y6yzIalFxtD4xgax3ypy8TLsw52W4tYoy
zLmYTKSczUFtMC3fMbHoSzBxQx9bCtmMylnvmV6z/N+aOQDoD1NF9qqX5v1fL9QZ+KiV3wg5WNE6
qF5duBr00OGF1KQGjUzMH+7P1CCqBiZzDXaMDEBUl2Uof8HjYfNFh4DNBuIjzyzQdpoqzqxliWE2
VExqGnWE/rXDRwqd/0pmtJI7ZVRlQ1Okgsohw4rTmVaNsGHOgzcrj46yNQ42Ohzu3sH2Ua/xgEHR
e5C9u2bpVJUEnHcuYmYxK3SvQegwCiTj4PKW/UZnN0Ge2b1YcTFQeQWHxUX0ldtW4oLal8ltEsZX
JQ4hzn/dSBuHBYMUzj0wXlTO4dmiAqdEcHeoK/FfhQx7AMBOlw8CZSRG3W08LRIolIbKLLlOTvl8
ORBKTsGt9OO6lrD8t8YSlK1mWjhvfqUpFBFnbTKeKwPhBl9NqszjYMREZ1xi5+g+x5WMeIeF7ECs
sFuQDItSWyY4FNhx7zfaaIW5iRqY57ASG3wSURKjN6zm9wbt+6l4gSXnsO3DJ9gYx0AoBTvpVkdV
TueOwc1is8fsLbHBmdb9Ehl0qedF6ReSCYVObKfS4E3uxBrgmJYkeHXvPQdM2h92aqWsJ9XEX+l+
3V9M43kqCNSgXNZIfmFTND7AZG+DOHOioQcHcezMCFZj6CfbwKJNbdz+dvSR2QLjNcPCHyt2Wuns
xsbeTLkFImhbkI1n41k7YQkMdRG0O6m/5K6pbtt9sTM9p+CqNsgEui2+wJh0Zh9g+eyu8V4TlzXr
x6dAXj67OYRzQIt0NRU5Z+JeGdCueotOyGh7vhMvTHG+0ZF/D+SXX/KiOwhdC5SfhUhyR2VC4+Og
Pb4vsI5kHJO0jRLoAXKU4PNRafi7PUC8r3sY8nIyjAVR5+5V0Ofgqy7Tu3P+ePwsuBrq4IGE7vGk
YZW6KqR8RYX7RqDP/tePCmgl4XpNYkqvnru0/bjvndU3nNlnACyzfUND5Rknp1T3CR7moktaOp7S
ykUv8fBU5ysopBkX5PFLoJbMO43SOqDwjHu/rNLyLmux7A/qwxFhkuxbIhhOlhysXTrX2/TihRYg
hAoZeOvjBbrB6N8ahdqnXUQ0XSP62YI3+0US5pPyyWgQ1IVMmfAziIVINbIeMbcYc6X7GV2XUaIi
JPXXRHr8Hi8o5VJrlnuRK+vw1ORIYJTLgrvrTRc5VM0WMc36SoRJRjFd7Nb8IjmQtfdRi1m34JER
V3MzZTtj6FtyKpKtheK4Zx7whclZApLKSQ19os35tWq1qJZZnp47OVmgwfPTtXXASTQVTc4ayGXG
cAtxEEpeRkrx/bcT3eFdUhK9/ow54n4I33GryI7HruYRdKW/H8naqBkw0VljD+XIzNfW60b43OTV
IP5A35NQx5QWfLhZuGOx9ZgPH4g6XL3lJJfJjvCClOCISkBIihvtDoPyCqzcJWAP1qS5f0yJOoKm
EAC3Vm65/LHdgAbLCa57w9cE0DeA82/NniML8qocIphCid/8ryrZkJQdCkfuze2gDV+IUrR07VLr
oWZ6+1fwESVAderW3IvCC96XXv0SxrAaUN75mkp5dP9W4CX7RcqDpljF3ttmnLK3PyyGn7IluNMR
skmT2QPfXajzK+ZVrX3F5LYie3/prmT9soi/A2WeWwxCSxDBQpgP9AQtCbbJpyBdxkCueG00CRrD
fKCZHpMRQXyFCfghVeaM2khDuNkGnf6ACvYUbvOiwulbN05NBKQ++EexLQONCvUeIsRqxH1LCncQ
LbgYxSQdAOGGbOXGETIkhX7JdQE1AMdjvFUMz1lDYsS3ZOwP8xbS+XIJcftDXUW9QiVdJIxXyLwn
/kNdzRTeHmTxsMVSnS4+nMrPc9v/25VWTtD8JuyI6HzCBBmlBIQldVTgu3rwKl0uYN5GggVt4PfJ
65CDqGTIptlJiQm6fwvnGf6OUci8Y9RVqXs+tSPjFgONosMxYvUUQOdrrcuB8UGjiLzyDX2XMZyg
kxY9TG9OTvH/Q9IZldgoKhS4oEHeuV3p8OB36ESJpAUPEZHiRCln62Nu/8lMaNCI4vMfUoXh6KYJ
Jk+nTarnDzTUrD7PSj300kDRn6/C1sJXZkoDmeE9XC36OISxI8i4MBbwKEuNiMwwYQDF5hksrS1r
CDmd+/ImqXb8w0CEgpRgg5iCAolOU2QihhuPjMtytSTgBH1LAodNRvv6ASLsATw6YHceQYMwEv7p
9Yw6CTAfszizsyvV62YUIFBJhFlo+zjehC/aHGUNFHioi3InUS0YZbA794GKBWcWMZJKRFuhpVqP
+xDxI8qMUULBZEryERnYSgieW4EmQHwys5cxqZP9Z0xbJLv4YZL66VLExdWi7aHaY4J362wXhR2q
44qb3C0jK571GtAT4sm12HSwh3Q/JBePt8mfGN+2GlJL1qJQJAfnjrRxKPQSkf5p4+dL7dgGqayH
zIrfvcGcXc/VKKGB5jKK71OrkeqFx7tkCXvhJBQ2TjTsas25w1GbpQlCL2mmPt7Rd7QzcTPIscbY
8LdiP1qRG/XhpQ1mPeFqqMqJ17JonCPP14pPUFTFS/Z63CDWEHUsEf1c7h3dYcQOeH36sdSzJXAt
0mKGuJlBlSwcFKJqnKDwYC1uNzil3U3OinXY+2gPDShUvN6G0AgaUm5MvNmZBuInCvKnlKLlHCRK
0oSj4jsjDZIZUJhRjNtMACTkLCf3JHUEp8SAMqQ51xd6Ey+iSW9L8WbPcumqPbDlek42dqRWrfmV
d/wYqxzrFanElKIOVXgGohIWyMflYZZ/vYsmoMtuzPEUBSPluFcshHTsxOlrWBy6sLeZ067nevs2
0nZBX+yfw2zN8s2cWvT32AXxEOGT/k45cN+pJZ0Yz3nJfrD1++7+Rohjlu33pB4ZGheiA8Rf3p18
NW+Hl/VzkimxFyhbjglgcW6isTdlWHX4wuM/u5cw4CSz+kCy/QvwuqNUr/IjniShvk3YWJISYMHK
S37XY8vIWfbKEiPtUcrQ05iQ2zp5zEFXjGWJm7rTqeAw6RZ+2MXkvmU40DPs8BqUr9Hsx/0VUWnc
EJ7FpBRvMYCun+ruzCLjh2DK43Y9YCyebNo8r9aeorlG64U5rS5YtvegynhkKK60psZDXv94Bmw0
NKJed86pog00s+QcjlYA+C4xoSLapQWSLRbFA3dKEOlUu1NNuX8K+w223fvoCz9uweLEtiRno4hR
LESM4ugZLWQGTfMfFPpPl+n7i8f7PNiP79N8ei/541M44Zv1WjT3RAHwWOO1cyydONng4mGFzutT
o+CrM0Y8PO7iLqn/LBfmEmeXGHTdI4kp4LvH1XAkdiPNXpTOkm9DsQuxRzo1mQ9cMoKZ5bGV+ss+
2EUpSa4svHqLhiljcePMmkYEFYQMu7rXuv2A2K6Pk1ySnxITgPjQd5F5gXyn2qhgUKeVfj4/lPde
5gvxSLNX5y5KeXV+7kucm+F2OoB1zLUDhCryw1uw0szPeFuaUgomyRaS+4FBaGE9S2lo0v+pgYuF
38V2NDC1WjqxmU3PyU3usdnSi1nOpTbVSMA8ETZHoVchS53Mbopjo0QZUuVjoEHgArATubEu0tfn
shDqAnS8cyhMQAZBsbQ2WDYkFUylzhArM3pCom0GNdkEtQ15mEMcJti/CKv4YO/ITOqzVcjBBGAH
hGPq6HHwxXt/oqsCcOskBZtdflAfUVNZbD4GJ+tXJsVqad2S4J+q6m/FADBW/Hys6xDAWDxVsgfK
JMke9bxK7b8C+APeeFAfeA5LkBQ6p9I/fUcpxpYidCk4Ds73Gj61lxH+HKmVPLJouTN44UGQ0SGN
4lffCcyNRDyxSJwyBN3NH3ZmFUv1uAct+aQaeKQ7lJBJ2f87uXznuz1Div+34irSCgS8ML4QNcxx
K0fht0ggmsBLxeSzK7YCMnaQYJzyUouctoN66yPucexnliMn3lnMPD6BBEtyyYCIRaSquN4pFi5r
MeUFAlmkHJEN0a1YYKgp4Ed6xH1ul6zz+VbGNApB5l9E3WgIzY1DNpaT5ZF5Qz1Piws2QzI4ywYk
QqrTRdHK9fHgMesC0KuVbX1VwubPO7AmIyDDrm3mq5olv3r7Q1OI1zu8UAKUB+ptSsuaZtCDmtqn
ve1J+4VyUHAz1lSbBtqYStSnCcswn77qpW0hjCcvdusu76V+9m66VQ/mtwx2qqRcs0uW6pEGoFSr
0gT37DvPMolC2K3ygfrUajSopAv/c2dm7IvYBlUxctzB4zBWL++Xijl82HASWFGxjoS//IqDMzN8
EmDp4sObRb/aCxKENSeQEJPL7f9aKA2NMYQVzGfi+VLdLzYM9Lm3XYFHvqc7UlTGnEPR0AXBzqBe
AxAfcfl1DOrsvdRwYuhXbOYMht6OX7d38tK3oEBQbDJKI9de82xmH3iM0BGaUsj9luyWbsMZ8uQt
tTKoH4g47PvwK4BqG79h+uiTd2jb5+NAD9wY+5457jZKhwpaAVfO2a3m3DXnu+CUCguQKa4pxBG4
GTF5NjZ7BwpLn72TGkojm/YwrtHqIHND5j9D8lMLvyCxva/eJ7WXV6PtjAuyDZhQpRWiBSwXDiwO
64zFfFi7YALTu5EUCvthqCYM7eYHRhw7nhKCwt3hh66qJeSXfwfcW9XCdVNJ1upDtc2nX2nZAcYn
J1gpaerDZF0jrsJhjoO7pWED5Uc/qxYkHdNRXRP9WsAP16a46UXz/5oxVicX2UDLRz1/JhwSpo38
U8Xkp0OaTsvnvVFfToTqeYVQLFUrC0TCtxKR/ci1G+kFpq5qSxQfJpszKittM/SaPF5GTYHhqaK0
4q3tAVQCqcd82iWjF2PsqhReLVR7ingDyc0UOUz/7jSWMq67pbR4L0TmIYIjDc3PCk9v4V1XdWTK
WuExqv79QNhINVQKdekl/0dwJgxOqjDsmXKp7trm2EWf8O4dSXUU9aozTAnDM8QNLWWiQS8ohUwB
w7xg37Gqayu3ttbRunWv8BPnjfePGj369pxBIBb05P2k2jpBg3HtUkuEJlzZee6i4jsnGiZa7T5q
GgZyAE2MYvcGAWk7RrLw+jCnfn/QP6SsN8PhDvmcHCImbucblnf6Hv0xz1hy9pchGiO9/wiN4RAu
Y5I7hZKacz2h7qBMGo6odD0vozt7bQiGecIGPK2yyIaeyuC8OUyS6+EapT0yIWconaWFPQL+lSIz
hUewaI0Wry6rmB4Bf8+ppKAMv76W9u57KWdzq5SM5KYWehSCuOKSAXL57S8QH8sl6FRvtqDWl4TP
nxRKibsCDgOHHX5AqWc2tTmtMWZBeCC7B9EGbyL9nuJI5XTrW2xsqKNT32hQBWZONBgwq92w7Wif
ROntSH6vU9SdNq3R3/RzZyjvnygVMsHO14dUsksLnOsCKrmZpp4rc5cKCRzh3ih6whif+xyNCOMB
2jnfItMd8uUm7bfKEuOq236Cr27VJe97S1btAy9tCFpn9hZ1Tj4dUq2WdUPtJZxrrBAr6/d73UdG
KPNY5jM6NHgAyX/WBHuxDVEKt1boxFKhOMvSrRYkerzyVPygBoLSvMRv7U7/0qk1BmUzPmOWxQR9
YnMgVOmH6iejnONOkqTwzXoH/koF7ZtcwR/dI6yig/79XKdNUG2KYEK7m1v3Jwkr8ua9uvFpKueA
Nu/BNLbu0avopbaupwV0THe9jIA7iMkwGf3Cs6djV6+BeYU/XjWXjXYss34aDzlRUbfIZtQqCU2H
LD/YrzIe5bxGr+ToSF5JH177sOY3W0BujiRPxbLALvMYOZ5OAVRfy6rhdsJHQ4U5EG32Pt3ZbsjP
uwv8k0sEZNS7qzM/HTe6GqFuWBgXf91oiLJSGZQQKQTVG8dmq7UfKAtLjyXWZNokdwlskpLUkDMH
1VqTlUY3pwKZIx8ppeZuE/UNRRxZ1pU2HvbysBEBeMwRPKXrPAJCL/APzHFJT4vdXwmkjB7Tu84F
SlRbDkSYYouMhCwf6bFRmd8/PBj2H8z3NzapMaZBwjqZEp11CuLSxUXE6HDKvX3G+pKMMnBIT1El
jvn/WXJy6HBg/IUFgARLzrjSS21WET6ufUWKKqzRnxiLO8DrG98r/8CD1q5I3b6bnGzz32A7PUaq
Kre/D9i9KWWJ/jtxlsDcnN6Sl5DAS6PctlsAC781ypdaixrlo+uHSCIELt4u2I9fknDYZnySKvx5
tmz6PQvaBXkU2OSlKOZ63dYecdTuuANs+yE5SykNajUYiHpLKmdRMb0bRkgCXr2VaatozNFO6aDL
604p3isqmdyB0qBfbPzLBH6ckttdwnsx6neIOktWARSEibW4QzVTWNnKvmdk8ZYVfxVKWRvW/Soa
0uTvVJC1tb0EP/ty9aCCozWoUUW6YexoyewMMXwGMediAOTRnuYgieUz8mmdqhFwHPoXEpKtGBVJ
UmCgFnwSpHvsR3trWNsXPcDxFWFi5NDvtXsXBChw0HHHsZ18xqkMLHPtQJBYm89x3UpLpe1SI9xx
Z8KoUucA9Dizo1qG4LIl8HpGqEhITkPMfpnJdezA5u5aeKyMUjMy7SH42Qo/0mnD48pBcJ5/ygcB
b7WgJM9Ver58nW7eeHI7cLAF+bgdy3JjjHzsHiIoD+i3BTlxl4FfwcqTJ3rMDZRzC1E1033hHU2b
V+D+kZ9LhjF839WJTguTsV1vfClcjyG42fWN08H4gJUjFj4RT/EPzudJa2qzFE8fp/HbKc6F9N6b
mCjNB+Wm3gGK5GZSOl2nUeV0ECKNGl+K/wOu0Dl601Kaw2IPGlWVuIQhrjPwLEXIt+UIKOD3tz5g
LdmtS9baNF1gcTiQ33JioaAy6+bUv/+3rz0Y990xbjGERpoPR2ntpUhdkWkF65VNgGQORzT4Z43z
C4zBBA9o2+dyCn8XNbaYAvc24+mEY8ho4yOvxpyaxYuTrDUGqNwG/c4r/n5lhGII8loUImR8+SnH
AyYDOvgPMZOuNGDC5eBn0ekBONLlHqX6pO0LX5IEwhUrgu8t9NttSMoK8KsyA9bjUefcVZ8phbjL
S/k9Q5iDWYQT7UlgHSgSV5wlAJFjKKfStg9p7jzOeqgWKOe3Qj8fRRjT55XCjSm1RczvtEvPVym0
Dyz8cmMI/itRC63L4gPjWjkzFu8ZROH15tRTYsPnDmRElLgqMv/XidQkq8MbCHA4RI5al45CpnL6
QUQTVP4zRs7pED/7Zj0X4F2BwTlqz7QNv88olycjA7u5UVmSo5a5RvYub8JB0VAUF27NFQc2JlSt
s+AwihBJziFd3GHegIviMB+X5DexZHeUSJhzCgQCUMOC0G4KTlIf3DWe5tGp/Uf7soh3tWDBzGau
qGlxZRPAagbUr2OU24joTQSGhAo1ElZp0GgJ7nZBruPo/eqAGY+nH0+2gnDk7t7zJ05UcSGGwzN4
ZiQCXaulCLPxBk2fPmytHFTcdbvRwRKwZwVXQNeVP+j6MVDtrRG54y+17MO6KVjKDP/wKT61IH7k
JPvujz5gq8B3VG/M9QzxYWSLUBJl1+Lj/1/x4DAr4vLZ7hV4HQ9CQ3dswts2fBZxJ88kqlXWAg3J
lKZ/ROHo/PXjt8quc7G9MR32hiR3cJ36hxgp2NXRb2w4YMyh/X1FsgLRboIJOryTf7toekbktgOQ
jk5fBQbhfce5qkNKO+rI2iOwlGSx/7pWBOf55iSbNKrBbYQ6oJLfmGRCCocs80m+h2eZoD7NwBJR
Qvu54NfiODNMDJ3sl0IgFJgvudjPvwlzxLLd9EwH9vN1/fE1g8DIgvOo16yux60G4L94R03241km
hqrEm6UzWbeCxU1kYGe4MRfK/NTZmNLvnGYh+7I/pqMqohWQ0Am5PqHhEApaJfpytjwgRgrkgiDt
MDGApWiwzeq/StnyNwT3MIDQOLUmfiuHzt1lNSVW7YtLOx9bHTSwTQ7Li8efLgc5zka7Ak/dM5wc
9rIsCquiXpsF+gQMBgWLnEshdhbOjIXv/I3ViEmTkA7hHXZv5rqoIZQA14BnaoRbm0/hTde6U3V5
WHNrYEsQ+fzFdGKvmj3v0rNCH7DxnwzNvulQtuPB0eP91xwvkJc0Za+DpdQfxDqKyKoG1sg2pvb/
atX5X1g8k1r/ahU+fYI9nivlaIhG1WezGxvpcObirJ18OJIulmAQjXGr9C4zC+S5CjzIj+XHPpMn
o9gRgNk8DgHoE3Tv1HLJsBwB0ihmABdUIKFQfIyUD75aGCRvlyRQX9wsondDsHaYz1be8ydsfkvY
w148CYA/Cm1KHVztHn1cez15dgY5NBb9Jd6FYStXPT3zAhNC9ew+lKzMeffB7bJNRPYoiLyTugEd
mX1SAR1qOT3seYepY51iQpp/kbigq2jbuZ1xoPF1xeJ/7NHZfqFFSFV5Irmm+X7ZTOsndhw37xvx
mbILqEpVQBz6F1kD1tjXBuIaSdm+lP0wH0yBYyfOtfe4QPmetdBdoYthmFQeE2EmZvQ1DKBrW3Th
s8fDxc9DsiM/E6uapmdOErPLVNYi6rLnSIuPXomyjv1KzZ8j3eqwCRsyBgLbZuoRmNPPiDU4x1o1
UwXZRYNtC6C7ET3ABFp8KSGWHR/cqwcBwvyXBlZ89D/WtLfkTvQCe7HMr+43GgZKAO8ERyvir9Ds
DfS/Kn3iGZDqQn6ArtBXMpPoT7NA3mTxqrtNRNN+hgiTahpFSITgLpt/7YE0jSVe0Cm13SOctHSG
T+Q77KBRG1j1CTopVmBj9Cs4CT1XsEPGLXv7rwOeTZET875YCj13D5Surjk/e1gVM6svcweGvBhO
H0GmWc0hBeF9wnJOECjHoGwpBW9QxqojPtUUpN35a04ao6O1deVXh8OIcUw28yKeWkDNh3xqWtp4
12ZP81wj2EFVnNsb9Ab1Anb9ZSoTq/+bu+hQBf/XlR9J0VPDU2Vtxogi9NMFXwR6fYcHe8fNB8En
nue5E3gcO8h7IEKrvd+GkEIEX42xljojrG9LZwbwfS8/GLIVLy0xSjW8t6S2xk1vvvvtvwSkmcPT
qIP7hA/wL7YF+v7GqPKG52i3aA5EA8vRJg8krSUxdlSl/EexmDU6fDMFCe0RyoHFvLLvcI1IBX9w
Ij7+BtdNCuNlQGbjCJDeHhxyWgsgGKJnwniooUn/ZmEgONUblL2OQ5mBVtqLVdfIXztvShzxiDR/
KR10Od2ViAvSMUsP3IpuxPWsG4OnSEg82HjxD7u+oc5XwU5uyzOpx+h7oLKCol2iTGqLvdEHHTcM
Z1ZleFNItjDxj31msH2T8cJLvuKssEpg88iCmEbuarOkA/ku7kF9dA+ZTLA070YH9rpmXXEui6Ej
2D1qpDMYxfRLNw7Wc0eHR/CdGZdXItCjaAgGZUJEL12EBGSlaa0T+Xq0jejjD4W60qjuZB6tKVv4
8NWfHjjX2JoWxQ1engVyPvlXVitCq6frgl90YFl+J9l1wgKKhVcar/T8HN1ZBTcTdGCJSWzULaxS
f5/l/gVp9ndfM0qg/r29lm4vDvCreR8OzrgBsKCHKxKxi2z78KPUSzfkGon/ttF11XGIN0cOYmxM
ENyFFrw5oZpFxI/R8L8M+WHK+6vS0FLtewySpvb6spUwZuSXlEsRrXmxGLUnn92Fs2atQBkj2hjD
RIRR4m21RESgEhG1pmU64a3yI+omoZ1VxQj558R+gXVIUsg9DwTkYLMdkbNHVDVYe09Lg/wy549k
fEz/idL1R2UPJRWpJHEugLnKzK9At8TEHR6fAlmfkHurRGK2VpNQAK1fOyyy8p59GTcrZqm65WIx
lUldZf/ZL7jhf4WUXsG8Ij8jeI/X4QImwz16DP3EiBMnn62+rsKipIW86Jpem4zhjAgMNqCx1yKN
Q7jjjsEyrr9fWqBVNLFQq1rYCUekZ2S3faRr1nsJRCaUEXObYJVD5qdABpv+ClBDK7FpxyHTJvVm
SGu09gPuqliZVidOl1BaSEIobHFhO+oXhrIpDEwZHfUcVQ2jYi/oc8ktl93DO7D7qGZouASSzPWM
vuuLR+hcyV1aC3ZWxDyVLg9ryNw3Z4VjSyIMyVev3Sz+BRZhd1VYETLwqKGc47wMuoWXI/DpMTl7
Owu37Z8A08Z/lGr7DVCsgRGEutw55P0H7/th76zxYPyxcNzBM5W4G/CCC57djUOrZeZpX+0EQLK8
wMxGjbK2SSciI1lelvYV/m+1LyIECCGo2bwH8QtBY6pD+PxVroYmFjyxyIO0LSRmAF0Bd6ZOQqq3
rBiGOGF9dMa9t9SqSHLyOe7FqF5mjhLXdYzfG6QvZvbuU4+Ilmq5KeXGa41YkndSqmTM09inb7CH
pEH+2jtCvLl3AmFbUWIC8ADQRTQGQCCpyhjQDfKUYqN9Nq/mb1F6WRFgasw6H5ZTPPEfRy9/TNT0
gZ9PCu+Y27QtTcURN7W7YiC1WJ92MBqn2FjllJdfd/pSTHQFYO2B36PGMhtoV6GZvipJP6qbTPuF
PXYKDmltSPBoaW7hXN3F5S+faCSNWjZtQaTiw2y3nOJQHK4UxEJbZ5fE+Xd+ynSlsZbQVesWZ8yU
1e2UsVZYSN+MiIvNRKumWIZXeNRZziY1cJStn7J1dfRT2yONDrWaJRlEFLfP7dg1GtUGc6YXDLSC
Q/2tDs2kdDX+2BUTDN87dMzBN/51BynmcwQamOCY0Rg1fhreixHoxS/p3f4CPjahhvnNT8TVMStQ
sGeFK9QQV/ucsz/0qFdAaLl2NXIHnD6b6mUl74PSu300mq4+2L0zIhMR4ssyQNkxX5HRigqRG6Me
ejN2eT3xcAJdV0bGhMLARI40HwY6x29SogthGbwGKKYHwV54MVA/Z0i7wwMDBf6tWW89Z6dMOfsi
jjGb0jqJECvN+gyvU8EBpHFwp8Mamuq3Av7Q4EpnFERItex0ujWMoGxShQMbdCd7sxYluu/ucT+x
aCmzfHMXD42XkAJ1+t+XTGPY+xq0H0h+B0v6jj7T6Yp6irNTCmiQXbr8WAWIvGoy134xFdrd3std
aNZxz1RWp1IPQRtAEnDSOpCtPvtMdnl5e3YxAqxBgUx1q4E19YKKR4JqKCGfvWAXniRayV4dJq2t
oHOX1/OFjDSsIYgAFNaopQVCQUqw7yj9DfYYIerOu/pCaXZIp84c0E6OM0dfghl0A//FLW2RGf0g
UhC3Peefy/ZsMK069EjhIn8QHBfNKkCh0HVgyS4GZnCrhrMBjYvi03aCGsOHTbUL+cDK+Dm4EHUx
o2xPw8s8a13sGXU33KQHCwjSgoXElsWJmi3MD5KNLDrIP6cIfIqGdt06XG48osBM0JX7uknb+UqM
Od2WdTblu65fqktCvR77yMzWl6kDIikL0JLtjBsTpYacYC4zXheceSqML0vVxjk7D3gXZxDLLMHq
xKixVe8LclogxYb58pfeHaka9BrxbiihTXv2Xdw8OKmuf0l0XF0YuI+EV7FLJ/zCnDc29b+tyi6h
5Ne9rWy7CJV6SAtKSGmOMtlnl7/5vi17V3qoEnXYCX0HLrO2qmJQYY9mmDtu7GBdt0l7jWqvoY+P
ljjfb9M8SX1TDmom+1Dc8cu6+kWFQpYiV8IUFBFq+FlnUAoVY9pclLu37soBIuLgeFm1gCryIM5v
2BlRNCf8q2gZFKicErWpLEhRK71bSa5Lm0ufSNkxMOWKJqZ3f6D3ffezspkv+XCaKLvNssUpTq18
Nncvj18f3c/WqZnCeHDvHYsAViPocLo65jO2dHHtsf7bkHI3T+TaC1CzdpzNaNLOJQn7OlBYyhRR
cCN3nKtx4pm8e1ebHxNaZIQUcDn2R775clTZzJj5mgJ1sJmiSNrpKcm3VFCQjbsh1c89CsgmVgUK
VV35jpKAa6IGI2A4Y/V8iHuVuST83jNA1vojkYEJeMYTXedGatNwhnsBNNA78SBRzD78tBS80FkF
BM9TNr3ni7763Lh36I9Nc+5qEMNDuEqJKz3vA4avlCODORbrsYjzNL8wqpfO/wSed9gk2glRNfuR
akb5DSBLQt0uZqMSsiuS/tzKRt95TEFCZ/oI6E9FCxOAL6f0wtLB7Citm1Diob+DG6WvdYJp/nxS
6LO4hYiLV6BPglt+wpUrmv2POp8ez6NAjuMu/LX2IEEGkE4vhCgt3i7NNbvZnCBzhOLMYFFLBmZ7
XQ5Hym7r8jMiSDPREFjNqlljlp3TxMBL55Dj1ap20KSRv4iqa1KP60E7+tHB24HfUy0Xkf98X+hQ
VMbhmWEdk25tdDaoGKRaCIcFN5EkRbiovfOmoLoUM3Jh+A84xB6owxKbh4ECngDmwuPciDl8geV1
fp3qySUYZC7TGe16hHAqWyKVNgWPrIPb2HjIS5G/F/AtvR2MD+MSDo5NII5Jgtc/ZXyaA4hEfg2/
MFmPxQ57GNeL3RVewf1HjV4mnYCcYutrsciniGWKvLmaHjB9Wuh+yt4BNPWkWQfkzqdakM7XCdGX
RGy2vALKYo3s0/8kfZySW2zvgoY/hE2dK3YUb0kXij7iKWawNShfy6QuwYUKnwON3i5Q7l+z8uce
2VgLLMmkUof7U2zmiCSrLPEW4H8w14YBQsOHAhTK3tDDabW2+88rIq7p1ZYnIfSnFjy8+uBYeLEW
VQjyqa3lhVrRcQME0HNeCeFLBPumZ9ajZnsqLK6id6lCzHjODP7o1T2Hs5odQ7lTOgq+r+cIRZ4j
HwO1sAhqAfunn7iUANDzCPJHwZY1SbvlpdZj/TBlp4PbDEdw9nM7aIo5kmSmcN9QrmJg8u5cnqwr
xJNd4zT5IY58yh+5KaoSBUPUlpElq9F0/TLY7o4SwvyzENIb+JihaW17avcIpVvvGcxZy0L/1hIw
yNFe3Zi8E4FOigN05Hvlp4KdFxCM65NijxqTQOkKTn4x7dTucTNHlkI5dXN0quLif6/6TCmF17lT
6EKYnUrlCaJFEnJXKovTA/lVp0T1zBwrr31FYa9PNBaOtAXoTP5FVJXg7IHBXhw6T0mOooCXNl3G
SdjvLuHguXs4Ol63F97YHpsM6GWZuAOnxTQ1ET//XaEmNSPktWuMusBUWd97fi8KlYZTqmJ84eKt
ZGp+yFcpGGrRddEDIM3S++AHrFYE+5B37cuuxr+zLi/h+wdp6nMmv+mV394qs3d2wgYXR+L51Dww
msu2hLLrrKrObKcAkH6u3U0UnhpX6PtOyEhFkliZf6Z6P21qqpo6hgfcii+ChYA6TjsS0lfkeIBW
y3gQV6t67Rvv9yI0yDxCP0+CGqkO9kwIMowuSXt08PvtV4A3U106pO0qy/C8XftvifTH1FYMXW93
/wgBmpIyN+uQ7NhZpvuOONTD2muM1Bv2NDQz57rXnOWivGYep+SltwHSWu+cuRkiTqDfn3ayZCCv
LJAmKjWrH3Aj6uvPZWOD4z0v1GXxHkAYRIs6spDRD3CTGJSEmnkcSW+rHaA0CoU9pmNhs44dT350
FwnS6W8yXhOJgSKUkIBCVu3KhHybDwWXGsGYQCTdQTCMB1dwShIoNPnI9jtiySvgxVtnG1VDyezU
0DPykZOSIxqkscG649F2hcP2xkVweShoxa1aEV048ixf9Q2nzIpyewNgn5v+wnop7PWPJolt5OY3
zTrmup4yktwcq/B5J3b30ie+Lho5bXHKU8IIP5HTgTpkaXYpZlBD3MVFYyaeWZN59h9zGEOfHu35
Inu4ujaP7grDJCdIncCpCgARDWp0R03sZCVQNcsyFPUR4EArecrEAXMgGiKQ1ipGwHHnl2R9syDD
idzLB5XObhreoxMq2MEP1YA2kcBzXYajMxXjj9ykiWi6r9IeY/zX+MKML5Uh8W3UZN+2Uf0o7Blq
WGVVwrO0uy06zKsUdkBSZYSmwPKOho7SaAlheO9R+/KHUZ5q8vImP1CrFAUoxHvvCLwIgNYYh8Ge
/8rnMGHIDak3BXvFTTTDE+1vkSdAUIYnb5eqv/obDE6CWDLah07H6PFWtN+c4x1MDirvg6Z902sY
Hs/oC6u7HzzdoROznv2IjWLZraOnWxh/TKa4hMkpjWmZg0e4qrFcSjFZ3ZZIQoGC2aAL7HgBy2Zr
CCtQoVcxFzSkTzuP47NHdSh2ncipIQ2JMMAJwbYsbI00jWpUMBCbL3XaWf9vYCd/lp+lWcdhtuII
XbQ2SEetVRIpZgerpL1/PWsha2LH2tvenKBabREovvAkfO+rTHBwfyvBGpa6pbA1azE+YBLd16IC
ZhC3WOP4lJwSWS97D5YQuaF+FbJYOlVWjUg5245LHW89m9Mlvm6PvIFAbBWmzS6vjByhbF2YW8Aw
jTcGvk5GuxUXbDddahCW1LE3f8exmyyLBvaJTh0TIFYGmiyllcPd5H9FQKN2Q9FX7c+REwsiHnmZ
v42jYY5Jmoy7Pkg8vQoTdv/MiQvslijy8E7qcDQ5T+SBtrr30hIyGqTZ9bLNHROJhwCQkLukzQUq
ivckvwyqfGVjCc3vp3bsJv8wgR4Xm3gdTsjeAqoFMQT/oPL5Z9zXwa1fjoSG9AXvAxQD+TiJv5Ia
pcsi06jgf5y1vnNuUf3HrQ10kLbM22d74GWzXXyk79CnUOhb/pekuMnvMxZNHxT1v9wtifL+eS/j
MuDOVZ2D5X6c1531IJ6h+gLb7FL5BABwJ2fuJwFvNUFDn6yrZPeklaIrWSC3vamp1ivCwz4l7555
N05ASEysH2XTIO62JNEsDcUaRT7jWBfjArlqQiCDM/v9N28lSl7UljLvmmrwdUax+LbO2c/BvgaP
5lU+0wxX/tdDAAY+RY+rd0igOVYwF6DXj/Oeg+EHdUegaBze4dKG62CZZZCKy2ItDbthx3yw+7Tn
OKudtmr+LBu6YoX8y6CRiH+USkN2t1DYvnXPjOhdG1Dk1G9C9WyvBHBJIEdTP89sWyKx2ozbSmkJ
NLEOyLXW0XwlT0HC7WaV5E+Sy1PdCRaKKPFGkQthSWXq3b/0Cl7BoC/Z2xu6E6f+0kz4nBFIHXse
VunztrTlXj+7LNtC0snug6z5as01mmDFnaToaShNIvbNBDOUiZzTvS9x2pXjVOlexGaBoMKc3LlQ
8808Ser+I9uA0z9mGkcG/e1cWPBf7PeY/HW8uimPtMYYZOFbZuHXA0SaB0gsW4YHgm0R1fXht1F+
XxFGGThFkrSJwFUWqLrWyEqx1lCerJd+mobsRgV0f8QLG7qLaiUGne6s+dzj0sGMN43R0JSwq5V6
a6lcRWWp36WsuHmiwcnWH3OmsSmWxicBuKCGLi4aHTXjO5LTjGWM9TTsYkbpynipPQ0gvSL+4/d7
/RcAMAf0yZNGK7+84HDE/je8KjPieDvmbxFt7JIZJpUHANns0FoAF9rrLGJ+lKEpstfXzsujCV0B
mTTzYqzqw/FXDuW30DWjvtxK3ESSMMtbg/DRTRxg9lLPoRGf/N6hRkRB5K9ghlKN2JxHN6OCSjTv
E8H1TtXqYK/2NjVH46dfF8S0sxJi3lyIvtGQPth8yQwUe+GQtuyiu0G/TppySc8vHf18puGZTEOM
UUe/fbtp7COp7so5VLAO0NMKtY6IbT8VcYVc6yZZEWW8CO0BqXpGUDiyua/iuKgXnyEWrW0dpZqF
8MlBuP7TEJMLE8+mYF4Yg8b2f1E2vMCwrFd2FtOR7C9ARGfsyxSpVahcfYY8H2702bhS7dRW0TGd
s/i1GI1VDPqeGAhGY6hPcqSCutQ54LnfFhxB3PhU1ymZqcEfmDvY4kQX5gws+dayToi0slk1qIq+
90WX4GbHzO333Uvs9HOhOwTlcaucRvAglM+baTQBTkiUVQsNb90rqTpwCvIK8ioj1/d3UUKMnsIP
7NI63zKBN2d1WY9a/B74DK5JgE6Wfwj3AaJSobywqAN/clyk6U4nWAh6hzIuuhau2Sx82hyGMzpg
bFZTB8FFG+qdc1MHy3szJm+KeH8V994F7uqDl5Vjsb9+iB2GuqFkFC574Jm4H5FjPH9Sxfof2Z6C
ZI8lv65UCBXSYPYuc2+YUnXJRCMQC2MhwNKD28i98fagUewJ7XxbYCyVbcgDWWguT7Nhds/8+bSP
AGXF6/5wasDVh1g5azjZzUJSAx5x6tTIGjssZLBfB3DfOZscNJzh1OyKkPcJJCeZgOG9zGpeUd2m
8X1Sjiqhb217g8ct4x7AXGVd3kMNGa4iwIiOH3SrksdaMifgYSgnI+Bj9jS+60/aZg+DGl52B3ja
d+axDLXQMopx4uoC+AndhCXy9khNWST5rG0b+zqGdFor2JVIpn+Lib4AuKT62WAUN8z3JR3lzjlR
iPSiWp3w2Cq4M7WSrlJmt8aY3lfxmeitBtFAXkOxk88AEuG2xDLgeVxuDmnXlLDzEqxOsJJ8ZlsT
qd7ULsBCrFAT/+lxpTLFFI46xcxO0xCM9fX69lSYY0gr5y9uaw8jO9dv9a5VP80N4Vp4/zDS4/3Y
swEwIPtvaQ1QRduT/MMNaWWLiZbaOISOdtwiFK/pQsHtiRUSEHwn8Wz7YMfbc5BLOYH3i+SceDhl
Lc17oVzzpTOAK89QgeZ1I+FeqDS3eRGpTrtCxE8/LH9LvUTjtU30yFVKPxKdFbw28xX8n8J9NG3U
RGZY+MHy0PGAPhGKMl68Dd8HoBjy3aBocgjFPZELJsmckHrz+oIluz1bEVI5uV35HzSt93gbulVA
/UfsDd19fgeZPK7NUex8wf2+nCmCXmUo1ufGP+OU3TN8DwS5ADumRksTgwZ/V0nzd76KEFdwNY15
Sr80JIiHmxsIGe6ewld0U4KJ+darAeOTEbIwcc9W/lFNWXmTHkHsiFPBQPErz+SvGbPxOd8d1Xn+
zhVSKQI3rUk/z9QB0aD8FtJDtB+V++TD4YbzXGenEpxE8CJaX9XfmYVzELRGGCa6b4IIxPDLFQz4
Lm/wmx+pJ9jOsiwrX1NutDbfTzAG6mXUcgo4v1wfuGNjCAjl7NNy5lVk013lsP7GfwFEy0FFkSHR
fLSyl0UcRD7zSnTdQw9lJFOG/pZKTjveBjpLeVDRrs9Z5rbNX4IZGmZBm/5Iec1cHJR9Mu/kbvw3
w2rAqYxEYzsAd+yKIImL/kklbqyNXQ3LSYF1ZhPzrKHdtiNoYdK+ndrRsYpQbPback9HSq9TTnal
bx2TzGim0gB5TUH1sfQ1AWsepGcUs7X9XCOhRGvLo2JYC7wdgaaItxUVWiQROmJAkM9MMqel5fro
+yo7/zAHM5MqoOhXV+vkRro8oZxVJyrqu+rRI9Asp1Kt2IRInLZ+2fwfYUnEBk/oSAQ4nxVEiHTk
91BSnCjAg3Yo2B62SHxni8vk3kTexKZv0LEBaQyp9b5hLeMKJQwaOSmLYEjdmHrQ/BXNb+M3r/hz
lC3s5Jy8yLc+iWcWs5ATWk5/QhekWHN85KFIUnFTgw7fZ7ztS5m5Kb6sNqdwYgy5Nlm7g2HoC4CD
kTR8BBgeGOFRr8Qd8Hxc7gBhfE44BueMOEF4kV4XoGT56g1FPuMZc5no3bEaBdfNeP6zzAECgfvW
OR1AJWPKBbCXJWkIDXPkqSIz0Ju7n5qPl2MuNr0tK1ey+3E+HKJZ0IPRjtK1SradkGwjFUKRx8NQ
tIB0HYpzapEpQtY6CjlyEmiqYeZQBr5QLLcYxvlyYWNrt9ncu6SntCP9dF82Il86BYlqT7oGfI/Q
rY2RrTAi1OnamfR7XF2WimIA0hLeA5YVxmIMQeQyigiYPDmPkzf0rmDfNuB4pT9f3AR2WwzQn1J6
998N5OuHgrCuPXC8hlMFUtU2lAmAH6FP0iQdh2xoMIuP5gBkvN0AOO4P5Z+h2x7U2LcvtrsDau80
5+MScova+xl/DUtkguhxQCCXuzjyRwCQEYHQ6E+LJwe+dJeIL09QB59sJiUc1Fu0Iv7pTckpaty/
CpAdsGlrqNVdbEpnQJe29O8cLAWEgWEsEHAQsBFW0Br0qicE2lgNqTkSrIw6sC6SeSHY6WY62uS8
FlG7aRDAqPNDEJhAGdiMD/Oiji9vtAsQrL3AsLMv/+ffJ+kuT4+GwsJElljdo6dCStxBr4XznY0u
O5n6JOTqNBis1v6bO6fBUK9A7YwdklqdXQ2aOdQnl5gBL3Vx5hfcityRCZ/jKJBueRIzJUgNg6kJ
DeS3JxvcPDhV537klZCz1e2+S3fojR2poR9+/xXY4GAjp1Clor06EAlfqgy3id/+Z74sMOZ7BK1K
pq3Nbr6AqBaT6mW0+KaVzU6NeE12fApe5os/bmcTN5JAjm+VMtA6OyFV4KroymBASuL3Ifv5Tq92
omGROeKvCytxiB0DCOxmozkNNx1xhqBgCnspyWsFrLXtyM1FUgmgb2AT6H4OiMm2BdNp+LejhYB3
3GIg6zkpoDQZWYP1uYEZQLiE/v+XCDnBt4EoZSUhbPoDpBKJ1O8uV07CPSX4/f5Gzh4cg9PGuYrs
5gbyiOr55c5rcknlyUv6D1wXnfLBRtgYJm3337iXF34Zb4zHo0X5AZwkg7ieV7u+n8+Uh69I+enm
FoIZxuA+9dAKq+R31n28V69vrEbTeuBD5DrUHJLnuNU/rsmF7x9W62tPVUdP1XRbiO86VWQqF2z8
lO5qIEtLctmkAwHj6IMylIGah7N2ecXU1OwAR5izJH6Yb+TjyfojGwn29wFxMVIZMcwv96lSLGs3
XtSFesoq6rlx20/0Af70AL7PhWQReLkY60LYXhuHqVv+f1r5VROXhpa2PW5qhaTxSkOo9GpRqb5F
3YYGLEVpZR6wFUIuG6Yxs+FTMIVz19staHNtvr2ZMhn++rtpH6jKTakeUS717hVRRwWH/DmzMZ+w
7dZ5AYX2surtiXhjCO6qek5tCziuBXD4MMFN/BMpVRQ3vFjtkBl29WaFmpA/qLqOYjjsFiPWVscG
E3ctGwb8mBhHjng8Ct3odcnFMSf7zvL29Hd22RUX8O58dKt+l2w6c2VKYHYAfPmA4TcKuPb2uy+u
Ew4Ufob+mgd2R0fTeyUtuzyyhhOkzYFFRxk4q5WiPnu6TzUMV+FJ1bEpAXSTHToOfcDajWV++++f
R8oLExjreMwcOis3vQ03aHXPKOLu3dvZy7YmKefhLJdODp8snM6Ik6hw356T6Sb75XPPcYLIyWJd
+ctydRu65laeF0JJbRMYhm9fXXJC3Ph2R9T2apfa7M2V+ol02RRlY3gQ3mAgaDy44c6qq1mS//HA
pBG7DBdtDoxgOGeEceBQ/UF2XnORJTdEo7YMcSPezziE9t4cEzi0gnUPqOG4IVa/MoXhpYTZKaa4
4nHnBU4I7zJsP/XMxjBs6RSomz4NjwczSS/G23OGuO1edrRsUPHnKtBxMZUT6pj5iZwGZCEv4Kqj
KWxIfyMun+3WPDMK/61xn7fya7Z2ALn9wp5q68bD+S20nhhMxuE8MsFOcM9FaoHDBpKThtoc4cvq
WNRYo8978HwOqcG8ayVqOI950d5As0Xof9fBvdh9t6NVbXAmNtoytV7jzBBL9MV3kPKmxL1GWQBz
By2RmiyS5jAjpOsDxj/dajFczfVu19WKvPcsjskgWTLgJe81NzH/76yjufSe4LxObnrOGuAQbZNZ
jM/yFWkeKQ8/7qWLlT2n+QVpLEGYi32lcllLz0f9vugpt2NgC1mdfek3XgLwpJkchqcu3800MRH9
9vWL8YNlwrhn+EN/7+ueZmN1aqqMLK0rDSk3mer3OEqTlRHL17Q+ArhYASgpnLj/F7w3D6xoJ/vl
27ShoseWLCEJ3k3iYv/S8ppmTztFzuFYzv2MD9Sep7fauCSmYcxqlumRYZDIHI4hjdeLrbQDAh7v
sxYqyCTDfM39IeQyrXan9DhK4TB8xLghNSAt2c0LZh9t86Mhgv95L2w7l2/YYvNx5lhwW1XtFH72
mPLr23XoIMeavTNkNxMGKdtgIe2Gs32zha7dvfQb06QCvqBf2YuZOmbAliUjSJ0eO2Y2jYwYwviv
YciuEkoCzEpOYANHtTC8hi2Rgfst5zXycyUat+zx5fsTcIm0oksopLeGzKtx/zsNiSBMoq0ezV4V
f5MW5PCtk9rF7iIGzjPQYqMkPmmDE5WtLI9VlQIokukWTZKpT4umuUwmsv/vmZzkgfqmkTKZhn5i
EGrJPDnIj2jJ3kEvB9gY1vveC0nwyOkcQlThjiiYiWP+Ao0i6qm3A1pPcpP6cAb4Dx1Thf8MWSDL
vXXWfGfPS/oDw6QV/zq46P8rq1QlRJnD2d1AKMtMXfat4O0Hd3nRxd+7/0+B2Ha4/425ZU9vX2CX
znUCJQdsZaVCpFX72hr3uWuAgA8AUhlpPsACCWEXgrODQ0mDLPwfM+yZAHDG5OtzzC0FALPKRv4P
ZwzGgBovu6cn5xIkzOkPM15/3JQ5a9fw1nsu0E3mI6C7qa2zza3/hprTR9ZMjcjLzXwl0iA8iJra
8861WBAByQ+TpWL5D+yAF8TEe580CDe9afIWrGL9t2K4gJI07RuaxopwU2Ish7rIfjOZoOPjv6xK
pm0Sdb7zdHLcxG2tWOEwQvbGOVTtCpn/x+X2F75N5DWvOGqmlhcVWQS1WRqKBCcsZbyDxwMQ02IB
Re2Lz1tOnxXEb52JW8UipxDHvzHZLXDAJwQ+/pMVUGw0YOJyIOYO1Tue3HtY8YtvTYqIUcgMe//X
rAv4kOve8MnxvVABqm9XZROV1SMFzyEG+Aw33UGGH8o3DTxi11g2VvQrqr0h7ALbqItWqnDc8VRu
8yyq9xip9pakcN1JJaqSQS1OeLt0fpEcQGf5wvqWoM/cyfu6uQPK/iSaticX3yDLUYGUb/8Fx6X3
8sJocg2cWjVjzPI6bg2fRscNH07bfTVmvjP8MffVcriVpOid3MwSJT6SfeWXd6cqNwwYa5GMAkm7
0QsULd0IjTbS07BxzVp7G+R9z3tT/isF77pQGWWIM21NM7ho2kqOKCIcOE8+yvNOGdpqwyyATfGm
IJMxv4ER2Ty0aBvSVDk08EGKT22IW/qVzvwiImGsv0oBYZq+Oq2hAGqkQ8nb1Bqsibu7MpAN/Rc6
QGdmgnVUoouyU+6FNcElQjKS7FNcg7baYsF6UoqfWI9WgvWFaOPDh+nSwtPXhfJsjpToI5QJAZsL
a89Bpv5883AaiYjpEFtxrJ1rCLXKlpWKFYAnsgED8FYqjCuHqV9VfXpSYuRp8MjblIWwZnvntBSX
FmJKd6qaESpwUjvd1FfEWcZMLUBVXdxFXvqnKXjnuQL39S5dS5xyrV8eSUWPxK7aNV2Nq27aTN5/
QcUNu0w+5KYhuq5Rn/ULuPEDD+1dfAShIFsvby9304QQ06eWdqCFqq40EJ9pYaGrUNq8bORkCmox
tkhL986+t2PbvVtl140JK4w+oPhd/J33Twl8vREfnDCoZBXHtslO8Vtf9sS+p6cblKVsxzzinFsc
B/X+4BRswfu9DY7hrlk5k1pKWqLnzRw7Q8FJU7doemCgXoPEJ8fiMsDzswCi9U5XREnRb3z54fdm
vAiRR51ELkRyKbC+kRhVXlbH70JdhcoRtyt4RLlYvd5mEZS4NTFgHKTbMq7SflAxqneQPpFCZtmt
qSfmvO9DdY5UdziHKouFUybRtJRjgaQ0dJD3m2mXBSYms00WI6fPioV5Vvyl4lBCC794YBMim9zq
7dfCGHo2lNx3EmaSLi95o9GaNUY2VFZfkEVgiolHT4jTqYam6OVGB4AuXoPbi3ezGdMDfR+zuJkE
V7nYSR8GPVumuVJs6b0rNHyzUOJ6suhQ7AGb2dRpjm4O4SmDhJasYPq0W0uflqxCPtbqPDBNOp6Y
DE7OMrZICxBVB7TL0XhGQ0fHuVMkMVXBLYTQtDO1xIPKDlg+g1+b7VPrUY8iIqTLTcLI9ZOp7Xho
w/jEfEonTE4MpVeGKd2ixjKKUbzJrUp7m5KpW7sKRZCLocB5P1v2JFVMX0w+wMucPouThvGqJp+Y
zQ5gpz3auyecCKs1H/+AIMgmkp67OEIFm6Yj0sDpsfnPuQs3EyP4KjhIA5HSyHcjRi/vfiVx9lw7
PaLzhNFCnbsAwsJ50fd3ucjllr9mwdjq7MsEGieO4ID+v7IqsfSc1IPM1r8iWhhOwdCKpB7xwSfz
/25uXIbhIR3H9L5YaZ4x0DWMrNYvccc5Tbnb7RR6c6XTCbpS6Lmcm6i51Sm6TOCaLoljj9t4dOmr
rQMGZeoF+g2Ie9mjv19CvzuzO4UQp95pI1lTVgesGL7Yfy3jKn32fUg8IwlwsAjGQX/uZsgaq9Hn
55Ha8P6LX9M11qW3c0chdpz6X+lZmtvfQ4Br7SI+daLL2OXpXH2hR4c+cwHLrBRj49jxwgjHkCZ+
QlTJkBOMO0j9h+XssmjzFwQF9WZBMijVghyOwWUODq3CcO5asBkrVsn0AiXm/izDG/S1Zoh/Reyj
b/jSiO7sGv5e+bqAAJimYwSgFmX59Z9K6v9veFlwLj56bF0sj5mPJF9gIkk0/I02/AtAs3Jg4Oyv
tD82sHZGWYeSJet83s/goG3wcRloMYw0JvuRE91Qv1Jf1ZT7zfRkIaecCLb3BxP18hS2BtBfcegB
sLtMUw7C0jLTR29n7gX8jm1NwU/VmgoI+HwE+x3mMqsLlQB/yK9nUepwRMqjDHmQos9xsRcg6fam
Rx/867/afxtdkJaoPUraE7jYjLcw3TGqwX1jBnvYYue1QCBIw+6nnR4iyEvKe1NSlco/hiKU7CYv
hUQKEYL1M2ODh7dEIMsU4oCPBOiMSDt6xq9D/W5FCwTfp6EfJqh8PSFNvdY2QG7ykgN8UKTJCXNc
hdYhsHnQVHEJ+4uesd6CjGVE/R+hxLwnVeJY6cwsY8stv6aQK4SFt0LBowabGQfjJ+wSTWYyO83s
IAqkdiX64g0lesk+aCW5iX7lbWoz4Oz0uf8TWk8aNKx2Ddfb+YgQ3q0ngp1vbPdNILS1RvaGWdIY
MN60+7uBiT5SJu9s/R2eh6KNsBPM3Qvqt18JVQzXV1RlasUHQc7T5uJ51XSABSk51dFs5Qf6Rfck
1sPeL5ijFTybIdZd/WYecS07YFyQRO/2yvgXE0HHmHzMKkQnOcdJtQYddklvIHxrtssLx+C2mdyk
wnN7/pXyA8toZwwiZOpBYuxj40YZhbnPOe4RNMRMKCdVYdVCfpwGUQxtxmHbxv78LuL5EClFfOqS
/N6XRFvdO+p9MelGfbzlI0CAxQm8wGkztA0QlD1LmRT1iQ+JQm7aEicaSA4oB1WuINOJw4JY/vaK
AC6rNBZmHm5xtjTmXzqWi9bD64Hqpra7HaiJoeZb7tp6Ytz+3SsUnFdV6BY31/02QMWqhJWbBM1L
FGfqirXgkR8ljDa8Hpqb8lJLL678Vrd8MwJEjsvEJckSYGXc6Fly5Qyk+/Xqui05+SsKyVTPPpY/
9YGPsJ6AOVslxy1kKo1i5wQxD/3HZDfx7+//6EhNnJ8yt3DEk5zmP6PZ3UgizucjRJkiLU74BtHL
pr3CwzhZakVvGEObpOycknlwSjyC2wTPqSIy0iGgwpGvYDuevwNeDBVb8V38YRClMFyxc2PJjLs6
XecZxG0VowqoYoogID2Hve2SOXUrVHXMA1ylq6N/nQrTlHFglTx2Uu6cmpts4KuvcCWNhX7ysVPq
pBZhWt17jujfit8ZiUvR2m9oZxSLCxsdY+sf2cIIrxE2v2hvqv/GcbyojF2MSWeCFlX8YbF7f216
yvJFksQZgvU3meLnJE3e5es4aRvhINceCrDm1BTDhwxLkgXScMJbKcOxTBrzVunSJVuRZK2OmdnK
YlG+UoTjl0TXYBAMP2xEAYDfJ9n53KyLIPgdsxPT9y32MHvvKpzv3ToHAS5kJp2OeZIg9FHHMgtg
k1qC8iuKEjIFR10J1RJufS9BmfFlCxgzRqVgMyOn2/KsYGowKMfKIbB3DVbfVg9+ECL1NqDLs/jJ
QkQaFnMJFb1StlxUYY6A1W+xEg8SKJuCbFPgXp1/b0jMhPBqbPRe7+sbKdhBKmTS4zEi7Z2ypu3K
1WyuOjEJ+WlZEPXqx+zjFJFcS4XEm7dMsnKxYwSyPnNG0AQRW7bO8Eb9prm1a5ktFxTXyi8dfyG+
jw72zxBseWXSFIRJo66uJvblYoEKIY9rWUtRHlhhY4++78HMAE7JVbNlDy2Rgu7q/Wu8aTr/Hcav
kGW2/ooIGnwJWOeWKgl3s9ug3GxjqxISfOM9TpIptmi+ahNxk9cN8pqKW4AzG7xYsyn/nRSjxjJF
hVTTZwJ4dnH7871RROPmwTtXI5tyYX4s550Vsjne7brzs97nJ3oI2fe2ggFpSMm+Wv893MbKcbVM
yIF0lQfddbcPqFQ3g/DFcJJmRrLLSjOZ4z7TZeGK2NnaBfN2mxQLiphOY8HnaBZq/2WlV0ekSdZf
qIZpCnNpPc4mqOVsGC816duYauWdTx3BEtf+zrYrH0ENHuDsN/T1M3UCJxO6c03Rled6Fss813yt
VKkPPQ5rMBwNi6QKNfiNGl8jm72gRTn4mykncwbq2SG9jTNWGIryzoNjoqYBXMeL0EUyPZnW2PAy
RshAgMSHMY3eZE0aCbUJCO6D+I7Cn5IscW9KkrebNRcDJIrL36KVKFPqgwQS6CpaZS9y49anlLj7
RXgNhWxPg09fIS3KCtRg1WgGwsIvJEkQTCXk8Zw+x3biyC4TLv+PtEPIzgO1fvqFh2vrI/2/GwZ6
Usg6IkrlKfADDORHrv1X+qrxuM9+MVKmteNK5f9bK4Cr5n7vpHs4eGfzjt71uW24WD2yXwp/deH2
O1BbksmnZg0xgokYUw+aifYRy+Mdcp8ig3pJaOUL1yuzhbVhI7noU4rqUNImAvx697ru7Ba3jorI
yhmjIIhTWXwo7jjc0Bg8xxPDOzbKkfbuaMF7I/a86Ot6W302nFZOm02YREXr29p6SNenyU5oIUn6
WgfC1hvBT7Le7lmwOBlkrnm326b50utaAgDd61924N0VhgxkRFvHOQRn+QgvzxRw1BeVSMrO9h7m
IXwEIjCMVzZ/g09zyGtX+DV9K4FidMxLEt4lhM8HIObTXVzPvBWfI7/TPkCdKTgxZxW/HZq3zJcZ
Wk4VO/eM0Lctg12L7clVdXCV47F/YHmaClZ/XqFMbgv4pBr9k0gD+taqDSKl43Dnh4LlblLr/sOn
Q2soDQAPTW0L43S1kDbCVjSQaf66VIfPbhdjlTe2od0ufJ+FKjHBfd6Z2NH/SMTmm/o0rauU+SZE
HkdT92GTAC4jq96nppf0NSeQ0sUqoj+cjFTVlv4aoQ2Ezrs3SuquyXBGRZwcsyzrMf/Ec1WcdoJa
yG4TRi1ly7+guqsbEu3hlrByJQx4dzCcJYbAaEDIVO6eW8fdQ7a3t1P4T8hshKCV4vdJPaks86ul
bIR8DB+5adOn8ppWG1YMj5KZQloBIFCL5Vk/5TNQrznntq0GVz/zrAVH2QK4nUlIRE8SW+M46JGu
zBzquvQzF4KTSL3KwCCiWF7pI8sHV5/svJHjhHxxFcoLYI4eS0SNNHX5jjDpWJ9AJaIUZOBw3aVn
7Z0zzpn2qPItCCGrH4bZ08kWwG4FNc1WUTK7d89sBvmsEDeA1mHXu+XFKFQfTSP0KW7SbKWiF1Od
oTlRq9XGh9b65pYbmquvMBLjCaQqLmVd1Xl991S1fqsN/X53wsNTw71NEGY8Zn519BzcCbQYOCJs
d90hd5Gu2gTXLTHX8ZkyRKCSfRp4f68NpaOThvOwDMP88uI9h9X2veUNbMEOBwk5RTU9wfojPYif
FN47lCO4yO+45cS0SXdvY0Sl4PL5ji7ZVBsiZvCO7vlFP/0YiLCiLlccZ0DwbwTQrAsOSd+C0J6S
ETRFC3WBTIWsalzj9U5mkh56zwZvEsHLv9TvX/rUavgqNkT9ilnfVNs2tWuudmqjukB6jR6q6BTs
JLoP+cVnXwjLucqTDNCQbTAxnwExPetD/blZL5578wIXu6kb64NurbdnMv4kGW5D3yWJQ2j9pydg
jP3gRXhUS2vOj1sVsXU/TlfYCIHlkqtQqpG4azrUdlEBQZsH/CWvPYvRh2k6+SnFP3GqLE4Ek41Y
IgF5T6ABGn6OOVFuPaO07h3+VLLn8y9nRFlvDNbREdgsS0se0BudTUzVgKyrufSEmun8Akcl8SA2
31r9QhbhzxnhGYRXcuaVi0V3oQPxs+sAVsV/tVI7yjgoxxJNfquJZIzQYpqkxsMIxSOqfPus5rus
vwKVIwx5YcyQEe+vBq1hwwNhKICQeuXMXgTeakE2gPi/lLMowvzxEVUTPJWADlWGio87lh+q62ax
+RrB4EVTRa5wIeaX7443gMYlzldjeuA3OG+cZP0zw+Ag32DHhCDqwFrq/ifR4A7zLDasXPnw7zjh
8OogD98i/rAjYDbTOZ40rdNBiRTCAZpcfUnfXxvtVTQKlyn+NAGJD9eR9kxPHPYGSN5FcjqE0wVY
1VF7vW4VZVjIlrB/fdqagxiUXPERzIsmcdlB+zL3uzALYUmHRPz7dCLhr/xWVkGT9pZ3DiVYki9L
LevDUGvLvasMyf37iQt658Bkr5XTmIYVcLeGHO163/QKEjKYE1fi4VbK+lrWhndgy2gl1Ra/6ZMf
CgINNo3J+j5h+DYzhCPFXJONUSOZtzp8sfXMNkV1kEQp5IqFMIn0eUxJsFYwDsGfZI1da0/jl+al
Ea0jn7Nr1VuIte/h/n1nekjFLafLBg+ULXptXrZZVXhVsa68FwZ97F61nDgxtMnlbuGET5J6a+Mw
z29tyKZMoc4WFktU6gK9F3k8kBkI2aNgNAmgyzBz0zOGsgQ37cdNUH6y079pPcqzjM+kQ9nBg0lS
t2qEWB0p9rrvCbzc0m8LjigVZKAEYex6KSd//ykTGBQK4XfG4Esj7ssnGEYxyWyIWvKcG+G4gmEJ
Mq4uDKUUCWDGdI6xDgLdw6Ay4a72a4pKbSy7/de7l2z5ghIMfsgX6v0njECLZI8GfS/6Fa9o1o1q
mGeU90aBcdT9BsBN6GqlsCCEXVAWeAP7xiJT36YWwFFS2N5WQZG3xDrT+tlEq2JiRu4JINy66Dsh
kFHgLHyig4tFSOFLzdqqZPAj2RkR6NpacVb+wc7qyqW3ApU/b3Onl+XPnYIeAAgHJP2B/MMNv0ya
PFWtVdk4MJDmPFoyA1huyDL0N+6/uPr7hPo7rDoNX9GZhmT5lRhZch4JRJKxXES7uYaP4poh6iHT
TppaGgd4oxddj7M54JnSyNMQnSR5Y3yykr+DXS6R20wcIIgS7cEFbn/JN3j7DT3OqmX/htEEr5UO
1tBRrJ46mJvu+wlA8xv4Wr6mCu/zFSnul8EKEyrFmUx5getpQq7p7VuLzJrYs4f+0aNCm+/HKxr5
nIvfpmZcCpbqVzdVkR6hKB0sQCzzayE8Rao7i/2AomTIjZlrr8tc50IrurQg0wB7Fv71oSjJJadP
21sEJJrR8uFqT+U2lmT7cY4pSYlQV4kbd51htIOeGQWb5+3rQ9xdu+AtA4VDDSN4q2XjT6t/5K57
+TZ6ZfNe8XcMIFyKdzKAWVzocmZK8OUfTP7cRkBsZGPG5K9Cy07wITghhFwkUUZY20+b9OpFhc4F
nTWqw4k0s10R7CFQusjcj7h3t+ZyN4h8nQ4wV0U+AqjXvJ1Dc0+MaASXfegUMIv4JXAGw0JcWU15
bFhyzC0i4P8l4BJiKg73itE8tFt0GfoHJAp967eKRa6bXzOTf8WaILfbwHn2fAFBUS8Azk3ZhX5Z
DKECxMmK0VSAYJ8ep5dkJ/12ArF/l4jABkzdKPkg1fIdta0Px61yKi2uLiYnZPWaEhmkl5fxHSf9
FWXSv51HMwui5gAYmEpZFoZrqszL2vBdgSfeOikelCVrwSvvZ21b68/yzzuWEceL5bhVuo/2aQGr
x+jKBNAINowjuvbBTMNnT4/7z0/XssfgQz04ttosk1i1kb2JoOg8ctjeRdsPJbEvrBazDLpWrBaD
6Qr0FhF4XhBeOJAO+PiJI1qUEp+WovVZaVSYd4hCRZ3AT9OjTuPf7fUS38lWHpCHaPJK+DNV8m2H
7IJ+rW/4+0zegTFhUjECtmmkZ7zZGegIG46O9aotlLJeAYEhGvKQUn2aRguFPZux/9pfb6Q6R45j
XS1GMj8dPoOlboX6JXzD7dX/FKIDUyiu3CsFAuGvtSM5JPy9QBg3cFn11lfTGooSW+UTUwg1CnLq
ZpCoSG7RFcbluSJ4TuhFrfYWozhfpj5MzWYSbf63HGV/FZP8EKUXWxStPHSoOkZ2YXua6ApL5IKw
YAt58llGjNOSEImGTaqGp95ZRU3uNZ2ZP1untVlOmGEsH2fIG0KgDySSQ4onEDUHYpjQw0lMvwtG
V2CgBpm3nIwNv4pwxL8cgYt3dEpVIF5X0WcmV7tws1a5rbLhgs2Lfw9Vk6Q2rfdQJgf79fcFqnrf
lI2kyCHV5L6teNzFWFzC410i4XJboLikuigGd6BAXZ0fqt++QVDf3AMdqzdjY5DTzHNnVjk5ktcD
8ddUF/gGFwmU4qIib+PtLp2c61/GB+1znFn3z3ugFqzINmS2qt9G+HT+mZvvxpG+q/TAoqaeE55D
11FkkrektP1daCDMjBIT/tCBRGdLC4R+cpyNf133hXjkGro8QIH953tdAkPC/I7ARiSVXMMF0HLd
ANiBGiQ9LFe24Ek+CUFysU8EUqB7vHJRNdmzJEO9Gs/rUd0Mx7GtauAzLqcBPlKLJ+wyz3L7V80d
o3jNzQy7jpHvNl1hj+ht2h+lLBdBa9sJOJ75KZQ81TgvMqO1bSBk03kC6x8f1Xsif2vmm6gQwvC5
LiFeY1R6VBiaM00dxYWNJTB/X7KpePFIvgsuIpERiBC34qtwvGqcc7j1LK0U6zVnkA46X4yQe1CC
vhi4ycCBVrULEjROT8zAJdsrgkeDGcA4GpvnaywGh5zCnf5tHG3LAD8sI9LuXYZDQD27p0B57HUa
pVwr2aVvW3kKJi5Vp2+LZOZoyAL9o9qtNiTGvnan30d3DQhcstl0E82lbggCbHqT9BTUhsu7V5DO
sepsAwdsG4sQjhzZ9GHQEYIeRQ11AicO8LvQm5TG4yu3P9C8bbhw0v3RfX8nTZLnD3eeOuCH9aEq
SNIpOSopiGYTmywz/jJKGHp6vPwVxSsKCkTExSY3IDI3w7bX5DAdowU//sf9TkNmzCf/16wt1x6h
YDgHEljNp44j+t5AtQ/NOlo7bW5AxbY+n9P0fgBP55NC7JGgOauOs4Fpn6L+/+YK6Opyl+kEda+o
gpExyKgstrD400Ayj4+g+uBfqfWNv6NriETnDnNtMfcmDjPI/3aynLT/sWFx+W0Lhdi1LZizADTn
SberKqVtvmyprI5bYT6B9dmhI4G6PrfJk1mZ2t4I/DsfgV+rwyTnLE53KhI9TtDsnkIN8IYok0Qe
ATL9jtGaYB/ldzgkLMA+62XHW3nDqt/q/DdGbvegEZV27Udaj3HAUyU6DHEU94ay1N5juAUrbD8C
AOj9+0K4ubZs4p/l3WeYQlThHbKqxRl/k+iNNt660So6v7pA9t+yV1I6U31EPZfAX78iADZCQEsX
TtmF0hxEdfrufMN0dfyt80IS4k7CU49CLt9CgyDmmFm+KV1fnKUCy4FNt4uRba5R9SY/QgKW3Kru
1Wxd+YjFAWvyii7S/qiLmLULO1tkG9RJfkzUUmuELXoyVzOatc57KFh3GRx5/XB5jShJqTmWD7k1
7G244dHSBZKKp80HDzMihYOlBucO8bZT3M93Cgfn8IJremnv5e50qAQyt6Hgp2/D7sTIlmYfDzHB
tZX2KlSMDqidIjC5Qo7kJ0EtjpsRcL13LyNHEtOA5J8aejvgN87Ke36iZa+vq8Xj+itQVWQ68ZKg
8irpCQtRbYHHQGX/lfb+qVlgxVWKT7P4p/tvatCetaigcwLu7xnpYALfcBo0QSHv0REYvFn+w52W
wFvnxuDN3ybCei68M7tWUbCa07q/luR3j1QM9KH2scuqMHF+TRHBQtKoH0Qmlb+tEcPjsfC7CqQc
YPW0H3Oj0WBZqTUvTTIK9KF0NcumlfZ+KTaqbZjV+cAIQKixRLxI+Dq1Id0NOXUAOl5CiHxi7UV3
lpiCuuDx7Z4P8DCV+BH4EzMlt9N5JohoAn7lJJM4ZUb3qptp02hU1x8yJwemFzi1qqzXRnH5MmxQ
zzNRcP8UulC0vsI1csZLT1Q03KUTg4dQCKvRorF1uEd9N6pae7F+MhYZOekLjRb9ulV65UmYFxOq
mNRqKEG08btR21B8aoKZLZxzeuqJqgNUr4SUFVXMHT1/H0FtQWuhM6QeN838Fp3ve/iX8ep2FFGw
D6yhHdWPxqRekFKP2R8T6nynB91R6PnSG/kgCf5Q33976gZxTNviJPDWLhZ4J2EdaM6ktgTYIuSV
plrmq1RE9jg0Dj+Ysw5nk6l4Yldqaa8569Xbu3Amw03IaDgK4/47TpDcfKwML5uSjWJey+rPWwRu
HpVgAL1xQdD5LNYc8AG8beZb355eWt4EDLzPpd+co0XZW5CzVY2fhk92JrQUF8BEJIcLFwXoBtaY
ksjyKaw9CwRGrhnVRPxNXR2g7cyPYlWBNUTpd6d2+Ufydtlp7dRxglJ+2v9kgIXTZcNYvo3o3cOp
pQ7qxYPTt2db8PUP20O4CscgMFzs3tY+JBl6RQYj8Tjq+HtIJ678R52iyppMu8t5aIR3jYmC4JMp
2WW4PQOKjBxairegPawc//0JtpLAVp0aLOVQSyNmQq2EO7oXmV7YyUbvdM+LQ4RQg8GF373JNgQr
qkdRKepJ49RL92Q7X6KhCsqZu/dqzvxvKT7FOpQM2Yr4y95LmRmuHIJGDG43PdcOF6mi0HvdH8Eh
Ha2Zq4/bxVjRd8+DmZtY43D28hAtMT07uLcc2OIy7BMkmnFx6vXA/oBdSFMA4PsOo98CB6W0P+hm
mduVMc8I8C31TvB0rTCrFZ/I4dZbi8Uo4oU38V4OREw0ADK/Ij9aB/1dUNnidqRBv1faC/Y8ubtt
c8B1hRie0c8HZFdZjfWkhRo0O5RP7c6aWtjgRWHxuKuGX4jChkd/U+DDImQPgoUoJx5dulJAZWwR
plXn22E719TThcxNE903FKFRdxcTwtnYJCNFxouSQjggx488pFewgxBZnw1BUXYzv1PM55pRh+RC
gKzJ8DmvMPBolCEcrhV2uund7Xt9Q1tUP4VG3+3KmRfpgUU0Mp/MfiJ+A7brFqLGHVu0TZ2441Cw
FnYCc6glKAl3D3OOCN2dPpNp8nisbbdfhrheaC7CaWBkBuJAuJC3hjbtltrRAp23z6d9IFrjY0ga
yJ6JKHnN3kxjpiknwUZ1+AeAMSFHnz7fW6dedM85pWujB/LSEeCi2vDLpWgnwLvW8PDNgZpOpebb
Vlk5cMs4RBQ3qitZelfoj4+UdsDq1hamHHUTNUdZS9ipZZln8b2hpAYcvdHDBEyGVfxkysbN33xf
dqEAwm/OY01/fFeXX+UO7rrH0hQMKrOxlvTMHs0NGjs3g30w/KqvTP69Oslq7/FqfcgaqKRcnA1F
kWt9dp1EIP0ppuoEaGLrh+4i07ISfQ8IpK7CMrpxdny/xY058kKQRAVyb58zCv88vozB9HWLx0mW
VK/dKfU4oTGaNLxCOZds4MuwVQ+ZkQqlRFKlLHSl4VJfkIcw+SAkcSrqKkjMI4Tdfp45BK0w12g7
hGEpgtGekyL3mA+A5StjdbVCxVZ0xkGJvyWFAeLuBIDwT9QIdBqDqES92Vd8KY788KdIRZnQ8gL3
/SSW3CKJi5evjEVWVU6WM+MhGsynhbw1BqpOdXM24z6t7aDVVRr8oOJr4wrPf9eA4fZo2gvESMH8
wi8Jv6P1HIL8bybKgeTRqXWAGRYEr9akkrwJ1ad3ik8bgZE3S3u9/ywUq6VODTRBlAvxg9spHu3K
XN2FWjZk5mK7lXbbKF/12+flF1SkwFx8ZIo+FHSpCDmBZvF5alfvUbQ4VQ5bmyBMdKQ3zCr5vdo/
W1hsaK+oerZXUAq3hG6DxRftpUh1Zh71EJiOXV9b8odeIe+ymdpKGjdR2gGgaOpiuiZ3NutLiwar
l022iEwqnRXnAubHyPuQhIY5xhjDj0DdHsiXKClJj30PNG30mgOAAvpggB+ItejqScF9hPV4d+KR
YOmBcXYefK1LkPP0MtL58OdV5+kAnRLDzXSh1HD8LUmENS0NakHvg2n7+faN5nxZ3kxOT3xQrcHq
45bKD8UWyYaKMTX9BUy0qcsCGDcROrLsDMJbNikG/LxCAQI7uLKCSEhS/tohj1aMzEmxLjY6hJu/
XsQxnOcnZdFJTigWwtY6Ho2M0zUoIC0tULHu/yAX/GkNdWsBVDb/J3R8ElwPW2bBJmfnRbb+uJ3U
TD965rEn0fTmwVDAyQTlxfXIDSchspX2OCTUn2e1g7OhtkeAbDsmkWWSdU0Ei3WAk6Up7Dig8ws9
BuTuWnjredV1AT3KA0+4OEKVt9tUK+7gMMQzyHFm9HebW1B3KA/XrJU+8bYYHJP85zXVNLxl6UBY
j907MSFz+5ucU4QJTRwghm0xkoqF+c1iNjrmjJAgLtAHgUVBnwgBB6i3bfwd41bnziaX0a49urA8
gqODtIpsdr3Dg2IW+3xGAT3r9E8gvTZMfnaoiWLrAIBYVFTV7z29zBtIJNjK8ZOVgq2C64WncDt0
A9CNkJuigk8D/S2rxibOJjCtQ8EsVrMB2imrT9D/FKt0LxMC3WYh5lTJ00255Px/ifA+2/F5Fxoh
XXykup32yapJf4y/bnw5msy0PmPWGEQB1mLaloxblJSeR7z9SsM+Lnxwvl95IAoDJplV0Nu7ecEJ
SWgEVnuheOsGoaAFoqaaKHcIxCeCiGh1ZlGhVQcWlPdD8b/Zq+/9bQglcGJOHasZfLKszf3KMmZA
r8dCd4Cfw1IuQTYMWvHED39e5jZ16r71UDsZ4UvhVBm4UE9+CT6S8lc6aDlDpx+b/C0DhNNqICXV
/6eVEwgGo9vlhekjW3X9oWp2v8IC8SVERET5Qktp0iv+JdDNV+OAFcZ+vdospvrNVlo+ifQxBwNc
4qY96DR8BPsI6XVG1+2uqNAtzmEAT1xM/kzqguQ3l3O+dsqCJzjy0tOwXQbuUbolcYb8U/vIQivD
1Ag3DQKOcBIagdelW9t4OTb0ddKK1F1O/8N4Ppt2tcSCOusyIUPxHp+eyT6VDesMNveWqCd48svX
9cLEsq5GdpkNvEa6Nr4stbYpqfs/iy+dWgQAe60nqdQ/l3iRKBP1qocGOFuWNxDz19XIkLLBTIWV
/RRv9hEfMLRVC5O2kM32d5gyD07mnHXwCJ/PYH2JFOM3FvSVd1gTDmfE3jYY8VExyG6gi3VSkOez
I7iBXDsCrHISGF8gswReJ+fkPk+8o/1acEUd4KxakuO4X9ZCF8d35OsEtAodDUKwORJCkcF8r1Kr
xUDpnDEi5v8MtrhpGL1RAQ4qRNkrum7nYjVLK1DXusruUZxcsmKkFNYYKYSUfkq7SD94YBCxIMhF
R9ags4t74P8pVV9CRy8wkujQBPeNqf01Ypq7ZeDoINLlQYumz+MhJXpmep6inZyGUSn7eXjihX3+
Z6LMusmr+PLYS5CIQM8xUpJM1j9RWx9HjrapWzeOKmTzLv8yWILhwgPZnycAutfo35IiJkcuT0w2
3fs6AVXDizfl/1BL95HOShhCJowgnf3e48oAOqyXrh5IUbEpM+Yl+b1d4UjMUR5CU4VXdQi18ziz
g7BAyW7tH5YTFHWErEQkO+H3wpEWe6wbI4qo9fCUYZFSoYGf03Au8xbR8Pi0r8dYTq3um9Q84q6j
g787XOvH1y3UNpDm9gesmvIQg9qR7+FicLQEM5qp0PXg/xVtNqCvHveFpScCnsngUA4KSQsEPLr7
vvVU6Zsxq++SrG0ONuCCAnUzPmh3l7m6MtXMHM/ApyEFZ5tXHYIym2rxTSNjfQnu+IpTlrb+i1Ee
jam+OYsoYeAX6B5lJmKpRJ8vcCTAyoPyfnlzbBMsTFcQNyNQ5Ob4z3fsJAzNdfxpH+QT+D2M+vU4
Rbe0asO9ZIMMUaMak9/Gam62oxSTwo0DdzkYq+qVu280lhnCLiiklsDojQRRaIuZYYCITN2WPB5H
APfyK/RxrNJzmZ73B0EjFz+VnNb0v9RYCilAWJmQ32X1WpDZ8VwhExmR31dXOZHjdiXEYnV+tU3r
cH6uhoNYo7iQfkD2ep+2vKflgXLviCA3TNEO1+84TbhyhF9B4NV7RggLBnT6J1JK91pYnOcaZ4p6
eE0QvRWQJaE0NzapUcxDrH7QGK8BuEafoI5kvhIFi0mKUev3NmHeq4fgb3o0Pe0+yKLZT/iPxP2v
4Peu+3y2JO7V9eLJoRu7IZfLacCnKgsbz3dujqItbNVvKqyWX24oefWv3eVUL3uLCmX14VxHhRfc
IunlkVns0GLtdJFQwBAc56m94ZODq8aaYHRVNIzW2cKX9/Jk11J85UDQJHjt1qsfpFi1VWyexCI5
4Fg2yb3diLpm3hkWFkR+gLr0JTm7TNubfME6B1NGsO62Ecc52/S7YALX3D3SCSYP5x6xJWPQiCMM
cc97U2fhnK6YGr/GTKpCwFDPRlgs2Xi35pzOS1jUB52zmIPP84grX46BHaTwLHkk/R8QDvAwaDIg
9qNY/a0PvAnEEyfDjeOSxyzTIMVe4euIVejhtqObTVwe4LpQS/yNfzbMK8yV9M42xoNy0P/hw+gm
zvxf/Rwr2TxSALsDc0a3LeibCiWkQHSM3bESbFfTKbcVumu3mhSbf65/7xuzzWpCPa5fjQ/BPeL6
Q7e42kXN8mRZ2HO+CZPJuW+u3RG20XExu5dmTTDX3pXzKeIuSu7CM6V7d70e+oITDHTvJJYhsi3U
EQMFQ7yrL1HuzJdFgRf6mwdpdeTpI9n2jThGp+j2UiyMsE0SLQapP1CsQnXD/b6hVrgMXn57nLS4
3YhBU6USyMFdKgi3aNdUWUOaI5OwT/zY2sznGZpp2RGBhTPife6PnN34HYmWikC4j0077cob6yKE
bRNxYMitVcOKTCa911G1jTWqkFr5CVby8wzV+ElkPszpAr/NEqxXCbdrK/J/YRTrTtk2IlEmmUMe
ZZWgaJVs4T5lWnXV4kyixGeIxw0OswHTW+9al00CAhe5+7IUL3jJhVWBvaMISxTU9/YUfizvWvfd
bGgcUiONX+5YuVyz518qaZSVqwJZe38wWA62DP3EpAeXbJ30sr0TAxHVwLwF1+twC0Tf76f8t0ph
3LOYlPKh6+zH/JNrJKAwUM4NP651mIgY5AUqDaQ4Lncon0UIXTNUr/MJcIh2XCKwdmLUxIjCOx+u
ri33NFCxBuJOKLS7AfWooL7AUnBjKNJvBD9OcDLYv6psdJP2nK79RfBeXfEGrDU/q5SA7JwZrzZP
gjVetcVULSPITrqR4QnExqtNmYY9QQpVqBuRZ5jFw2+fxEEQa9qOxxMl9jpFzR2WklsglA6/BXFd
w5qZE3AqHgGxSnZpkcHDYQct1XzJmFin+u6JZZN8H1MU01QvSlguhnOaoGGQDhuu8nPw22BzjSJg
K26kJwKL7QfcYrF7P07jjDTHgi0L3bDjYbHucgZYfy15P4C2NM9LHvaveWbMyuBcSCyVjtdMx+Lq
2XIH56TmtsJs8xWfBbggr/2QmEGKquK1wJdKgPw3vlUSpw7HsLcvH8cDEUcTyGIel6Ow+PWh56Am
pxXcY4Ih3GgoA2rEonxY9Zgr2QSpD8F3qXwcxOeMZRCGAwkJ2MZ7QyKJ3HOfkBzUJX/2gN+9LKwc
MQPsnHQbCKqbHgi1xMKJVtc+N+jb1zTiRnEAJp/JeF5HqQlqYFy9yzZpfn7vw/Fhtz8VaOtwcL5F
t/ntIB0jk/7t6xm16KKEOuh8LXyIepc2pL0HMhePeykXyL4zN/IEWXS0avKMLoFnnjNhSmFI0EHA
nBW+zQK2sULVVhS17bpqTOrhcjvZWVAj2of9szvspeDW4N7b9q79xihLqlet8ntOuqqNPrDJDogn
GznDiCtPqSWtqX5oLWLOKc36rHs1r6ez3RH2fVj27P3uQc+tRh/iPLyUciLd30Zqq5osPyrXyogz
ZQmWrxIvcpshxaBRO4I0HUddKJGCAS+B+JiLv0+zBjVRJz7eymoN+JaXv9di1frVIWsZIGM5yQWc
1Nb/x8aUCcHTpq9JOpAeHgNVwcbKOSSrk/VVQ4B1/imNxNqolEUfVq/pgmSqoYVQspke3oOyZK/W
Zs4uOEuFRIARumloKWOK+O/ul72vTG2Ku+jeeBd3nUu6oWRlqtVsjmFmEeTA1AaLBxUgQkeGs8qh
doeXfpZ128c40o5N/rPoCkQSfN4r8XlnnUSB2NzmRa87DOvU8f/u3U+5NzwS8NilFPWaadc3nZPc
s49yp63+KAe7ySIpA6H98JpmOBFy1vpy6XrhiMWk8Cx29wUOyLPA74UH/2q51IPyyHaicR7qKCOt
wkUYGCnwBU2ySCLPoidE+XHaj6KQCJTadL8nK+AHQeMUiitFMKZX72fSq2AfpCTCz9G2wn5doen7
MctZ6TresUt0wjSr1M6fs4yAizVRxRW1gp+U6Fs5R2aTeztnUGsdKl9sgOf4d2xZnKK7iVDHFypG
fOKhb/+mlWYQxgqnSr/gM/RsPH9VftKhDQRCtEfWfBEWxf8pHgt5ByaCeJIAsXgZ7Kkmv1kAcCok
hoB3R2Z3BYpnPQWiIGMUWjWnx7GyzbjHQUOMpF4aEw8nt5H0BvwbTq4648WpdW73KoG5xknspjUl
YwgeZ9vL8fpHoR8nneiOcMFZDDKyfQ+yyJHh9eMMNPif+zGnL0gsjfchXjwa2+w2Arky0Jmm4TLd
U5Lieg/shMABu+dk2jk5k/G0w/nSepwyLtvlNdUSlzIbOepZudCzrIJ+hFJx+L4Nn8GvY/EoH51f
AlC3WMnjbT8sItUJEWKcaQW66qqPmbH4PA7Jj8A++eRuU5zLwgdGFtoaade4q0W3BhJu6IFDSzBA
KzcG8GgCWom4C+9jjbR7YSOt/vKt/R40xbiEUjbIuKZxhgnmch3XPtsqDIE6iRr4b9cHyv5eLAQC
bagEgD29a4VWsjlTzylnaiXw0tPJIu7GA2VN5vfkuW0V4OIcvS9Qd1LcHLs64IaG/wy/SNXvxkgW
ziQb6VLOQMMq/zwzrgPIpvN9vUdOeSNsuL433V0dHar4u7Z0M/Gz6yL0hTq9Lgpz0VJEZ69H5u6y
rCFv4PyektuBeDG1bhpRaHGUVg1wv1dtwAHFaTE6iUO+ZKWRpC36FNauXJsbjp+8p/hoiXRWu8oR
Eh8P0tgAMdB8sfLygFSbmITMqzSU0SCNvTXnc/C2DZiq0WaGVsNd3YaDWqYJoGHeltmgmusejRXv
D2BnnhZ28WuwKofmZUBnKc5OzShelCpMzoQYLknWj6nJLwHz9l1Um5oc9Q+H4LuSvIFuuSKUaPOA
8KcVk6HFgyG98y1+bAUZF4rp30J64FRwgd5d/HcHP/1DK84anrFvTEGm2VqxllRoaU7uw1O/nQtp
ViVrYGg7kW8njCuGEJ+2DfSdin9QMCUSc2ynK15GVBcl3bvPRYR4aqUDExsvM5DU/1+wfY83cngA
Db88QQuboqTtGparGePl+AAaW4G/y6CU/aadLa6SzxHpuVF0R58i46fj9P+GMR4sTbslnE7Te0FW
Lu59MajU+CJe6m/H9WPeI+PWjRYtTFzMpnjmbvfw7fV8TOGZbuPK+TpfoRwE33l8z99AGVNmxAEr
z8pMEuPuZWa2cwn932TtMIdfU7V6yjhP+cvuSaX3889kZgDI2OvmUYMQjI0iyLEKQkSzdMReLf6m
1l8CJZBg9y7wZSVj70b1XFtqyOkFk3TNPLAmn8JEuPrr26TQsELlA0q/EHCH0WzIJWV47/1sSoge
0ynWaLF662zG9OIOYyr+rXJkznVJXSpIKb5oR1rI/UfkeUAzg0fVAstEDwzSrNcA9UlVzA099HtG
OzXd84Sz+/bkhiXs3zxoc4dWpEMJsQB78gEXG1r4ra8irqUSLp4H8ApcZhP1daeB+tQle9Dr12hI
lH6VSkncmBUJWaDSludcC5gD+DGUoRszoYImKGJYs8al4QmK8oA9C8m74FZjSFPnm6kHY6iAUmhM
JGdcuNHNfeWshDrk9UyK39qcMV2AikBkQWPVFfwhdUlrG2unN1oZqy6n0kWSLT408tD/y2saVl6q
FwrQTFFcS7O/vk6PXVlifxqpFzl6I1TOkouEhLPf1vyvuOYYmELqZ0pIWtEa2mbH77RUcWwgvjRY
jXdmCJ6TL6XckmIRy/3rzEUVsydDXzOzpFNKX38gt8qe3dpfdtWO8aqy8XsckM6HJuIim0Gttflp
Xn5jkDIzYzNLdeZkgNR45RGWrln5JUseT735oBzgBmVGiidYhrekoE75fJUq4tmMghAuMi9L2TJc
pxaelaI2h3U8QnaalPxJOk41bAywZb8z06f8sajt+tE0ihPMLk2YlJ8LHQKDVAacQSrF9yKPrgvB
ZHdPl/6xb8itmPuDZZujdXn2ZbefJFhhNx5jGFB/tg1ag8muEOLwQC/TiXh96sW9lITldSH3N7xX
X02NQHu81RTGdcum6iWZ6p4Cme1wYMsWb8Vi/nes6+21h14jiF1kChS0kqgq17C1YJHaKtyuUklC
e0Q6f34bJKb+4f5MiGPE3DiJ0wG7bQ5kYG1wlMEShCicrj3di172T1Lpm3UMMyI7ET46RKwvK168
sOe3SuSp3t7MY4DiDJTsDRL8j/P8ro1OdZ5OK05AbB9Ywf4p+42RmN99mLCp1RA2m5EDQ1JwvH1S
pWXvmVmP0h6FcoNRQwM/xsnJai8piu5Dph1TMoBO5CgQhaLNM9dunMfx3a7pC0Z/O2VI3rWxEF1q
3zXc4/Z7sYr5py6dVIkq5+eg88763dCsKcVS+xGLKwFWvhwVc6NW5bMMTb3khFIjNCuaNJY2nyzM
qZ1AYPvsv94C/7KBH7d2cRf5XtuwCyEH/HMTMP0HBs61EtVuqNkZOc3YplZ3iJidKjW6/31Uuz2C
8sWjRVcsmdY+KzeMFg37FLy3Eyr65le4QxwtIVf7NfzPcfc5IB3i6YYdlaskBxgaf8vXvooUq5PG
WxEq4y1ZuCIVjAG9ckYXGCXXNrIhDzJZi7bI5yeg2WnTPB53WF10LFTq6M3U78fb4r2EXWWA7bps
oYYpAdu+ccsKHQjRDp25WKHbBOAdAdqC27uobNFVLrz81ZLjhXff9oM7iGpfrXqB3/wFtXe5d2tf
NykRmEdmfiYaMAAoOCtsIp32LFsgbMI54OlMVSkf7XlqSwVgxzZcFgHYUReS2yj1zrskuE058jTS
JK5563oCo/KXEPv7Dyy055OAf9Gh70oQzr2laREDiC9z0AYZ+KZ645DPsz9ao7YwyFpermcS2iEi
xB/eOZPW/omXESeStwQAtiymiLfDixBje0BIQBYFgxVn0stvHvb6niGr1aE3QQEjTr3kaVVtN6Uo
eksVuFbgw6HdV7/PGFueLprtw7nX1Q2Cl2BWFgURw5K6TpYW5zFtIhVjTNPXWER7O3JQ8Dd3uXTL
iixL2xUxhp/3xQRm+z/jdqZRuNmdEaMp7zI/7eCjkuxod91rMaTPPhIJiUSp/aQZ84NQNtqUR6uL
Pf/kUtRHJa36pUW7LVzRP4iC6C2++YOZDx8yVqKF1Qu7WDmcu37Kla03VEWY26wUEnupy2bOgmMW
GArSgYvRQUJhUTWeRn1qv7lrrtMUXnzje9XWbLxdTwPPqVdFur9Iad8BZVtTs3U4ImAbWcYlwN0r
nbyPeCLKm7PQgGMAndWkjTyangVfwQrB1EhwvBiJFpmrbNh0mC8fqlzwKHev3HH7h/0jwwuGt/VB
zj7Zh/H0Hj1KLQ2zpuuUTGFAinjCCPNa+EBOKzWf4xY5hZX7v+0afQhczG8y8EHudPv6Jy622ZI4
e2zG1c+Iw9QqmQQi/UeRnXQs9FCNDkqZqppCGyiw2RxwBxUDXsDz+fgyI9gOkjAM0V2YGMHzpdyk
V58ZqIs9/nvyycHp7tsXlaZn+Cil+BYr4y0J9b1gzcsAmX6AbkAQlx1ieRLHWaYkx9f9OF605JWf
FKl9DcW+99GOEj7wWhzzFYjl+pxAenqKP5cFVkLZGJU2cOA1APU3X66IQq4PvpG7vadt0DmBTb3p
YbdAVUQEfH5dgVAEEH4SggCh9sg4J2ZGSMd6/jPFGRcYXP40AeifW3V1EW3cic8MvDCh1YnsFPaw
w0avlAHZ8+SN1O3fhPLbhFh5VHJSoxTKypXxj1gKIyE6naezY3eZ8BmHNIki2utdE618hDe6AxEk
ilb++FKgA5+XJKgGtOMjxXOWHivgygpATbyQia6EdAooHgkpOv1SnAL+MYD8jSA+VyQSYvZziAoY
YEzYEPlxl0REkUqI6Qp4jaqZw1P6ai6ddlRYSXXzHVOvzakQd0JwM4MV/vaKOxJDjSqvybXgSm4z
3R+SbuIkY71iLHyJs6Mig0QJGeJlm/DwUu2vEyKAkjqHZsOcf/FZoBZ0bljOTDv5b6PW/4CRXz0g
TE2LJsUR2uEkBllB2/GMHE+U21lCyGzA2yU01gSSWsx1chQoS64V/cRpFL2Tdvpajou2CYN4dpVw
acvizUEkAPRsmo20bRE/L0+bfkCOWBRxw6OBOUayqR6COEAI8dbt4TBpJ5b42R/WoxmoiFJ+Vd49
uA8XomYZk8XG42vqqii1hFcVwasuClV7OvnB9zkvi5Q6hGe4HDF1QqWSlXvN4Lv9Vf8E0ba/QeuL
RTh0j/WBUt5QXQzF0l3hTAhgI3QozugVVrhuddDGFqAAYf3AHJpVXKVp7bGDvoahpiH0++4cQCqf
IrA3M0uirQBten7+n/+nk3wJrl0Itb2HBLWOPJly3KsSpngLHDxEgMlwBJCjpvCyU5AObOI9e43D
3XYMF42cu2ezrqsd9nRAAEfZFrT7oO8L3lbmvQPnsBCEKCXVr5TJbFgSxbVEkjhR/Yk+J1PI/WpI
H18zFhfoIoJLsNb4GAHE56jFxJMmrZji4+4VklThola4K+NNnk/tjC5WQtp5mgXI1mL6H4nb/ViD
UE1u32UYN7Ti/urElrECxv8+mm9zuaL2LO9HoVA6R7YrYNHoUoP1bI93p7dw+8xYKMLM/R8GT+xj
LopkF8/ttx5xDLNiQH58IEY+MmVbu4JNo+6BDhv+8FDMq6YQr6dbxjPeKEmgqpL8ZvInsIk854QG
JVvrhVEBiL/IixZdRV3JBaN3wFUqfMLcdzAgliHO2eOeALwuIcTjP8FBoVhZ1cuppRuoxNQ5KPcA
CbfOxF1AjhP9riyjC/YJlIYjpMt84nmAA23der3kp1BnW9eKeqDTx4UiWj+kZCLQ6EUVkF1BDsnr
n1XvbGg/PX3D2y5MWMMizu9QKvxWt6CxFXK8vLxO3vPAw/FTZftrODHGRhlmg4KU25z4S1om/sHY
jFs+SSZnIsy13xwJ1vxnqn17JcTrZ0uEueGUnUiXzF3TeUoKeTNQPZEI5VjDBllSomP7BFU+u196
x+haIIdrozAMxJpvfSb2TUfqMTErLFHiQFe4g6sYnG47S4ArHj64/tUuevd9RqKFG5k0zZASBMFb
i/GPcZWLE4TcvSbffaMjjUPFz4vR94TN+idy4FVTgWJ+3Kev1jPHoHQwFqoCP3GmbOWecaywbuGx
gslKTzAzvvByFNmrEI/yoStbnohMt0sDistRSzac+pNwsmBSRcXEoCvV/7RCbRGFBYKd2p3Kxq5p
u8HC3IqgIzp8qxA8QKByFECElE/Mkfq2neDWey/KMp42z5XAqrBlq0PZ4Q6f+drfbJIXBeIMF6Zk
LJBWd8p+Pj5cVLivsslgciEm/NrDC12B7dlnEMxC1CpW8DEG2NmhVFn3Dwq7QsiJxyjpfbsRQUzL
2EPNeHwQTaY0tq4gj3phnp+dW2PvqyY1g3jbB9UBqn7qfEK7SHqJ9OmatHlrwjaeYSm5sgyHNqri
ii+9xJFmN1crVYxZQlqMov6nS57PWdRjxZwZDmG3otBhL53CtjAm4zYlsg3lD+3Tk3MUQ8xJLAKF
JvDF8mE+uJsA64WIW4for/iVWVBPeCliuNrx9oRCfkSRNlqijmtYL/Bp4b+TsMRDXAVZZd6XtoHF
k0RY4kYhtW2VaKlbibk23rTO9ErYtprRgYamLxE8jPPn6heVAcOzrZqWJZttrH+AX0RzxKBAaJ9r
DkY44Lk8l2jm9+Uqjeq+++Hf3Iyo3QsLkTKhhbY3ExxA++9j4jXzNHOswl4zZd37Upad9BZSPwDX
3TBYe6arTHWN4M7EPvOcZ57HFa5NAvhirnxsWtkqGCNIxiVFMkI2gQOzNdGxtlPjNHe2sQJCdasa
4hhltck/+XmfjlxAWqzHaVBqqHP1bRT6TlrgShYi9esdxJDyDgd3aM59j10wpLFLV79oNHYrsdec
pL55Ms1wHH2TL5KM1FBJ8bcx2zo5N+I2w9U2s277qBX2tpRUynCtmuARY2CpLF+JDqua2KTw3Itj
GxEpwgkwmBzzh7wtLgOLPb5pKDnfJSD2mgY7yHXmO1meROjq6TFMsLd/1NtyJ9H6RMwtFeFtXLrR
Y+R5/Yero8VolUWvOEaIikw6i2DmOnuGhQnAfRd1+xN4Y5E3i/dV8VhFBdeS3Ino4F0XO/KgeQlJ
l0SZgC3TAnAHFixRBX0x/z9vBliBC0knDXyQ8CKWwPz6Pw4vjosAYgpZm5hweQZf/npaKdSlsvXL
PI5LrcVR1q6xnAqqiT9i5bMYYKP+IrwtXnssivlb8L7R2sJ2uuyJbAofqQQXJ5aKFmG/ddKvuD3e
k75ixyY8V+hIAGJYiwBtBoGwAHHowL6QfCfS6dtAsE+uG0iO64I9lkPZApfma+ZT/6HHOFVw8KwA
PcB9y7Yh1G89vpjfjwcVDGx9BIJZAnBR/wOgTIqTmRBGnqFr3JEUpX1qlNvwiHyse5jvUopy1Fay
9vyLgi/brBsqw+mhzj7kaJhx5TwCiSivUH2SO4WI4fi5e2ePdYWbmxqAYSXASrGDyhvF4KMKhsuP
BR/P78cf9n4fAOqogTuf43qjDKMTaRAkIKsGBGDiMBNCjGfUTLF7De5J8j5T8M++hByNGpvyd2ky
Ih0G0z+QnSZYAuvWbSZMAKwxY9Bn0IeOj8j3ZiZuo5ZF1dOV2JWUI2IwKxNJR/5cOpjyVb1qZ5S3
bkutCi1uzu3wXnefnQv0pmCKJZp4s4tcuM+GzwMXd92j5LuGB7HqmPiQwe9xkgrAx49aEqWAqwAJ
yxhfzK9Q3P11YJvqRYlYqlvWKONetsTidi9J0X9uNtJ0zKGFggXbL6+NiQ/LOHVjmfwigSlAb/eR
hLffecmsnKzEa1HMjp+4wsLIwhnQWGh181ZqbtEZ4KwkpLUqu4Bq9bzIWEAfktZZUSf3heWJwLdy
yroLDnzIjHs47Ej5My3F6i4lNPihoInMeXcIk3UVLV4xJ+MrHSCDRNW4dPXhO+F+bQPfIC8B4IjU
7yq67C1ues4EEHo4D5++B0r2ENuob1ppvmzB18BjNudcCcvLrZOpf85eKadTcVcDFf6xsCza5YMY
dijJ0u2rM5oPHRJFAY0j1NFFM1mkRGuBym2Ni05CVH4YzIH3bZ+xr9vlCrU0b2sLXqLAGMeg+Llc
PRs0a5ESAME8B/04nFu0Zukc7+dziFrNMzBY6oacmgIiVFTvTNPSojrYiLnnfRyRK9FtQsOq+GsQ
YiwWbNvbNY/6bC0aNPXtsYG1kZs8sXNu2q4lyr7Czpc+3QR4EptUQVQ5Do2G194i41yTzSFprb+S
UEshOKE/LfOdowMYcgMJHzY/Z/GADeOu2DszA6pYtWQ8uLO+3/AgEyN09hdiCQ7QUFY7sWs8k7W7
qIEa+03JM29qoh0e9aLcah0iRp7ayZ+LLqxP0ZyJ2g+JzKzwO8PU6jS7yGUCPKHAH6fYSSPB9ev+
5pxVDHd/uSkYBpn1HdyidoJK+BicO7EiFOY2HIXTuSjSdYJguQxa30dJAnMnFYVinZtRvMDS8MOD
fo5VeWGcxiy6vyQLhYTDuDbS2Faf4gFiucvESReC1iuu/CdwRVq91+kkR/wmXAkRZPi5hlfjjAYk
uwc45GGPJZZRrvenFWwZeNTKg/921TIZeSAS9mBTuEMrLvtahH1CKad0YZz03RIQen7stI9FfLl1
wzqKqNRbz4UYkXx++EfQ14Xy78ZxbIBFuNWhccCu2XoKFbLD6atf5trMihAzis7NLvyA02Qvu3X5
iwa8ehRNgW2VnRIjjp5tzZys6KQG9AEQWiPl2ovKm8hH+SJqEDzosiY3iTlhrzAy7+t7vYOlok4j
6yria5A4DGw+kfXQMNs4ouWSj5MT7YnGDJFV2x5sg9YnAqaHbUcZPCscXPjlSCWzsCB0K1runDWO
La9ZbTAJskBxIdbFl+m2GcMVMmRVqtP4qO/ObX1tlVzExeo0AbtDi+HQx9e0hpQ8Qoq+jef/KFmP
Mo1vhvVB8Z2AcaQldUIk78z8xKpzw5NZKcmI//iPZJ/M3Ea08GwEjoKt/+lJ/2T3zLSYR43hZPed
DqeLbE/8ERxq6rsHzI2ogoLTKpc3mpXVHWbDcJS1Yq1keh/jn493WENQeQHIZ1vR7AQA/PIHggpU
qiw8bI/jFXzdiF9pmPNTw+n7RuQRlU7WiC1A2uNk0NQ6BIHZRHY+1ghlNLrgxhfbc8DhbzIsaG2l
sgmyXrfz9tQqtmiYPfv1eJ4XmJEwOfGAyLbtTCwlVlqn8CSpuuAxo+iKgtjubLZdhsRAiTWfI29M
c5Ezya3S4jW50QoWysaPs2/M1AIU7M8xS2IbXlhtS1bX0xJcZ6cDLYEYoSWmBypwe/5v5Gi/lG4c
1jbg6pB7GiOT40MTPdzMH9twHQsOWKps5wYDICQdDgGm2fhQMIhSLcWXNdIJzptc/vDP+7L11Yv5
zXGEAgX7t8YaSEMAq8xflSVGjyzJQnIwDl8OkSHgj+wMU56+PgEihL6w3AaJIByzqXpf4Lz1wFP0
Ky6G4F8AQ3RKXDqYeFjCmiBzZgLTOVRADFqfGb1QMotXdOy/ktJ6z6RXGEDyWFrYTuHizqmOC1Xb
pNvaY17FP6REvYSpL9RLs0csPvlFiexFxSGJkTjC5+hmEW1GcH57hO7h1CjbGxnHiy3FtFHA/al2
0tO3BN0weVBcSLYBNQFZ7HubMtwezqiyyqVMjo/6yMrtDMq6arbPn0xBB0HSl4UEZd8Jq+3Df7FN
UJOgoQoUBlU7r9bZJ3hFy/xft7r+wKnRW/bBZKt/XHIWUw7QXNYfAYQiqDVaghQx3wPWOLRbDXAv
5tjwJwRgnRfT9JgLnVon3w4vNr8WsgUxswjwhbVl/fcOZ9ql08wLaRo1TSq4pegSBS8XPTzn9slA
qzLALQoqRvZOxm9DFSAy3OBxmijyoZ/Lp28l/I3/l2YNb3R4PPWHHUCSty+dPHx+mvEJ5ZiUz1sn
tDZYTjadBHzqchz6Ezv/8bK/GslXz/apHR5TsvIfvl6OUi97vn7mgP3rYPTaO+bBgVKO/BCqyXN9
HVtbfO2yO8URwt3k24dEu1sDc/jJvVe4c8Gu28/2/Q+3ldh0ew1OSNhuPC1s8+Wi3g9ZVdzx6dPB
DiKtJOdu0CvO5s3MQ1qOeyB/NW20KpsJW8F7zGxyZo/1iGDdH3h4vbeQn5q4x2M6TzHqmHe7317Z
fEn5rL8rWbRqXca9i9eaV0MYxLO/JwgooUibLcfOd1PK4cKIb/ms+lytQ5CAHUiKupgZLAGDXtyW
LF32/jbBR0pldl4V8OLMakhNHXyZ7Beto11vpItY4p7Df4X0vWALwMC/drXzavwKzWX+dibkcs2C
yMfLGilwXuz42OEwrTj+VX47A2dxyjHiiBNXXMFx8reID+A5WDUL3IpJXCfbWpY/1HltmpA7Gv0a
E04xHG/0mtdbyn2wu1+PNqoglR1H3SVclMNGYhBUYOfvb1NpGg6DFxs1jJx3DcxQL1De6S7TCiDn
S2MV9tDkDkiQRBzspmiwjAhqWDvpqFIqLldTi+AA3q7L3VqSVKXGZTaTgaXmCBGnFtaI5IzXV2+p
bjUphMXTiwXLFGr+asiuOHuGait6y0nrunoALJm9MZal1PP9V4eo8++hQK12f7YgP8nrq9TFiaOx
nalmCYqUE4ilrLtjJ2qjE9XIFafZXHfpUNGSzSYZ/4huckloW6GD2VEpwgZZfPBTMgFWgmAr0lJi
QdemboTd7i7injTiWaWE/BgtCa65s3fo1gN5g6z3+6bi7sC4gnu1S94vxNrua4Ps62bAQ6HTEjSO
Qxg9+NH9GQp5muqLdElNphJ1+cP6C2S//a2H85r3XaMB2GQbzSfvAyQFIDq3Bn6xzM8/QxdPre3T
YlWnjiPuUUL+lDOVFsbBJKqy0ASMB1ivVjB0Nc5nspRkT8D7ufCFOPKPSxGTFTBvHcKQstVWblyZ
FsG1BIdh/yjXedAFiWfD4CU+TNDW7Beu/CgExA5VqLSQNlsGSAtmZh/MiGYrTTOSAYVrGXOq2DBM
NvViNe4JXjqTEgI2PVTrtsJtWFZc+70HDyRUPRTqgzA2Q6xD90lYKdJB97O0pIBNlbM8bP1L201P
Hp+Y63glYvkCs0w8WMAL/N58j1e8rLMAiHiIaUtgX2YCSevrd0VBFJaUtiRgO6JFny96GO/J+Iwr
yNn2+di1NVkvfCz3a/DC27zaB0KxZcIcKk675oTzVMyQaUIVoRv3JgkIQird3WqemPM5nuQwQ5eY
GHgp5f/LWVmFCZ6CNRzvbOpqn/aM2yeP/Tn3n9EhUrEopVDDNUZGGXgjaAMfO8wuuOZXFcCmcMOh
bKEi2DzS8lwM+0eXwoRzX2AuUlBoZjLuKX2sCIfMjwhJ2vxLEnDtCMgF5F67ssBQRLDA7qxHZftk
NdtwT2t9/WncTzfd8LHAY1TIqz699UF4XVFJllHa4b0bD4H8DFKCgUB1vxUZWz5xB6yGhEoZSsLD
VYYVOIWimc7z2+0u635mJe6W74gI/HVF+EjijxyHgoJuXEM7CXt0+/UtXouIU5Qc1+zrgGKuODe8
QFN1aRoUAyxfSW+UBaqOtPak5b4tIQYGsvOgMy8dzthT26AgE1VLxW/bbsnvlF8b+aNNQpngHnUW
ARbCSW9K+DANGpisSchcpj7TN2aDrhytAv+bRUdN6OyBihreUZmIejlN0Er20ZV5JpZsGIr7KxGT
7ltnzxTg0OYU8MJn0jEMuuwzZdXfELJk0udYj8wAiuEfyO/6fker44gDWULhGiKDz9Ia5ZhsbIDu
ZLKfAbMB0tG8lqG6MJE9K8W9gv4bDkGiauh5Bkv0BSJO8vHJEmXOmQKPODcWJ+qhbjSfo710nMfX
mDYtec8KIrSPByJUULnpbITTlEnsAdTVEOJCZIsP+bZRap7KwREr9KXNtPyCJfG5DIMCqBG2pga6
M8jQi9avC51jDqRKd75nL/w25WjofSRDH91iAePEe2XB+Xo9KYG6e1txUPVx47aUkx0l/rFea6qP
jtvtDKPSsLSoEtz+wXJd3/fej2pyxRfxqqKiAGx2zNRIkmYsM6Pq1//qN1h6xd50AKsIIE6DnUaE
0ofoDwSKdS+oL2IotnFP5Dc1A0pZILeaJwMIgG/mcY0D2v3PPl01DPOK17RgbqYUFxvPNyPeLMfW
tPp379AKFBuvPr4+DImHo0c4+BbH6jBSRF0ZQR/IJDe8+KPY1Ml7UYfzgIv7QlnN4tM9QDrjIRgY
jYe/3poJaq33/VbsYOmof9u90TAUZBJyIhQ4PgRrdZQWtt3r6LsKIFQLiat4OE3QlqzHmF159M1k
WMmyjYjh2Np7yoY8fEVBPe2YDRu+exEJAYchch0ia3F57Ry4EkC6kRWjm/oCbWgTrjaEzsVhJTog
Na6hbUZTNWCPyfXTe9F/MHCBR4Lzd2zwMl58UEbuRDVPmslVSYidfeTZIq4nyrPKe9UZwuRJXDYi
gbkDaqGxesuLeVC6jRWWvrVZ/jq1qz/NauJFf7E2FdYkV8CygZrvGhakY14y2vg0LlERd73WIFdP
BFfwdp4yK23iPRWf4fBNddJrskCFZVA+b3mOpCtjzC/vGdKeVhRw1oh2QHp5c6kBQgEmARuVF0Vz
2Iod/WUpTL2ZyjSKHdDQDjYpIpg8/Vs4hnK6hyrQBfwO1fcCcM2lpRrqd+9BoBCICow/wzwIaDyX
/ec9bdkLRxWuG8W7wJ2Q/cbuWnZdSbRxTcupg/bCYMkO7aQd594jKhCyOI5b7qOgLnaKoRKbeVpJ
+eu4W1mjneBmkfxjF0fAr+MtSEsL4zFjOkClKrPK8VCD2DFi/TnUOlEr6jaduGuFyIBoQfyt+PR7
oKuQQ2yOKxF4lqNHwj8yO2lrJnQH56FclUC00WkWf45E9zssaaVYLP80SY5GpCjy9i8arILUI7Rg
7ctVs3tirYJL+xTgoeQIOs4DgU++91yvNpiKMTH3bpAS36AyiEnV+uDWquGGjWCl1gwnvgxvGpWx
+QUlzl3GZZuFlUwsnlqwQ6Ru7+shf+2mWjXcgtQEl/EAZ9JP8R61GCDzGGGngQI+hiByYq3moG0E
jMCRVoSXxar8hLFf51K6Q53oQ433yn+FkxPLO8eFZBWAs3MnyHaHrWOVdYjgETc5+sChSRQKLW0U
Uchb79IXmfcXwHSCFb0fkZYf7sj+LCcmMzKGaVNHGDABP7gTpPTHp65RvX7pjDeGKOSuL9WYxKyh
B+6/g710pmu10zxZuAQ2N7OraQuRWoWSTs4CdLqGdkFHJRKuvehUC2WLMISLDVPuLdGaRCOqQqps
JdtZP1/JZXT462aMQFa7WRlJfsgtMDL27PQ+3dNhdxeot2/043pTm/h9gx06rUgx/FdDPjs/PDPq
tVJzEvD9+GWHC7Vb8d4jhNhVkA//AhiT3ePEnRQRyYo0lP04ZCZiZjgRPJkx42w9JedmruPrjM3K
m3f0GXHdLnBuc0mKzFCLXO9IvFYQFUNjcfa6xOZQIoDBz/JnuP9htT81FHtR//6oXkt4ozCwJrGV
Exc1tbwjliAHOnO+qQ+ca0XF7Osvsplnxkc2G79QH+VneyeB2pOpIqjKf3IAWuXi0RC7EmcAN35C
NuZEun0sI2SH2XCKXET9F3DSvJuFkqZYwB/l5WNPGE01ZpyAv7c/TeVwYE8BTztw44z4j4ZTyK7Z
z4TBXLXnjUVDLBWRxH6qOruIf1RjSGC/6xlFcdCTm5vnt1olNNhA1mtikIBGyS38qigFtyis9Ffr
X1IYXuz04kH8JkpP+q7cED9m6uoETR6m7rhA8zrCnSWNQcgrCK5AgeFZEmyj1ZH1fIwSFwW3kXyY
ct+NHIYLCBsB+yoS0DzabkUTWD3vPJRv/5n8GxomUGsR8g8d6ekX3Z/y/4XEWG2Fh3ImBl0AMf9y
sAzMb1onmJlGRKkeWRkpiJs3cK7ZkqYelEJ+o3aIMbOBbOAXgbZjsFhOQlU+N6uwPlwBgDeXbF/w
3MMokvJSHr+fn1SBIPqlZGX77Bh4TvUkx4YSGCSAUvI8q/13p6pRZmIgRtdOrqKoRrXFo1rsoYFr
QzkPdjuVahCUBVwlvSTJAPWuXiTKK1F5MOYd95qHWI9YWrnPeOBkQybSY0UKIepHNYyHdW7RwXEk
EBNeniOv75q+I4VAoKRdO70tsKtrFAyIlkLVgks3lDvBL4o8uvI/O9epFTuhS7b8s0fkYOzzwaLW
+E8Ubdih4owjaNhXPKVWQsEnAHMRlvvTgHMFyuBeh27ZmOhb/pkUo7pAwYwInYrOO4UD0Vp1i+PE
hVnJCFyCIiacfDapRUJRgiF+9bhV+kOl42/inu5WC6QHON94la7szjPMl5fArsrBgNVZhqQCBlUu
YSneCLZHoeEKDh+GI/zefoMjxqYlgfY5UVd8+WeECQDOveIuAVkT5goyYI6lZ9F3gBm+wffKOy22
IHqkXygJYnxMhZeTWXHHqO65A0Lt6zTSWypDdfVQufpEUFqirgt+GXD5ZRLq/9yYey3qall7SQ3L
D+ZdKQbqIZUwvZLeb3sIV92oVuQFEeBSIGylkh+Wr9Wz3KPVLYe3S0V7R65FbtU+WL66QmuMZu2Z
l5klFSsicNvfzMhzJul7TL9+p9KeUBzc0Wf10NYjcEEAEWfv5DwzJ6tRt9wGfcEqR1EUZbN7S/mn
kegW6aIKxMettcratiFE04Za5VoAk3igRuwaGlVcvi8Ulh/fL7E7OVObFtZNhcTKjDGWcyCGzumt
0PZ8kO2Lzntit5Icw8ya3Lh4harknTqef13EUQMwU3ojTJuFNwrMbw8khLo92CmbdSfAeThzxppz
DdkoqoS5UHYzBpe2Oz+0KsQ88vlyHdCNmrH5BddcH/C+Xay9JKgTNI8+SzNpZ+qthPu2W7g+DhAu
4jMyGpkxZY/J6hgvp6d+1UbgRQpP6y+c5Lqa95mGgh9/1olx4BFMxE6YEPkIdJHOINjf6evcZ87g
jMJM0gzAP+mh+ZWZUPK+5FABmk1G3N+tUqC/I7SPm2zjek84z94z0q31XbzIemn8eozIDth1LCHB
Ye7oWLUy6EKxTZei0hRgTeMr8EShnXxtBZNMsAj1GEu8VxC5VJnlj/aSKsX0rB+l2/6euYRByWjv
r4zyXqD5X+4KgR3WiTqo/IK2mbbx8I8cDtEcYzX4dLsNNxBiXlbbyNkhuxVwRAsLzpuIiUTnUp55
wgutT9O8p5AgnZ7WiATfaCAXD6a/e8S/rR1TKaxyVI0Y5bOjyxJxqcjN9LqZSmHBNBkuiFBUzB7i
YE7eS0JH8z3FfXsDD9v8nOI4o1aX/axI5cg/Y6jqYeb9lpwazSlY++E9qNHPczuuytLUIhyalnKV
eJQTrphpU/z4DmzfQX6ScCVdBSc3yyJrWUX91VaGa++4rKW2ABdsPeahItUeQLRN82OORqu57vzK
jweiMf4u7n+/k++HsBPT3RoGd9PBmRSyQK2/foRhZBMwEF4v8pdLXuJZRcLhKpuzfBdb/QBl6Kbv
hGpk/PLZyqdDntNc7EHR1DZ3f1urfwppxmcJ95mrX4i971OrpGZi3ujcLpd+/dIlVVbhbJSh5Kle
mJUSc6gOI2S4FXWUnYFQEKsAotc/3dHWtwtPWhgZqXoxzh9Ifr53cWUz9l7BS6Y3Ow41qzkOAR6g
bnfoWHVAl2CAykr+m/lEANoI5JvTc6Xh/0mJxvu8qKMsfBJqr4K54BmwlG4vQoe7lK11XMe5gp81
DLavR5ysYTNQ1IyJkRoCI/gFThM7vUNtZf8AgSLsKqINY0UzpFhD+3s8qS8rbf8m8ULGi4Npfxvp
n1A0x1agE8RW8Jh0OQW2XWXC7nCuB3+Ox7RaWRU1QFtzclXJtn2ZBqPWSXyXBAVHKfW1yahfWo0j
dl3oKbOw2tnzZwDtFlNRBsUe1EQF1sfbTgSTGXlx54Y1tlru+3ICgtSD4ECqCbCdG0or2eqJ/Fq1
kq+mwylt5L5nfs+Xf4Dc5ySc+pNBVbZNVDvxwh+XrWhQU0jAiuzi1Dt2RRjXF3NC1EuhlmnC4/dp
bW3bbnBfTVHM+HM8Vh7LvPgB/qorY9X9JaT9bw7tCEsn/mJZ1V1ijbM5Zmx/QwcoxZ6EjQ3PyvL8
jlAzuW4PZmlQAJhRzi+Yp1ognzifKGgbwaNR9OJ5I0CdN8NgNQ5DiFhMHQcyu/XeKaS//wXLhAtf
5U48ML+OtoK3VPu3OuOezs5SgDkPXYVTgpkWocdEyTgADZ0grfFW4K4fPoV36C9PgsgtIj1qkGOL
FkhkqvB4m2Vw1uEGxAj9nDu3ZnrueZ9sU6ZpO86wluL00YdaqhGY0dQh4SNKVp+pu5HJiKlsoGyL
lF1QH3bP3aC9t+hR37KP5dsYHcqahyEy5C79athnZ1obc6wJtO1Y6cwjgyBg5GSgWL6J1LdLz9zs
DSEAnDKbM32DCTBaUYsh3NtRiAT9BZxeg0U1MlkVo0q1IQX55me+ydg5pjz2B0kZx9Xh2mDH7THw
VzyYHgDo8N8/sJcmR19VwXDLMQ8I+BNlHuZ8thrPSCLB3fS27EMtVqcaYHq6mAwrKsF+NcdQL2DR
3+RrMU93iu3rP3t8C2Gvy32s7lCCNzsl7pXQOk4Hiiidw6MI91mjLcjqMXLc4AGnhOfyh2PH00C2
L1aA948CkLwp0qnDNv/SARnQspFP8o1wEOn1b9kfF+M87TGBEVcPQehIaPclYMPtLwwzL2v+/siO
17adrB1+R/yZenCspn1ocsha9j1/w1WfC8s37L8rWq2MLxft5Qk9TS3z/xjDGU+isdJqowcFvRPH
yuMIPBJEqAx1i0O1aZLLfDA+aUZjG/JIaYDAn2PLe5iGUrBQ1oFjplVUdjiuWPa1kE54b61vnMa6
1+fZ7tMGhSnLY/fDNj9QhkPyufENG0SxzhIVrW/NIcF3/E1tBvyPyiG4TsqCErE40yAfsBkaAPzl
NjL2dIOurTG3QBW48MvbwvXUBprXSXJdAdi54FSUI7rSwVeO3/K8GN/3zdeUsupU+lGiuBv7Mvxv
VZvAeOx8JoQPUF55D7id6YqWGceBnyLaATQN2k9uA/jT9j6Ar34Urx9cg7tyl9W76llMFgJznkI2
4CJnbma148mrM7CupNAMB00ZzOrPQxB33bt3Nl2N0zgqeNrvL29DnVyC645vi/ef1PVAQECZ78yg
TpDrYIPgteTYsARdPSgIEvFNFOEjxHKAU/p0TpXeed4fJaYctml3UvrgLuHnfjn+/Sqk7eR5COah
VuEfZwC5o4D9a4b1QHAJ9ockmp0zJJbFvGibE0Xumdgkq05BXD1MrheICVuQPYMLtZvXDnbUluZr
Ukq/H1EqQyjDsmqpk4cDC8X5FqP1GdCPq98KUi85R5HA8Tly+GdaRvqA5XCuUZQ1dV81zBwF0CGY
d6DmT4XyesdARMQMpyRBhTANBqsFfaV0Bu6/hMMlR/F/zReSRLoqmMbDrnicnZ90Aj3m2tvFPwJm
I2t/tXPHqD72xqsWEJHTWx4l/kD1AyavcWUaWh19q5YqP9lVqKD9LY6SDq5z+km2Eq+dTzChBIPm
NOhZcUiEujQ+/pSGGBnYlEGnsN05Qwkrt76XkZPLcRCaVv1X/HK43o8Ibhg3LlGJe70U1gXcRCcU
kAK1t44Iu71EtB/XRlKEV0jMCFfwYn2XB0ZSX8SBNHpEIwRNYyHNp5VFbb/5CeIW/DeY7yPswPPb
rJtOr944VkXfbMUsKadiujzGOW/WxeALEiaJfgqKPprseaJB/bOyoL354jGZzpJbQFmJA005zwb9
YswwAvJ//3YD9YAgr8cHGTWzyChIo4lUMxjNl8iKMkvqS8iUOJjpkRwC05ufWtaP6rdSwlNBMUbK
wbTRHyg+i/S3xQ3LKV5X0iNrX2X+kqFzvnD7G09bKQ20QdhsXfEwEuVHWXHBH6br/UBcSw+NAoy+
QVKImrRX8NkslfsKsj8WCmLBow4m6o1MHnizDVF6ZxEKrfIx3Xxq6mC/wmEOtqpeCUYvziZXT6oh
KFCQ8PMEF4LAiBofMSXt/57zV4my+d+hkjFA5tl5Os9e9mw+dM557oR0KHwE35OG0kS764M3y6ST
KDCNxaAnLiWx+pj7tR/bocBgR3iM01uEbbH0ntefsdcPko9uWx4FMqcCfUAq2YHZINA60JM5XXt+
JOyBCv1i4Budf9r/MC+6HrAjoTXmUe02rQw6yPSTjWFuselxS1XBv2AB3GXod25CQ3OEAN4uM0EW
MtoTQ0GGhRTZaJlz2geMm4DNONGXrJEb0Dkkio8wGBp18YK27YPwe5oh/fPf3kGZ7V0O7RxSwIa0
WZPZg/uHoNLdlcw0o4XizMD8mu0Ib0bGgDedMNbXxYGGgISXM4WR90/tFRS5994GrXISm0d13nTc
RM4qQ9D9UrPrUdwIJeDEISt92Do7XOwSvW7FRj/Svh7FHwfRWjlo+ZuJ8QVhXNLmqoFnQafOHHtn
i8s8je48Ubc5cDgrKLZIj5VZsFYFElu53AVS8bX/p7TBUFtqwWKZhAKEUZqSE/EV5qWiLGZ/P/YD
IXoW7Sa145r2ofKfzRug/2PY2lkDvEBYHJiCqh5qxXGpQDdJt0PvTIWq5TRupufB++X4hGwELU06
CtrjnRmcYwFobS5P5f8URV5XJUTi36Q/sxUSyah3rzdYYyw1dh0tAiOLX0LXCeCJtVhUsxMDHZPa
olwZ8OFi+sYla65zg4J3nhCV4GFVJOOmSn9rtqG/zFUBdD4uqJNPRXe1ygaD1RlYsXkD73bjpCgD
VxoXMo2GprbxJEz36qnNqSoORUaPvYobqA9ePrHRMpZs40Fpp5sj8UO+t6V84J1mKuxntcYhvlF2
kJwYvqAii7r6bRkQmT0OUX9kVpYttvs7V3YJaL8x9zPHbwUXMRm5M1/GDBqZwM0GPjHx2Y9utBYh
uqvi1NJQ5PTnKbVHV/K8oMxGSk2X82rBT7k8njJdnmklkQ3IfADby39cXn0PivknTywYwovJYs5R
1w2A6sm8cm/i4X5i6YtE3ScyW234KXJodCt2myvUuus4eg2q4Op5k7Nt63wPplm+79NNOqZnauNS
tPVTOjKa5jh9kZDF+l2Mo+FsqMuQvpbTUYcKPKCmuMw4ba60aexmv5Ybv1x+VeB5E6BV+t4N49Cq
60HrZlr02ImyaM8PlWSbqjtAi6e06nNUtDyyTUmg3bt2qEXZyxltuSE4N1iJJ/KGdzOStKUUtYQs
7LGZAwUi7pFHwzD8Z56U2qvqQzJDrmxZxJLc/gG0zINDhpYK/BL/JdMdWrPMHLyUr2z91rNho0U9
k2QR5S5hJrXDtk/PMVEk0IdWmhqBrA7agiOofbcHuMIy2rwkylwhbuKMnpTIZX4gEl4YYDSLMer2
r8pBaqCaLReOjxyS/SYKIjo/Dn/0IIiWpRCbcPJrBNA9d2Iib6Lv5zqHSGLETnrEKhgDHZImEJA7
+/lUHbjJokDz9SJkrO4SdNL2UY7UxXqs2Felgx6PqKaqz5F25fDAsKf7IWXvISKHVz0t+XpuISKB
aj+C5Ggnw8DDQqioZk+Ie3CGWXfFZHzn/D/8Q6uFa2ipGu9HNZjQTaM3qSNiWKYdIpi+j9gd4m8r
7Cva+OnGnjKZSwl5HzJmJ34g7z5vyC03nVvaxT7dUGdRPM94za/yDcqdxEQz1pzGH/cUh/hVzLGY
m6EutfKbJoUv4BPJyHpcqllJKmMaogSLR5H+ZnKoMa8XR4cAR7qzSj1vL45S02BdZtXPtqTwkvfp
P0/WK962WpEidOdq7GPfUebyDXgZ2QPWVuX1T0056HSXYKwteSw0vpL81UlfbhWgaliyD+kEtdCK
j5Tjtv28wxa6eY/0oBym9x0+1236OzsnEkzSK3bv3MEgysz/tELeGr4eINvFbqqYC+zMtFTHHxRE
Peg0j0ZampnWC1GLRlHEHJMHDKtCdK9dVovnL4NrLMnj46+QORnpHi9AQZep948Dob6YSr6xvU7p
lZI5dX8vkLqSzMXF5oi2F3xT687V42qJA+thIgQz4I4r0mnMa/PWEhD9YQD2uxLI1e/byu0gFuuw
bcMp7Ur8rMm0h7WIVuUF8pqHYPm8EIYmAfmaOlV7rP8s3/6EdMBOYhu/0lLFYEgA8YjvXpqm0CKg
2Q11qV7BbAQiQ6NaDGauqzkb2qk256quV/8dcpxNvG66E5t4NppzPORZi3H/QwXtw57Vuw4KVG7n
1ZnZvg5X4EU6Brl6XzLjShVNByGZ0Q5q/mI2sJt9381VMi2sX2D+ZFJDFUmeQWIOFYNlfOhH8klT
VZX+ZBUWscka1VQPOmm7Tv7iA86mnE+JaJUhStYDjglJLp6iiE4wMhGvvTDKKs2TJ6OikgTfeBoq
4TwVN6iczLxdtZ8RuGOAY9vtR1yxbKf/Wl6XuQvvhR8juxxgejdyN1JpjfnurYVpBwkf0F7r9udP
R6TxCq02ryTq79XIr9mmWAqD3HgdeBz9R9hi9w6O/kqNtfjLfw2tSQwpZww0+FC0puXkgYDJo0zt
Wl9xKKXpiSEan5K13OEEhNWbV7c1yedSqnRDRNgfcNkYBYlC1lcGCHkp2iIp27aiHcs2ri3i6VAb
GMU2gEWKOTPJSmgkcz1GRN4rSwZRaZzrWmFghAlnonBG2S//EI5GfVu00VBjRAkQ6OCoHI2oLQSO
DoY3+ThnARa5B0ep+IUtAN5UsaYU0YqLl7tPp/lN24Us1GkEwI3YhkU/Nb7iV/6GDfsINaitdGlL
WMdiPJ2VrFHkNUxSKUkHJdv2gJvTc4Dh8s36zl+Fn6dAJUerF5CNePd6bSLG1aFjJdBDgyk8JuQ0
bxjyIFi7Td4cIRzr8DLOsL3yur+U7+isDRHUc0kx4vG29K23jQdTXLfTHix4/Y/WZOF9AhB7FkRy
l9nngSuef+aEeLxK/mj1UXeiyn+sh3vqs145ODv1LNpEKEACx+EBzQlUwirTq+uuECpnt3i+kI+8
WaRK98IjR3Qlz81k1CvuoYCw4Qfr4wINdHtrK560TD6HrULdgEwj0xPECPP8pAHNXs5tacVGewHP
h771nkW7OwolS1ZuQRe6YhUcnJ3MSqnNLkbRkOGs6fgTPOYSKW+iP/XPRi2nT7cxrWVXl0xgyVLX
Xf+GA0AGLmU2mDHFby4Yz0IFXETXsDDX3SE/m1QUCbaPYfg1M3v92NAHb4Uxan1FcT1w181dY4QW
bHfT8BNU/VedERUrNVMS6Qn7kb8xAGqisILpii0HMZv8oVaGXHMeXDGsoHBKahRjvmyufwdUqJsf
ilKGdOeEc+uqLII+xTUH9ZtCbLqp61E2bzgCLCOlL11pFHFcg3HexxtXqxbLUDqCoHMKtwfbGi6t
NAwZzgThfGOfIxLc+gYAqJvK1yVsFCCKD1JkCaYzHJWB6sg34FCBbhHS2+quYfB3FnFDRhRl8W8e
qf0TvcAPYO4HUta7sHQEQsRYBvHBJ6OftBCYCNaj0AptuuE8BwaGoEJggp7iTxjnmXB1PMiTAGz5
TV4rIqmCxNDYTarlh0P72SOZwxt/ZizQMU4yZPUUC3H8TOwSAbl1AJxp4Ik+cwyUC0KejMm/Diyh
aQ2DNO8rLylFI0jrwiSayfA4BGXVe+JvHZh5hhsLgA0MUJgdWcdgIeiFGtwZuLM5p7BRi3Eowcad
RiWotRtvIfMA2+j2HsbdL0x4nNfCGpeRWj2aoMNXgiRuQSauy9fZXAb48F2jOFCtz25nOtjsXPxD
DfByJ5kaXa184BC9TR+iPlZyS5ma6ddRNUJZjmKowJvYV2m3aQCz9LSvBGWb0u+1UQYphYP80jj/
17VoAn/LO7u/pQzGY/SQlpVtpLLLvTB5wTLgDD6iHbT2yjzdJFCqyjh489PNHFGxd5TtEBUTX3Rf
D1KbkQXDTyYTCE91hW1iXpgIKwCgI8uN/UdzFW7BMNMMno71Sfneczy8VVY5kTWheegGs6MR2BjQ
UrFzmTz+ms83SDOFrJUlcRz60wA6QbcZK/R1a8pE7EylLyohB28AZRuH3Ik3X3DC2Vtg/UHGnv7p
3Sd1nfUqjuPNV1LG0W+Fz//zUmApua+CwKW7Pl6hI8BsfkgyDbe7iaKcewAMmxfX4IPQ6MYPve7m
wo4j64cbp+a3jfqTDvygB5Fc0Ds6oI0r6IxdbjVSM4QX2IU3XHRjyp8NFrPg25QKvlwZxljIKDto
DWsL7uuUgTXUdpAuLEMQypOY0rR6GshwNoYIgf2WRfO9shWpGfeGzU0P7KdxILlSwtYDZ+v84jdQ
wTPMy+0/ORQupupQjYr7F/VVi98lE9YquMqOucWEHpfGu8xPcgl1LGybDCMYrlA0L1YdVAE0xld5
XSb0CArRv6HAYq6sOQ5gwHYhRhA9eBPgX5qfDGRZxBI7BXrDvAYWwoZ3JnZIstcg05iPcgZOu1Kp
fPwGYTQfekP751YmZWn0NX8iNdEl1Zd8chcb/pysVSlwoMKC6OMyA6EnEzoP5UafZnDahRsYAxlV
deelzIUFivd0focXGgVqFDibpIWlW1Z1aQ0pRe44cg+KYYKG3bQONQdtlibHgfUe39w1J2iTpKfk
c/nIzKSoniInybtHxysS682Y6mJzCL6u+zJVcLyUPrA6DTA3EC6Wk4hfdZtIndT/kzD2hN8efVE6
TlZmRzcH0/v3kMs2og8BlegdzhblrAVNp+zL3JQyAKgmDRDfYh/Bjjh/dTZEtidK8/mAybV/RVNX
TQVfhWv1or7U+z2iBU8s/pKNYUqeI2hsk7MIkzRvFqPWgI6B2hqNh2iG+Mz807eQeUdwyyBMlcyx
jESlDY6doXgGEazmKu1g6X+EyhIOcR3TUq7bi/bH5OcNgvDHUCcDFzDJGgc6S9mswuFkRtkR5rej
bXgS5tvwQhp92S20hyrZkec2+U+Bb9/NugjZ1nyZ2dze+q9lCB0H3w5a9zjzUWY6Vu9oX92d42mI
uk0/THIiDR7RhwseSmF0806yU3RrCkpAW5iFfsa1jNbYksXbd0xrHTTL/4Po1i3qolrHBf7sMhjh
S6rbg5l5cDzDPVOgxxocQzbEhVPRP0a5bv4lTzJ0xH396I80BEIYUQr2urpxaXqMz+IyFi3cg5+T
53prCr+/d5ifSReoZ7jiH2mrdU2t6WyEdfcVW7bLvEUWIxuo/74Cvz0VnIxGFhXvp4Q1EA5rUF/m
79YKP8RJnQhpdNBoUkJwYBGQORk0+RRHb4Oyap/IbPE6R2NrKm0hR6pvXT4qv5ImJNeBtEhPd2ny
3aGBiVniryG+alUX8QnHhMx27yrlzzBLX0AFcBGpznPbiusH7hUmtZo/O/ZZizOAFpE07eD7ZVE0
3w3eoI/XB/AJ3g3s86gw+rsemp7dHb94mKq6nX5rxXa/jVVJlvyYYBj0eW5hJQ5vVcAScjiIwici
L2eh4JrTMwRlT2YbPMvnqCoOYdBWusmeUCJtmZ407XzSb70RVteplkbwf1a/y1mHj5ftvh2FSMbE
E48YqwLdP0okZCSqZnpAm4Bb8y+2b1N8cGAg3kWC6ZOBi3FmYzc5gW3dCf+C4eq9QnvigZBFnv9I
F73d0Bf6g/L2JKTRNObEjvE5JijwcXzkJl/u5f6PfHQZRRtFJRE168TPKed4wTs2EXB2fSNQ5OTD
VAqDpz+604aF2rhJcfpEDxyskfn/3lXOpwaEjb8Yyhy95RJ2EIiTLO/HdJbUrZL3jCOdtXazy3+3
CMlWdXpaH7lPqssiyaBIZu0Tv+cjG4OHYzhsBCnacUNPDUFyygb7tfuAernHSx2FdNmi5OhGQIDf
+uuWyBsY2793weKTPeZhYmoJbVtRNfPnhBMT9EK8S02rjVkre0Nvn6lB/9hscGBYeAQVHtTGiuy9
rG/wcxrVO12geLRoczzeCBj38z+L8XBkKR8v1FqVlKBF3YS8uWGixAo3k+/V0U9jjWCdUK9MMrg4
qmdksRx0kJyWMaKI3OCLu9V3+BAA2LAd6O5sdMyWDzmYjItJY1L98L6N/wzWz8MiAmQGIt8f4L/o
i4bjt2du0pgHZWZoUVz8Qic/P4lemHbXtwPoaQo71yfqGGTwrjNTehjfYoSRNxuWrjmwPFAb4+H0
70guk+DeCZHz0Ldwfwd16rKnl3nBmra/W2uFv6+KsTmbH9qP6cRf887vUII3naQJ/4wS+bSVK3c7
PJ1Vk1tAzUcLpdKZxssyqUKpUO8miyzTRHWuHi0I2YJBMUuSLy7cRgUs8JbuJVjCAPiPdVj/TFZm
rgUYE3y1SFfIV2adWj+kJSM/tPnnMYrBSEHqlG9jScXqC8OHlbtVGArM93NE9JMxfWQxNE9ZBqun
wfVk10Raq5KUBdJERYahExzEdf3PuVsLmvZoUkjO+H1M4qIwD6eEVhVYVH72mGiMcxBJ35ztdm4A
yPiTbzgzH/RmarfQeIVypdsQFk0iziYyx2+ZXopqFrBZVmpOnj1dsmoQ4csYBpaFt7GPOH/Jq6X8
l4irTfWCsRKMxyVG1UMADmezgf036sRVD7d7+KXedCTiaiTqNsRVEVrxkkuiVWZFcTyROPqmjGMV
94EdMN7lc8I7KWChRi6Pzlt6SDawR4+Lyg/4zZJVSq8ci2rHv7UYgCWub8+T44ucot3J4aKeEoJQ
q8amR8enbsY/6AyxKN2HHl4nSfS1oQ7b9lzS/hVFEAVu7kCMnmSsFrTCRmFL2JY8nLzYQT1nPMto
XlrjzCU3D+XoBzd7PXMyiTwPNUysH7AxddqlqG0A93XzvowTmCy+2RbCTMQRQWbeGIKBSmQh/tCy
b+cwRgkaBIvU9j23GldZ0v+wR+/fu6kqhSwMRrhWf00Tf8dOx7FKC4508Vtf1vSXxqyr4uKiEn2S
Iz6zibKhx5tJP7CmTE6aNajvCwTnJDRecJNTgshMUYp3iQJZd4ujUN3zRHB0lihNBmYaHoBV3hxV
yZqVx1rS4/3TPscEydCtlgdNTVKcFOZ+KtZku7U/J60eW/WMKizHqcce4Lb7vUP6rWYo8PlTXBLn
QNYn0Ru4rHstCzHfNeS0lsccAfOilC7QY6/38VD5qKwlBPYMrwzg/tu9gnTrx4lF3zlZJj3yZnrM
RSUb6DW6XVBf4G2dfSFJhi6vR0duHBPQooeoQGi63xjU+lb/tvlQqggqSUpQ91sCk/Lk4HXCELTP
ZpS6/HgGHeR8goBDCzGfVpY6MI3enMMUTR/q5axF0htXFOIdfnj2d8UXyD1oC0WXS/kE8Hrx0x59
DsLEOmcpBlSBTRXFEKyUnim9/qI3SCBBqL+6FEP99iyjLxj1EeGgLCJ5IqBp3zS+YgdgAxYAPTsF
o5YwNww76gRhgRIpH52+8IS6BKqus18QlUPTUFGj2Sy+gy9qLNCdOJrdtX5xACYqAtc0cKv9S4Uu
NH4eX24mRnx+rj8GEyJzf645hwP7qzcrBswmcae9ofbYlNwfWKZxvLHzTcylj7ZgTZ8FOR6bmLyR
8mNb+j804+UbfXZjhSpdrHOq/LFtiBKgaPwi7dkVUzx76ih+MSHrlrFSpmLt62ruT6PCEODVSmCX
EhdVhOU3OzGMi6L5Uc9mQi0YdHiQYZWrOcMxMeDeU0/CJ89aX9wVnLbJd8qOBxRDmqJ4xrRr8WIt
Tz6ELb+F94cyQEacRjhU6DN7Kqc/k+c95IM85cR6l63LxchVktg2TG9qPUyrcKryoYDHqXEpMgGz
t1no9syAr7SU+CsHYGM7862QjaQBueAw9byktGaU/LZ9mw3i3j/kAhNcFVfbSPf7yNALJNg2Dklp
KF3/AECqfXhd4LP6YErZ9scrqcZoJm279fF5931oxWdH/ufQqx5mff/qyUweJv5PNRPTMHoudxSD
JKtkCkBH5x7uLoEvc69XvEAlbcvJU6aqpw6cKyAoJYLlynNufcA5L+g4Nw+x7zMu2g2iz95fHMWH
EIz+AhAlejw6gHlnCce/ShXQHANpPlJM3HUw1k3Z3bm2pMrjcwZnz5yWIZlN8cfStZsQzFF1URkl
KHmsFk0aD9qCSRSgwrelU/FIvrG03rlCpC2Jt+CbKIcYUKAWkJvl6zg02DGORDrA1Kq2IxojajsI
WaL3EaCuQe3jB4GToCscBdzY7m4dyOyUNadRbaX/phPqBF9BQVYT9usk72EalVekdVmgKeumrCAV
XALpcYaLmYkvx43YfTLADASaQbTTWyrFWgXKi8IuvRPzuXmVvk9/m/9NP3ML9O+cxDpAnU9vkGNu
kVgSJ3ijEMnX4ys0WC9ROWxg9Bh/BhH1hzjsIi4qbl9MzU9lL4c3pGvdcIHF6q5bQxC5aZpnqZNY
QrhRbclWYzatNGkucwYTK/Qn1qooA7A2uPOomlF01xumqKGifBAuSLfRmScSwnMjkBGv2nhyjf3K
XG/IprDIb2UnaCkpgSUDxdDgnlkpHu2IWg9Ss0+gNcotOQjp0qyfxpuLOh+I776eXLkDuiWsbchG
Dd5mVZtSr7KW3Qr0DXD4+cUdlyGd4FBcYL0CNqa2Drd05P174F7uFWKdOdMT1/GosWtXD13ZX9gO
H5bKXPenyteNRqwOWR9FUBljUfhDO3AiKlOXwTnIr3I4vsrserVJrpbbxl+aJ5BI9G6mR1KAQHT/
JGlWTYuV0o1ySmU4rqF58Lt0idUVzfIO4smRYH2ha4hrfMUdSV/fi9LwvqkhFOtvtkKHpqVeogoe
G2s7ZAvHJKZ/unSaTUZ6Co/e9oilZdBYraeD5guT74gCcR1BFhWpSb1E3Bb4EPTvbeSiVHvimIpi
772T0YvvPon2aCOgDLMguvD+nxMxX6SKZydRNS4MZWjJAUkoeO+/H5QZr8Npd1IQ6bBkYrlbmpNP
001ZGcRPrvk4wZYXLvkiosTY2lSUtY8FfnvO6oRre+h6vaTn96BpVeibD/MMCJE6kpT9L3jQE5ZV
l5asFjBGzK1tiPFMPquZM8uHMn3OrLR1bUQ9sXtKs/8sIsNW1nzz6Sl10bRc5IlJF1ce73HCnPzg
A4g39XL+UlcZrpI30x4UajT2L+ZW/s94hYbMc9iwtrAPGqUlva3Y20lvt/qqORidEPf00kObKe7s
0u/UYnuXmLYBALoGh91k0RR7TNvXPdphTbkhlLuO9cOnatMbDVcXH5RKLi9GfTeFkB4ZmDvMtCoA
G81J9EsV0D7X7TM4TLE+KtdHMc5kAq4uaTzhhgIiWgeJPZHWsSPqQMfT3KAimTmP8PPN+IstX1pT
HH1fquiRGYogWU5/B4nmG0aZcTp/dDG7iDozkmHgmrf5j+SvC33g8ruTQx3tiXPD/OQYsoruwol+
/SFlgcygvsFzmv+uNbLBAQxjB125gkDqYQY0bD5bGGMGwEz3+S34COoTb7eh/kSZrmdrprCJm0uJ
qM+PF2I9q8Zt0AlSGD2QDoopy9IJW3vVsEb9RIVX462fEPiFT5Mn2duqp7sH5rpBUSG+5etdwCPR
xGWigajHIr9ZPK7vzbmBjtUJB27SNnW1FuWYoB/oIIHGGJr48DZMeGBNduuj3s4ciPlP58ghOXuC
8yjP09975zZ+L/NJIQ/HkKUZZZENlU9EbRVyAiV9gGr88zObk4LJPUr7BuqPE0kNj0PXWhVSWImu
N2TQaZYEo0d73sK91KJDmrlr11CtEiCps8MXz7c+7v08fbhE93oTIvM5Tu89xB0H25LihQ6AINcB
z7PEmbyu6PBj/34FmGnW1iv4ViLxnUdnBHF4GuCuiwEI1EiR8vCc1qgoBBTstpDafJ6ygru501pd
aMGkyS+57kdOloF0KtocevNcnIA2nrIHvxgcHMMAqQjGoEam63CUlIG9sEaPqYaJ+i5kfGsLcSwr
iS4RSg3NzgbMahZW7syHN3Yr+rj/BCV4nQa/NRmM2586nyhkJNdnVrtR9m5P9NP3fm+r8qrTCDx1
wPQBJVv1Ct1mYa0OP483KZCoESB2d/8WijiojpWMOiIhuGjCEfUw5dCG/39jKLFikhPnYEWT3deU
B0wjZbnWXxYy2wsyjjPE3kYLdIWcY3eOVhvHgUkXkPtSTET3/+Vdml5S8EOmOTnYqRc8m60bWuGo
EFQ3uSoPltLV17JQy6oyfZ5QPYElHwAVqNc2QlvL0NqZa+tKj4ec3kABemQvj4l9dFHX294BgYwR
NYBlOg/F4Q0UaVLQMO7LWtIlJIfxtmqyiF4dNHXRzzVfeGjaB/VW989oCW6hPB2A42PYt3b2gId1
hWPI7nvInsLf8zDHkOavGxNQ/nyR8Ezq1jA7+kro2+tnQQz03+8FWiixK5Clei+5ifTEQNXGH0a9
8+Y0Ln6PigfAELgydInky8Ai6hLxKWizbpk2GrpyvmFgfIj9e42VdhIh1RsleQ3JifyoNshOfVdS
cSOyWKgNuwC24nYHIN54icxmTsbqxE/cJ0IOY+mJ26T2Wc9NYjcgIrzzxYT9684TiQkcLNzPuVCf
/LVD1ak3I3IhEHEvxsRP7LCySAwIoi+0HfIXTNosMoYJsItjAS9wGREtB2ub6e9orBaQl/88CrQw
kg0pTkg+fhbw95GSzEf00hOzcRl5pGfP3dtZSSVQSUAuAshWw0mQvrOtWB+uLx/bp0CLxzVISFjY
g82Bi5s5bG/875YvBvn2KQp+Olr1e65/ugv1TnNecwyIvqed/K0R5ieyGCfnKA3tkNbM4JkSzirs
N27y8v3IwwPcu48yuSWEoeSkPRAIVnGTh6mMRTrc098228Qp5hdLA6W/OOZF8btIb/zR1o6ImDAV
etMy+zG4Z3K2RHa385ju9MbRHoX3B6yZyJDryxbGlMJ7H+t0rBpTN8nBKQGxsaf11zVlCkI6xr01
YtQkfVHGD2HWJA3nqoD598LjMPA7AG/6k99pDlCPbz4f2fMWuMdUdimbhzbce3/EgQx7y32kTy+f
9wgwHdWkIrpY4hU8IVxFl4wPfhkAk0wYgDN4KirlV8rx0r1UpqPELN3Itbd+fFy5VC3u6juT19D7
HUy4x9WNO3+kLzmW7xzv1SCa5r+b/Cscmw71F0frEP3frPA1dWpHV2m6G4Dcs4dsu0lHfhI6ApFO
0Mz3B1dvE3PVAcRNWtivpuyR1MOUc9NV880fcN2V35TRSONFCDCKkpi27nBgy4vCI5iyd/JsD3/6
Z+W2Jp7NX9Da2E8Ae7sQwlMguccWSJdooRYVLQyI3WVW+uqrNDqb8dF01Z06kNxliuzKz3PULclP
Ic+ejuxP8kzlUp1ZTO782HAMKaBLcCsu7BZl7TqHY2ejl0iHjDOGlVvNqVAzOzTQaMuqCr6hpLnA
SdgamullCXOpSrisUrzBG7ukjw45acu3NNqIBELi0y6l1SdqyHMyf1vsfcuQzRoa4xDd80KH+piD
8OdKkn41XNFe2qKEyGRBgNho6EK9th1yLrQ8cR5sWDziYmqzYFGBTH4wt1xyj6wDdUaBO2xS6OqF
9+dxeera8kVR/DdghL5XF0xjlqI81nMI2etj5QUm3syUG0AX5Kcz4d1fniOSaC2bXLTnvzCD7ydj
sFRDEi7C5kLWtYO9x1byw1/S6r5WngIcmmkEnO7ANiQg/uVSm4OTzhRYDvabzea07z/O/WEJLYz0
wAng6jkfMydlPJ7i2qkCBGHh6EaWyvnY4axxWzvV9knzYMSYP763EZmPtRiIM6z3bETnU/LGT7ca
OygM5Qrhz71vSYKCjDIa5EAQIYi0F7xQjT++o1kLdIYVq2Fh+7e79vJz3LxLPNvZSA3dC2Hk3397
WT5klIZXH8+YmOB6Vv+5d4bRsEwZtgjgbwOgOVGgbT2rV1tJe2dnD1yqPdHq6ucNMZg5VZfxrjHe
/rEeFGzBYX6icm7JX6xwYWu5TqJvhNN3+sjrFT/uJN6ZjiQh4mAk5VBWEI5GI6ZXNRQl5HZMVVW+
zDKxf63RHjutX4Q6AkiE7rG/IqLJtk0xFc30atrkPIEboDaCZwe9KfXKxUkEPCSOzv07IHerSLhY
y2pL7WhD0qnzmHV+lZw7G13s/0hNoSeUpUriOBmoovFWaY8btIAvof9diKCmmxGSjr77CzmoeL/y
91ocguBUKt0TcOADiYPouHprJ31zJJsWT/EpQDt9n3DGHr+iyDSrxfkyB7I73CGxgaRoexUbgaxk
FVGxi9rkCLILoTHZrs5vc0fO3fMCHR69rZEHu1Cbz5UDVfRJ64Mc6XTyTpgQEUCuPscRkXSIBby+
QfDfumfFwN03Fm76dkEjJU9/6T51TcvILy6f8Lr77XAuo9aNRbK6N1j187CCiGnaogOSC760Prvg
7xcCxTcFsZPfT1thwM1gHdPKNA1VRrzrkmKLk1mTzyu+ht8Zuty/yHtJlakV/GFagExzuVMGHYbk
9Y+YczEwa0TYgi87M5W6nFOLHIrzJT3frq9HLg2DCkaT58Nf09bFDG/UHkYDmY/qNdVvJ6CpzI2M
yd4Qy7yW6V+xdk1MDIKRYlPDNDLGGMrbaNBUwGAX7IE+mCGaSbIApZ3U0AycMxuHiM1rz4PvrHbz
3yJ0i19eqt7xRFOhw8lQdi5grSKHQTT6cQlAi9uJydGfpMH5uwtcQBY10wQX1Lh8jYRFFxu0+Gjp
9xaK9uekpAlw7J1E/WOM66MweGZvQ9tGUz1AmD+LVZjyMw7rGjBj4cMd9vK9P2P6grSpVOTJ3WwX
PMDEa53OXWKdAYxiPnrP/DBjpDd5qlBvInSn4ONfwIoqzc94OA98v3JcDWqQg8ju9/hX2XTtenGn
ZUVSmBa1wXUyAkNTFcPR5ARBw2ZgaZPL7KZN7ttdxbOsCe3LELUcEiIN2t8Yu0nz3pgJrv2d9MEn
hmUyb8UtjlB+OIDkNKad+EzO67+9KxomiKs+WvdGsWUE8Dz6TIspje/vMH2fYdppJWZpfyID+gto
YIXey2lqwx9Zm6t6zEz2aSKXTTszQwVvw8pzM8Jjsu2A+VCAAo69KlS/D4/wzEoE6hEi23warHAJ
NGX8Yf6W6K2PtPLI0/VTk92mtLaOSp/uwCwuCYiQxwoTwacHDpbdzkVhM6knz3zunGelfTumr9zV
tE1kqVCllMlRTsNZ31x7gpfOXp4p8N/LZe25dzF1FQ2KJrKJJi3aYsiJgFzz0M19alnnSayWxXvr
uyuwT/368HF3XzvQ/DCkZeCeJZJwlyiKwALdHf/tGRzmWTlFMbgruIKV7kAwWS9jrBmbsHukNOi9
GzaaYKAI2Dv3bnpFPQpLbYg7UQqmrsiquRwKCGTgtqnzUCFdRR4vfG8bBLkL2McPASrv0ZWkfZRC
bg3fWBbpcxNUHtY5XGEqg62drvmEXYAoNGJQei0rL2sOu67a52SPAKTS4mEEb+ZWyJB3xP6Ihts4
3hdKlySvvGuc4NCT8gQ6jwqPqVmvr6twb4e75x7CHoqg05/mi27pPXC9iCHn8lLfRaktgyVGhWtQ
lV2jG3pl8CUylG16Rkp9MbrT2m1t3lJOBplMLO3u/6vVgQx4hDCD1Qx+4tat0sOdGpKH7sCbZ/3V
hNe6mA5JXtmci2dSrAPPzqWImwK2l00IyESCQQzy6CQ8SXRKtb+K1keE+jftHyhC2y3hrLU8URBJ
phv895BfyYAdPLEo5tM/gWm8zRKbDiTtza+9w0M5k4Vyhk04Z9UROFiUQdbgKJDno0Nc/V4fpSpS
O9gt6N64TOO6WGT53yZLIl9IjjCHIFwzQsrUdZFkwMFmGnobXpQWt4jKyx8Vb9LfLu9ktfln0D3L
LStdZsm/gwy7B0tpMPLJZ7j/oQLw00uQKnOWSUw6R2RwCZMbUs7VrboF9cmpFnD4GwSCXmEQ+xyA
j2DWQovCPeJzcTYw7U1+jBrDzfV9Hsd8WTckHB+a/x2lKz51p4NIgGkdFc2nXopTn2oDaJ+ASGLM
ieBeCHS56+OLTK0XbOdrkozJETzTaRm2ngCRRnqaYH3rrhqTNiGuKok0bxqA5DF8xs8SEEmG72/o
CJepyn5tDS0i5dzda9uDE3wqUmWPK0G5ph3tFuZNAXHiN+IqU9ZDqMc82T+lAHgfKqzIcV/B41om
RndU5+ZBLE0PVqjx/IlMaToATW1gF0qFb+tDMuJD3UqnCAztyjwDkX0KGfZ98JoF2j1GnVu4kp2c
B6TqygQWKTaCQo/yo4eY8Z7XVvwtru3mnbPkivyaMLFNHtwiw4SI4cLa21gCV+aZ/zLnlnLaexLI
/HX/1OVFm5mwjd76eZUHcFaBviLSWc0XYqAIO+YSE5Ws1ph5JHYEbLdeBnalEPOrenZa6CGGC2rl
+yFT9ycFNIHYirId3oDEFNEagldMGPZuf4SnF4u914YYW0XX1pz/Il5/1AUBK72n2K8eN7olxIcA
h4aPsHidjexaufEtcH2qAX+EQ3EfnHv4y13VQIypWlvZOxQ0HdWN5CP6TxaZYhsVWFIKlwW7KL0r
OltSwM1tlN4ZrWcAsVWTlzk3f+gYUHd2B0fQV8/W+qPYJP9P7fjLDeje/XMYvgCSOpMu7ZBWoMqW
NoAmcSMmbileP/5n7++XmMa/y4ypIEgAqhJlPLGOedLS/mH+z85pp56GEECirYljNEuoD/OwVT3U
L4f6iqkF5G2B3r76Qs73WOSg1nuYeFs2qsD4eV1Ty5gqzEt1So/Jy1G6qdnLfOPcCGF7gRRaA2yh
SKGzPzwAgwGDHjM9qbcPsEGQ261hMwTkkkmdjODBEFXjOHNdBbFneGJUXhFuoj2MdY+Q6Y/m6if7
rN/DfZ9vPjxSaexlgyXdCS5jwy25vjIOYWa4hHAPc1zWu97q5ibl+KY0R+Msni0c5k34e/YKTPnM
EyrkSpGOcVGEThzhB0KVEziUJv/ZqmB6hWaWpMFW20qgVcr/wMTGo95NDeS0T6FX1g61oTTO2K2P
TlLnvlGNP68VObAHEKsBR892R66RMQVrOJ4m4l0DBZOR4iuoOU1KPhuzvwnTJBqdliWNgZ7ZtK0f
7LdV2qdM7ZGwQKAyAr8+tSi+1EoBzrE+mWm45UQWn6f7AKrjw1B9unOX9nuolxmXMXOXoTmQ6WA4
9/FuRloUwecv47sZ03J1LOs1bcHPZwhdgBVrhp5vDsl8A6fhqr5A62jxqItDZUOANOgSXb1TkQD6
QhqzO4yQ8kwOwryFhs4t9Eno9IarNMWWD04Si+PRv4rH2cudUgqJ/lATf0Mo5mhkVNxkeEbBTwtd
0ZtiwDYn+VdAZtJTAFTpmyODNg1fZMskzCyXamXELFI0YPoWVkgr1Qkkz4NQIwjbq54GD4Cjq4hu
e44BAAo+XSpYtzhViHpYRj0NflKg6n6ovNwk9/ZC690+xVodU2hPd48xsda3n0RH/8uClpZXUmth
3SRKVXRb+s1JUEllRRY+HreCZDBxionKeF8wGfkswOMZ2o3GAQFzQ+EBidj91NW9O5OzF/JO+fVj
W+CZ7So0NN/V56UK3PoHWQUJzA0d32J35qfs0Ypt+TiGU/00LuLU9ztHqrJgjYaJwNeYapHhpzve
z0Aw9PRzC1Vyc39qWQC+uY9ZXzSkmQzmxdKQ5AXYRrDlBn5IqlFF47ajsThjNuE8bKpFrBKCTwgo
TYYFZIc4DpyE6LNy02tRSc8thHJKKpfAVh9keTVVCFVY4g/lmyf5LDJqq+uq2H8vfTysBw5xW7Pn
FHUWfpnebTjfsOvtuUgIqNteDkjpTyV8XShUCLbtLHOg3b0v7anQjLKkdKz2xfLj4zYKOTOJptnK
7XGQt5i67zN/jc3AUENBmsKxm40kPvI2erOCWg/4wQmeaG5P/XweqJIS2YROJgEJO9fQzuVZWD+Q
G0S4KCUwxZtqTMIkJxsxzF5ngaB8Ncfj2mWCbGwUNr6JE7177JvIf1/cXCfIpqKhY0ijmaj3Mwqp
bxrobN9pfsRflUCnNtEhCENLTI+Ew7zgNSfqYLIz5L5zLp3NpXw3oOabF6e30w1sam7k2ox0zjNE
M/JlE3ADTvQiSRQNsPfky60kAosG6je3pKN/XbsHESjH2SLy5pZxopLT5sM9SB4J+x/Ml+A4xoVc
gLE/7qdvU33Wg2YivZsr4zihLngcez7aWDmdzpn6hMmk5evlM4e5AiKm7RWobgj860hc4Z8bzW3j
5ywaEbLlgCrFICx9ydIT688RsxxgOCFZjMxNeg0ItOax7X6pRu7SRtxeg1+U6M2X8rV7ZHPPcGCo
C026LVP7cmMhmJhchng1+KSHNmf8JskZSC8vyTXmQFvvqTLtOzaQksYg9QwzQ+APca03kO8+zzaY
+rpGvbM2BdlsIIafpNkdCr1EiOgqKhwW0HDuZpDbs6Xpy4OQGlGL80GeNlgLPM01FOzT5exkDh4b
nEYP1gWk2h6s8JujVMrfHZxeOwgZvn592MVBTplODYrXU9gBt3TsI5V9Ma2mhnt01t2S0nTJkWdS
Tfy9NjJMMseOP5nsQlm4iBbFCID4xi8sC9PeSJvWdmVYphN9T0DWZkcRivg8fgPtqfpXLHhsI77f
qc+bO5Bz2AnkDHQ1TkQn5AdBilgNmynLq/EJnVTyaob6tRVY0S8tmJN1htFzOo57W+5i7FQIwYSd
R6BzlkiUsQKdXAGyYNjWkbUROhjOiz4HBZyvLUXJrnhojqvfRrdzWVDcs6iAjNNS7SHfTpOuQrv+
gEpnXy4B02UzXoeK+Fr6Khiarm/YM1g4N/+Mmt61Da2jKAp1r5t6yjw9iqYIB7BLmS86bC94+St5
qvRdsXR42nYa9F6ugpowEHqK9V8COKAnaEdzcxvL/1qocLnRobjRZ/+7OFHKlTVL3NHdFUUn90YW
HR8gKU9rd1LyhENKLSWM96+2NBH83BHqzpmpnIDmNzx9DHNhfB5CjeYvnEweFuIKhdRxUawmFo43
GCaUo4tTddvNiR/iPvF3Rd9UM9h0HszOMZW0HPcA2J9z+U0XurG+KjPj9jLEKHz8vfMKQZ0uJkQ6
yni4XkvqfENNa4m3iLw3Xsa6qO6AxKLfJfeR1H7no06jA8Aea3TRQlu/BZv3KC4KwCwENzDcHnWr
9og5n+FYYV/gxfNPlJUET5noylVwz1wxvccCfAiFeGnfrtG7rBb/n1vXgR8bm2pT8FU8ftXbJBiW
7fkYoo+Gn1x4Bp4DptCilr0kdoThlb/y2YkO/ki+mjYMphJy900AbMlT6cqhzmxnc0UyiPSt5ENT
byZkRTGuY+ul8eAbY/YtKo75kMLw5Jrszi+Mynb4GLfs2O5hjQlJvBwV8uUF/l2ijgw+HIXc9/Jw
MHE46y+Cwscqr25YGQflxF3Pf38g2IPMIxdR+WtsDWsDCfx3j520IJjOb8vi/0DvoY8gyFSaMKia
Pl5dzyrFpV5sVhkQP7M3hPolTIKrEAmmgb+PSA4AzJ2a70gh3wRQvPwC4J/fgM8C3SMGON6bxPaI
PZqWFxuhSTv4WNWn+EYpxNvS3o/m5RhMgyjQjjOUrc44EuHiGOmW/Usd5cxlKi5+KxJjvVokTtvu
NQ9kMSwdq6VBx2zK4cjk5hr1FUwQVxs57TypPIPkyr2CqrEV2kW5DhpImEFF/WKJlDzASLMUEnbq
iMTgjTIWDnQShFfgqd3xI0f3YpX1hrRcUO9nERc+8TxLUmpJVZKYVck4r+b0eKQmXOEHTxsPCHH8
PtKqIs341FvO30NKqWYV6tb6t2IgtzOi04S/Z3VUoh+ryf9eJOYOBEJZxnX7finrdlJou9JKC0qn
ZoFDgWhhlAYVCeSffa4gIqySfgFKXfcZlbM/YalIlbKtxqGB5mWBaIV1i52d3C2nKNLvoqel3K9n
Cz9pH3x6lM6INIOA1IJjuqDrG8Qk80EUgF52iSr66FgWVnjZJVyz3nEvGok9yghEu4i5B/EySa9K
hoXx2wTD6kF/cozgKI6Wo58eeHe4HBLNeGFE2lFckGar64/bH3eHND/JrSJWcbutro2OfLqfxF7C
iPvL1BweuvPei770IOl08Yjhk3//FxiDX8ER/6PSKVuWX+8tU5zMifEQGZIofzjwuqrr8lb/Uqlz
UO5sNjzGOP5px9DqTW/8I9kJEHDcEWilPYgAWpw9uFSWd3psOE3pKs8SRx0KhwYvyQ56LE2vrBWl
6BnmVS6NOEKCZqQlpPhPm5tZOVizhgbqv9HSlsagGzHf+Hc34pifP5QC6bbMRbPfRLMRUHfzrnxX
bs1pAGF5/CzXU3WE7ekpgiS9OO9nX+roRTYtPp7efvbGTkp4nhWboBmshNUO3t3CEVTV7ktAvqIj
KAQy3MyVkQy1idGJOvXJGE1/PXUmNNl0C/rUXVAT0AD4fsBtnzD2BLCDN7OIrweOl4vud5RqrPup
gR5rI2kaCJYTv9KMHxBEAUYsqDyIIv6nrfrS3AhhmuOvRUWq9FCnD33h02Nig71TtMr4J89fUdL9
b20lKEg2N9fnl84THNEwyD5IDihW8xZ59aSwlLfy7TdGY9LERT9ENwV0qm87GBR0kgxEMYXdInyt
Z4J5ePVgxopqtTsHtBkKzKa2eoSxUQEW6yTRtPHmxTPgZdueEhfRZKlTz/7uP+R28bWcRmXsBZ5p
ondwPF0LwCRi3jzWjruHyg8IDd062HJcSarrCDakTAAzKdo5cR4lUuu1JcxD4EGJWrognAaGetYz
PAwJqhtEQxKJxbVRY0MxIP4XPscQymeOY4/ZTRuLP5vVDoNmq+vdXXsTDdhTevdnvsTTqdLuW/Ys
0S5EYQehzBAvcy4uJu5nIW2QWGORnG6uucMGAq+XEr/JDQI605Ef0B7tKbvZ93UQ6ojS60phLrVE
TOM0qBSacVaFCIh9M0Yil1Cng4/r+FjnjQCgVnTRG/p2RJupOLqUF/6Co9dSgVBPkXZXvL1AfgVl
1wwkxm+k4mi+n3qidV+3jBZpEHKlcTe0Dmc1LxColARqSvhS8h4uScsywIwALFwGv6FcLRy+OCss
nDfXejTm8QH3+i+tETrJ/UTJn6267rqDUsxY92c0z3nx7ba5wUvv4qA/2OuenBMNgVvOCzbPrqPe
05wjNIUMbLc9hpIqy3ZtHwtAax65DC8XIFX5NYFrkySTbcPUR2Cm6Tl9BT6n0+VnNetvYS6tYvlb
TbrX9TWoAsRzjO3DP4tUHJXB5nBmpihcRmhPeGszhzdMeoZtyhYUDUz14z19RJJDhJpZ4j9Eib1G
cxHmG5rBlVJMt4EbZ7ThFzsFoINw8w6+c9QyiPH2EBBc82rxNitFyIzHrWNOB3TwLOeX0Tk+syVh
YwpRPnE36tg3HethZkAynigTVXSxeSiq/ws0LR0vwu+3wlRSnQxjwrOe8ZLv9aCSMxHEzhihxTj8
pcHHLDWsN/PL+2QlDQqfJkLga5Anh6VLxhomsfu9dcDmNiyAbOVYdDtCAuDC0i6K9rmvw9vOWdKx
RfjV5kZG75hBCaWBnHWdholsKV3RgA3Q3WUGE+5nvKZP0yK3bvCgJke/UxKj+/zAX/JbGLHXXpMw
UF2TvCuPvB3x/I1/1SLUcB0zT3ro9WD2BRsxtbsZfmM99cHOL+NuERbeLwfAGUlOlRm0hpN2t3Od
A6Fq69rVaEmmyRNfJ6ULAsxFyl+ntSDg6CeJZQohJjDC6OXbsNOaBnFB3t9yj98Gq7/j7AqeC6RJ
c87GjoCrDTxYbxkfKcDf5uca6J3kFwJc5VsW6Eq6SO0onXDjkNKjMmUa0SPWFG1DzT8PDrIe32zB
K0W8eoUFfGY+oqU9BCH2/5mjXb5wJMhT7GhmUW2sU3RoZvVwAaBq541uvJ4j0vr6sX3Jisq2L4Eh
sIUnse5TLM7Sw0xm/KM5lLFiaGB6e2lQeCYI9ll0spJtoGCyLpmvwPnCSBpzPrz0q8l/xGtaFAtY
zCM+S2KJDkOJbrtHOn+7yanAqvzY1s8cCE5Xcz/HVbILIzec3fC7BVrRSt86wksNfsrTDpDSJcs6
ScW8Kc0Rgyat1RNjs89K78CyhjpoArtzfJr41RWxWnnwdfyF4vh3AeT3v/BUDBCZr/8kP6kW6B5+
rr/OMmclxc4pVpBO602IbUapoEWMEbliJ+P8Y7BM82Jt+RSzynDuY3xQtsKByIJzkUuXUE24bEwH
ZNc7PEJ+VQWbJN79kXmJd5fP3doZmyX5BVIFcGBrW87DCApfquI02Uk4q/cb5nN89uchtNuCKT5q
37TGNeFgtztHHf4EFbX8RUKaCkiIWI2qVrW7g94c/dbXWTcGKILaISCQge6RjLn9f0Fu96lDy34C
PH5lslN66KRA4EgrtkFs7rb+eKMgDsUP3a/nr1lVf9Ux9Xo0O/94XE/MeSSF0AD2Juua+3CC5yeh
76L4E1OGzR4dBmNxjvwXV4Rzf3CAxkxo+eews+phm8CcWW/8NAaOTstMw4Knqn4lQsi7++YYbtGl
Hxi2luhojS8R9zGA72ip1hZ/VT5H5U7K5dmSqXP3ZpExkipFxxWBHxvjgvj4hRn9eAkCzOScEUSK
oxPYfrGq/IOz4YFcOrVNPE5+zzsMgLy1GzhoOttyanxW3EpY4cx+0RofIZ6hhxY9jyIThkLBcEzV
HEWlTXKN6xK447VDfAPfJkfcFSUn4moQTHGxstD1uzxI2E0DCZwq7SSWR2cpHEpWcKivqPVVRiqP
y57ft/w8MJvKC1rqhb189gGhiQJNbT0r08W1tyhHXFaP0yupxVN4NcPoD2vfdJ/ecQ/PCLi5HbZ4
PGuVqAByviBQPjJFXJj0jCjQpVAtphT6lJNByGwsgpEE6P93ytaKDktKnrKn73Q02DD/fP2e4SS6
Mgu3DEFMDFzc4vWuj39bCfBXIyUPwP+RFPO55buYX+Jiq5nNDOayXd0WxT7KshlL32FK91RA0MJq
kjEecUWEE3VAvo8Oz4/td+TggiqHRvyABE4iy6knXr26S1tKqfATc0uC7+JuxgsGVVXDlNdjZGcG
B+eKwO4swzvTVAqYajMtWbsXSs3/sRm6d0KyZeU0y4ntAeOfJJEuCg+/UqTCyQPbXP2t2kVdKbbM
QKZOxt6Lf2Ffjx/6YM+GLuxsgde+3LC2oBnO6grdCi56pZ4XbR5aBi8SDNhrnvnG+J33LJCrTVbE
H8mcuVp4yTp6HY7GyV9oXWe0ToKlsB7e7vFA3Op2bqz4XVnoh3jVwSaPKzl/taW3A1QpDP3N9yAq
NcyIOeh62XLzrl5hWdR+bbFeXSaopTSTh0FcEvbYrxJ21LMv5RETWMsbMkpr1EMPmVYCQJjy99UF
ehYvNMM9wTwyoDSwfeb7mNIOVt2eLvt//IUoyy83SESOitOHWtBn6g8yjBJOsY01tkl6zKBKrSJT
ylSH6dX2SAjrHaciAOAAc1Ej70g6VRH49+6ZXylJ7UOgpyNNFIBrOMjPlezt5AR8FV/S1aydEkz9
a6r8JNdR2S/2slBJ62BdjgqrWvBAYsokYJ7i14VJxXoCUp7oAS9+59DlhpWhreoxC2zKuFN9TXDz
CM/X+qmjrNe4E/uZR56QALMIGbNixIxZBnnAhll/8WfC4fp2mDSQsZX+BkrhOV9NGHk25dh84cvT
feb3l/Y0KjIByEaKZzDWIklQkdVIgrqp4hIwd6uNs90G5gmxeI96H2i2BsjTVywHV9XfBHHg1Ea8
6Zon5QxrLUn2CQwncQ5+oqvq6FdgDp5yzHoO0K5Too9YZDDfA7Nors6cEAnJKqgtXHPZHU039aDi
Rn7Gee4HXIAyfJt5iQD7l8hjW11c8XvLkbZ4cPZ1MFk9sGO0hiKx0PJfYHmgVuSyx5Ws0CxcLhix
Vj16j3+SVsqqZZhQgekWfj4pzgjDTp46KJbyKFmSqj+QJjajEcpsQC8FLDi9hWxf2vKFL3ZxbrJq
/7c0gly2cH5IqlzQvjt+MujpyNjteleKeZpicuUtNq5nIRh6Uf2E60ydVEf1rPyMkUFw/wfgFZXA
jihCVQP+mIrIIfv7ZrHM0wPf83+6p/tvNUllc9w6hSaMccbocW2eWSX6RVvTz/QiSGf0cPVbSSk+
AKuOWLZDlgb5j3p7SMzoKeDeThLmzEQdjrK7JcE4SfG8sa0OkBXcA9g11Ko+UbSryILLYqY639Zw
/H1Zjbeh+/p2em/giFromeSwo+ATP2buuPh+nKyUyWBt1LeTCMohFmRZ9ix9WT31bI07Ip2tUWWK
K46KuBiHXBY/Us9iUdg5BEzS5F/uQFFJ9gtzKER94j/ASOoB42BARU2qSsqmRxlaYIZ3AgNV5Iqd
RAuh+ztg+QioUWvsyAidwhvJiJtIKynLHz2Rpf/DFTbUPdmWnZqgneQGJmR0ldltaiL94DwZ9KLM
35anNkKQm92ggTtPBH3NM6gCaDnmwdhEL1ve97zPmkoy1121shhiKLgvylu234fI/WZa+5SCBn3o
FxQQN0z514yPA1QgiwtWi2X+1u06sJ+OMrGy6BExUzYF59oeYhHp2FESDE31V6yxIRbwXHxSB3M5
pQdpemJii4DSiAPAnOmZ+3o0X7EfCIH0G4HHwOz5JGN0PpFB8VLAAbDcZ8bha687twpN2xMmrLDs
RD3pArBhxEfJlkiq6Nui6cy4UsR89+DzmccHy7ju0G7WxYJx0WylrvcIYJj45GAYB1ZbBm5i5owG
/HIg4i8MvVNQg7gO7UORdQDbLJ8qjskjKzMoFMrsWknN4mrGeYXoQBL72TmzyiNieWbSvtvlRTxV
3pCp7Dqu42vJGzQsIiTCnZjTxihsD6HhovI1O9WlsENl9LyJPvkU5woBzv4EUy6tGNUoZ7PYHbTO
Fzy3/1VFIm683O4I4L+QXv8Eq4djptVvqZwmt5xfAkY/OxStVffTnT+Fqe55M9uY2gsvHc3kXl9H
kmW1JeeB1clsvkvV1fZkLknhNMYAT2gEdFAXYgDIeztC2jGp4IWNiVhDpq1AXBASrZF+HCghcmOT
N/uph2WwhtAA0G6qlZUXpE8OcyMQTRAigUH02n7bsLR8v/DkxSPFl0prDDTqeyW1hNrcGbIvO1NU
+zhL9l2Tw7SXfo6++ok1u1ESrImpFVC9iGs2lXkHb8112VLCUQZxhdfd5dc1eBKNH3MsoRgGo5oo
LcH493lCyup4QH2FHTTOaxbLgk8vpKvXbuRihEfNwsQXUjF93/eS3oq54DZW8M1QBYtjfm9Q5ZVL
ysbptw8cXElpJ+NdU/Zi44KH2O4aEZX2dcUTGAcyxYg/LI7WmcoldAFzjrBvBe01L4aIHRVYUI2f
78uiH1RHUYN3NxVz2EhBdx4IysjmhMUlE60W8Go/vaNoezqzuA8zLXxSz3cEwx7BO4J9P3qvfBxE
2VZJVhw3O6JJvTJhR19t7OQSBi9ExS0h6gB96obFPpv0A9dNLGv0RMkTnXP36hEkgohqpJggBgKV
clnRSgUuzN2hJ6Z4nNFgqj76QPwKurx+/zq/9z/lUyd2LjOuSovxgarkfpwZPMIPU7/mJp2r00GL
oW9WgK9QrVmXtgOEO46W0zw9S85Hh/uthYX2g7zd9I81KUBa/3BqI+Q+5upqzRVZCLuNR+Fvbncx
0jgUaPshz1ik3GeYuTOeYZBz2+CoHGqSuLXEwu4wXvhO12q1PZd0Fm645zkv/AIDDwQ8BO3vLYVR
HUts2vLuwJETJcixKhUI+kGEnEeFGpsbHcwQjeML0vNkv5lqDCyj86qfvo2/bnLgPv4VZxXKcfX+
AE510Nu83W0wZFGL2PQbI05ejiBUak0HdTP82FWCKjYLBnjPUAJplleU49ZrWCXaGhLspm+JtfZr
3NgB3ifaSvnRL1xvY4LTUX0GDXWZLqhQXvRHVS/lSIUt8cKOsY3bbJN42K/Z2IofYH2Z1pOh0nr/
gZRdp21Vzczi/WE0PVPs04jnj98bzb8tp3N1afUi10gdMaO0tKBrPSZgaTT9tYNZxW9G62qwlbcS
YqfoUbyjKSkWXXFMsBOunGaM6U2J+ht5kFkO5CVAnlDdMZpmWHZ8ytUWuvzM5ly64JYG93AEnRT1
DTeMWnoPYmWvwF8nyvFkrfVwBokHkHgF8uTOlbEX78di3zHh8nlkCa5PuQ6GMciM7SeecQ5/1PX3
DyWTNj1ZDUDCRjLuloERnka+AZTAFQUXTHfyHh/7sBJa7enOA9dBlIxmHxhPxegXKRGxIPP8SW5P
m8xO7ILN8kn7aa6FMroAIASRtDGheqmYbhhxViN5/jk8dQj7K4Jx/jjeGCLi5s6QmIdYYHEACHDK
I0a/ad9w+djA4ND9kr5WhHhnHzXcQv8sxQOX5AVtMmCkBbHskKAR1TGMmEmOSbr0Idd2XgsQg7/M
txPOONkAgWl+88uLQ/ekj1W/8BC/qTWU5ST3c8YkY8kSMBYTc+/hD4+rWS8+P4FcEATBZM/e4Stq
fCbTZaCeaQ9MGrxJZltCoTkjEiT6BgT/yutrH+lrY8gtuB/VGWDJC8cUqYfufiObfRJ7zvZzqsF4
8Q0j2XcZGGs+n09GMa/8KaMAwOIq5q6D9IGbk+ohxv3daMuAU9iaiWDlX2ehRYDGW2f9VmNARazB
KFWNQsPUKfENgwXXX8VfNwBbvgECQxxXPPsM5nTQ+dD/yohLZvS3Mh/9qUR7zCGMDbVHxP+/MXxl
1Wc+2Zky6sgCphgfbjYlbt10fofj0XFs/A7meddKs00rQ+IcXznPRh1u2CLwKmNxTshYBUPmD51T
GBcX4XiVU3yIrEWQlLGcUR8rYno7j+RyLCkqQ2uM7whOikfP+3BNyx52VOeh5GiVe4jAuEH5X/TK
KooBr4rh0Jt6DIUpslkdpJQpjLwiFjTfTrfxrgKRARnJwponBIJ+9+eeEkWpi2F7XlaO0jG1BsVB
9j3G6sshQuYmnhy19aD4Fna90LeddzCpP6wF/IUuuWweKNG2m6zdsG5pTFOk5fnD+4oDcn3N/1VD
o2BDRmPg20DMGo25P+Ia0uRFGEMRB/gJCx+gll8kEeGUxXVRV8zGGw8Oyr6fa4F1IQYcW7HEifRC
uYlFH8yu82VJBOKKN6BKthE6aVy0jAb/qX/sva0n4GaNnzqwgb6TWG7eVKM1q5XN7D+cuNGUNJOf
hWUd88LxVmbGbFGfRgRSStCcjtuquhc+NjDblDdifd0Gicj4qVrlX4ckga/9bnfG6Lrbuuvy19hk
9dNUsx1VD/eIhP8A9MwDB55HruOCzufB9r81N7IhNgIOXpjdJGsg6g9tFe//11I2BxEBxGnBPecU
mS6JtYvXiWZ96WitZAyBGQS17HzL7uO/sQxbQeOloUsg7ug0C301F0aRO4UyvH14+PCjzB8OLqis
rM/LrDVPOU+pfGHlSin0wCZaRDw6nwyppjL3jXSQ2s1RpCnae4yChBMhbHWdSnW6vKpLWGbu+61T
utVm5M5D4Xe2OQT2yihj/ZIX4ab763Gto73h9PXXE39WDXuOIEUsVITh6TtnWxs6HzOVT2NMftpW
MHH7r6OF5pPB5CH+DkXg3za16mVVlfGB04hI4tpTRxqLz1NbW5b7Uw8C75z39wekQ1I/qURrMsAc
Vu371TDO7ZZ3Qbsm7zhDrRBNwgJK92rC07ccENEeljsrLrlT0rBXM4DzSUzCSXHpD33QFq5YLm7v
z9iSGGwkuhmPErouPsXJ3SjTkHUTjqKsIcXn2IDmieUrjNNJ4QO7UdgFaE+ySJSWj1Jj4CAOM9/O
EF6zaHantcVfPfr9a3/7Z+Fl8lV8M4BlIw/5+VDVykr1oUFKS1riyGqfV31+JiF370/Q+fsDWHai
eeifPqzfccdnXT94yeaw5Abzx/EMRE9DWr1r4b1rGK3Lpu0UOsXviyIRTXunZkN7PJs1dMK0nBxf
OD7tSyo2ynhHBERhueejNljXjNGmTq8xb1IGg0JHbyZUKe1lW2h1KMZkOQNjQBkY1k1SXkyCWbHm
aYiGMby80fZbbY6h1aFO3xjhb00AukUl5Z/qpfRa6GYkp7YJIuXaanRYtkH8L3MDSle8Mlk/yLFl
EaSwYfz5CZcOC8YCNFlcR3ihXdjQ3B4fgYR8MM9Jr4QkmeJ09wWl3AR8OMxpbVVjUkBT/11VQc5X
biVxGnjGPwQlVDVgDR+qrtQ67YS5J0+eYehaqRlMOi+MmWhoAROpQvCzFlmAp6m6raCih/Pq0e9U
qDrrTIbCko03zYTyjO/nEU1Qjod3IX0vA/gMQtlmAe+3zsTCeWcC6pQA/m9DaByBx8qP5jHmsj7S
BKEgWqB6cV0qvg16o20QWr1W7bZRjd0jhY9u+K8E825n3z3W49QTB7kqzhABUlH2Il7QiBhycDoV
cUb+MgJxTQRuxz4f911OnxpWO2kcCQUiozshNDpOqc3wKz7azcaQHHyjDqT8VAWn6mQExKBKgPxe
1/yoFaE69dQx7+3st3aLfulgVfulpjZzbJvtKAzbxgKa2qhDVcNDeCHfy1QxPP9WfX7xIHHXyH0y
KdcgKji9+H+YiGqbYngGuSlOzoKssonAt6IQtT1P0hAqcXMKwzy0MnL7ej0Ksi4d+/S3v8Nnbu3F
y82JRK6cefIeX0xNnD/UKfG5dOc+C32lwIID97wqhldVIYhMzTiWWCm2xbUeJf8Pku1HAY5ti8Uw
cqmoCAxRnHBn7bsbQHczyspyUlRCEjoW/cbmyPVupbv83T0fgGfnzigcHE/8ClG75hLhUfsJoZO6
R9eAoo41+xwxSp6Z7z97+IfLXZu06Zir8VptT7P/QfSDF1+8SAm3ic7kHyggRbTTkuhPt2ZtS4HX
YptCupIcADcM0OQQkgiiMo0z8NJv7fdNthrnceM/iCDvbvMQni7n/+YgeRqd4XAEDDjVIFlx4Dap
mAVQSEF8HqhPusm5NwJVd58uHcuivGg8RYjZt5ISaJz3MAcxkaRA11ZnuUupbAFJPSu71cYpA12y
0L2jCHqF1ZDiVQSFjeRL1Gweh6OjIDp/zWKEN2w2rTkQXU0iVQ9G/ieuUPtWbSQfRP0f5FBskJ03
Vpm66zjQbd2jeXd8TmoAOi9/cgTWSsjGyt93pdVVzcMdfpX2nBITQ/VngRW31F7g9LXsVfw/0oFh
Xq9jopSdstKHPfLdYC9thrn53Y6VPbLXVitd7I3XvjMNFlCKo1rnyQaNqcyv78vJrb2T+vxvg7EX
fNh/S0sYI6WZoT/D8RdFSPWRowwezfKCNVC2UTgXKn65vqTlUpUhTDPP/IU9OlDudYY6IfcjFb2m
1a4G5LNuq3jbrLu9zyt2+Zzddi3Ny1A8Bq7m3Ql8BD0zhBnCCDDML+s8nioBGc+yOudT60hyUwCn
CDqXbe6qo7qjer3oZYz7GpUWUZzjrwrFe0Wo7cSAwkeXSipv00/odsIDuZsx8oyVDbKZqG1sR4Vl
Uh352XrR7PXHPcteU5DLngL+jHD6+3tOaj6RjQnzVJZkddN4DYFf+sQ6kjaLIcqZoj+0Nd5LZDXc
+Vre/i5xeTQwTQ5o2CxYTQeNXdCdMzy5iJ9+Rx4ncM/wcGpOhwA2OVctcOjI6fg6AZrnbBDuMQx4
bTgxYd340i97Jk5RoZxYe1E+Viqy/oxaMCXKKOqlcc9ofxIObRv6cNNu37UYWRf9wEwztrcefM3e
viTo3keAo0HZhJygy4yzGVnwNaZOk1fjhvfdwxURyHQCLHE1gLCSfm+gPHR9IYtqX8VxcgNRIRTT
pq8Dd5AI/sgWqk2+C3Ei7Xj8xgBS4DPrnygYEBNE4bXnqW/haKn/IsiGimdF/Zyt2ctq8FBW79tl
wtMiSvZ3p4v5B+wfxmwN0BFYDornrTzPQasdzyhrTDfdiZsFxITWJmRGTbEZCsNosy8EkC2H/2Et
oNIKK9sEaEObK7HRA4p+A+TWMB3zyDQ8rNLIXReCQX3hQLWd8CNc7Q5F9fdf7KrcVszNN13Uiq04
IkGLjFD7xSJBhKpLHD3Qn020DMUPiMLeQ4lUpqWJ16/GmRtGN9gWRPG099jLumxybzTb7h7KkULv
wh2odZDbrpgyiNfnN2A2jeD5tBwMFSZc1t1mUVzmYcfCIXCBeiWWpXVBMyh5UKT/KTWkfjf1FKOz
Ul+MDebdsxKmLcUX5rrvi0+n8XCPxrT+JBqZtHB/8rB+JhHbRkZZVEkz8mzLTEgo6zlhJ8+eru5K
pySrav/Wkk3X3z61/q4gyNpWBUIAVrpoukCZ63IgWRf4YzQXoUKVCfxQikltc4MqYTAKiuVQUvXe
oU6rkbvB0THMcCFDJgW3Z+K1WitEgJjbSSLo5s99HuHX0hbmquaDM77oaMY73dC9Sf8mzErfGdZV
ZDQXCSwUG3KGmEbxDdfOjp1WAEiS9IjYylJZ4de0TRwA62/ySojF/W6JaPLz5HxUaAgoiGKi/L+B
rpHkmwarLCeCSbSR66i/S4ZDgRkkarq52/Gj9DAmOFMlNOtoOkKtcgASwd1ztQfsT5Clo56eSG3J
Lg3eplnhvVZ3beiwbrXt7JN0M82lwhU/P8D1QqdZ3p6r4eldLFIKElRIWznNFlAmoj4qdPmzajLJ
G1cqINGCc8CaJK/90NXQ1bhjYgI+z1d1o63RmUbvf/PJSkJ5q0hiayJi4X9s4Q0X3PAdUCViIaNe
5ISWKzFB2CCExzqNTaQ9E576z7SE1lrv00ZQM6lcCdpYLuipA6eagPf7BYZ4ZrG03OpTGmObmH8K
8kuJJVzZbIDzG0if05jlVZkX+QaILvtdtMem8EMy+vX+CX+cVkrzJAlONgA+TEbz9MtN4bsiMlN+
xjayRgQwlmiAMB5GhTWGwxauNhLGbmii9hipZ3DUFSB1wUUt0yuMXxeOp8EsU2CAQnKG28Bb9Seh
xes9LkeYyjJPAKZCDjO82uV4ujsPZP/OxM8p6+wpebNvyrHuvtfel/RmEcng/KRjWDnyAliDI9vz
K0usL/60yNEAYIVwoidaT889gJ1Wqg0RQr3jUY/wlSDbKqY8y4r1nXHlHzwkKb/ZknCFKdxMs07i
Vfmxl4s5X604TJMqGr5FAR8BfnbIdWG67ZCKeZJkJCnbk9U3DRPmGTRVEP+OVMAGR0JE+OIESoHV
GSiel71UZFbMAlksyOhKz/5Ax6+IidCm3JPB3g+aUwiTdtAKTV/PooeLBZYzpuJpZJ+r4zKX2II9
GMSdijS2Ja2tQ+JgEj4qeb6SrUwzkH/b2iHJAm2nANKr2y90KsGBOFbxd99AnmzCH1ooxUW5y7PC
PRhLrh+xOPD4ShBZ0FtltjXhDa8w/+DJ6V+G8tltO9akKetM+KjwQpKLATuhLa0y/Ln6iw286G7R
cyZmmXk8obwlbHT7nGzp2uQbLos1G8/h5RKjWF69P8AAVLcOwjPoFWzwHWlXB7rrQ6laRwiL3la7
UbDaULXl1aW4w/Wz/uw9A5tamdHwAGVxrvRJ2w1RLO/oEjGq7A1/aSRxzWkY7MIzgow9OCsBvWXM
1trPT/xNQ5vIAek8G9F6bkVvGKJcj6SnAuHCsp8vTCHeL7AXoai2lRagJJwUZWTz1rbeRJ6NFQnr
FNYU4OZuICOuipp2v1hCFQ82x7gVoqYQCdQcwAI/YEUhr/lJoldMZWYXvSrhD6jCrEl6qJ48tvuF
f/56yt/hBlXjFpZ8P1fONBaUxrktILdqTx9DAEakLnHIDRVLcPVh607pcpDg8zMhDqOmcTb7w9Oe
udkbNe6K7QxomxrJOFB9By4f6PMKm8wyH2/A5fL8SdjxCIis+k4e/8HLLAaql2f18Pxu/tBiZTZj
RM66WBTwXehlyCqCMutD29HjYJUT/p3+W8327dBAS4IxIt12VjW7S3WP87I1qU6ewaMRZnMarb9t
DPMVgv8Nuzz+YBNHjY5edr8e4zLN+h3OK32+RA24OvqAQek0tY2BNrxkl92HJp9krwWwCbyi7j87
umyIcgotZjPivZz34/BlAOvf4vJLoObnjCzAo4A9FJqDwb8HNSz8FKsghKr9DYj7CNAuXJf6ivuc
dwMvK0V39zzuN4SsSW9aewHx/M7oEhYAp/mQWo4SapPmCxClZIUrHmkdUxYs4taPXTkXf2JV0cL6
Vr1cy1YPrS6VBnxP9yvlAwO8P9mkdkpbx3jcFKZiX0yRjriOQChvx/ek5Ha/xcvLbr9W6VO22IHP
k5FPLI9wUvitMX71xye3EPjCHnQn6lNzPI+5oSCX35a/VY45F7Ne1go/jyAc54QGbyQXoRMAxkqe
8KmdPkn4Ousy3y/YOhBBt5FZmf+JIXw9pauNqQBKchFjsbDlG6nwGYyRZ4br5LkwBCgCZVdSfycd
LZnL0ZURmewyyKUnTCPC1R83ETiVQInaCyWZwB/ecUpWsVHbezQCovkvmtxZqlLzE2JzGrfHPzxR
uaFToyLW+mXYg7zrqT+39m2OI+clM1msUkmQKzGnhR95miJY1JrZLkPA4rvujsW6fQC15tYmz5s4
kmI+1d9XwikqXM8bryKgnW4i7+arAwDbTzhivg2eQaR3vbzHk8bMWZpm9fIjoGtM7hBedzuKqghv
eGea/7UrFgZtzxCcQSON9qQQ93P0SCLy3H5SywDbxrL70edmFDXq1jQS3JpsZexAQZar5tTKVJAc
TdbvEe5BJzTSjIo2taKMP2J4QhjOmItFPukp09vnsYQuh2vy7HsRglocDLfntkkow/9w7K+BQ/2I
cArGBxDxIps7k7RVs4UYDWcyndM2tRxEmPSzBCmhsUScBF/F30S5TCCudZdCUfjD+iOlzk7iIYUm
vE1rEbvcryv8vRV+K7QB2cj3daP3+u1pSMXAtGg6OYXF8D8YhOcRac2OzADOiCmekFcQrwvVBSDC
LJNI5dn9hhzPf9YRmC3hOhgoB7ZcOFtW/LQetdnaAcxZ6JgLwkhYCtb05K6sw6pg5aMgryB2aYkp
McmFYwhRE+vX/tofFlSbgC+AEhcosbe6XNKV3UZfCtG/4i4fAcxGjdj3JjnqQWFAGT+da02ynB30
OJxwrRYxL8/AzTdu0BczAJwNDu7yyn7SKRMtvJNSKBKaPI93T3u5R6SDuoD+2ULYy6cvM+FPwilE
khLjsJ6SzQxCwg1AQB05vy/Gx5ryi0YR5zaE0ha67ECEOUGqdNrGaMPLUG4UFo15rPv0dnsdzIwf
WOI6zikS5VBi78UsOTYgesLBk/egB8Awk3hnu3H+Vqgy37+0Cgbt9RNKzrSxSBpZf5g2+N0xC4Ew
vF1n8NAXcIFFZyjYIfJb2QsQPu2pHQndVO8NVPPwSWd0IapQ+tR1Et72yBQ/FX4PC9ktcqvrxTWQ
VdHh8J8eHUW1LEqQeeEmpZMpMKNcVfpVROWfr8Kc4/DTg1/tBxNGmNSwQAQY3AmqV+3Tr5WGYCs3
TtFIvJ4y+JzBNdUf4+ZcSMD4B5kKI9YZu4BvtQPinpkkCKZq9fpmWfoI2Nt35+ewUmGUntaeLd+i
7R+CsT/a7M772jyA6FnGrtmxsMimWwy677RFrvUjOR2U+ZiGYbb06gVqlWP5CVowzAdNgRcPrleT
u10+zy8llhTsa/Ns08LdiksIA3/XAiZmGuT21hZkqOjQrZGUmGlPuWrz8elwtOWTrd0XY6AwTzHB
R6Fos1WAJm4dEn9UR55j9YiDuWpEtKV9Uu85UaewbGVuIcD4yw/uxeelkoA54jV38nkEVzOFlfeC
mK6azriQ7hiLWCGmIvhQgifyJ/X1O3ogP4atNxXBSeCqls/GrI24v3PoyGDZPHtn4GgPBgdP2nyw
iwggChql1Dujwjl4wsmlEP+Vi2iOmKP5Q1vddT3Mroxpg+fxbhwuxEMozGD3tJbpZHXNAEEANbju
Y/aPoPOuENGvZfww2GCQIBVoavQtUCSw7IwZslEGQ8tZ1PAIyhloR2igsInNXRqMKAdI2WEB7nto
EsGXh7zp5kRuf8epVMn7km6DE7taJAWfpkByzg+zsqIHQQcJfTU8dLRkP6sp/G+1Byv3LFxRUOyt
iaOH6MgIBNVjDMxa7jlRMfLRtwLdWK8ZFapGzsXeixTcSENOcnObfr7WUXm2qzQ/tue2s7MY90ix
NMOM7nXt03vhS08BrnGq2Yw1QpGoEEpgUzyAAZrdDwqZKxMpxjKms19Lia9rsrf89lr6pqZkZKud
4XYYf8yRftWcdOSBtJlLyl9EIiSU66ZrJzJnal4ptuMuMkFYZwq7hp9r4ecC9ZVYELCalJUj9YGG
y4lRnQZOIoxy4ZIhdRX6XJqs+aDmJqcGCVKtH02Qd7hbEU9Vu6QARndjVRY1VWsZh01zktRDRmdI
xbG/aRuKn9v5HQwvvp5WdX1chU2kVVi1rtKQbqXlAu+hBNr3N9CRXin3FeKbKL2ORDTrW3eM5Kc1
XZBxD168JLQgoywZLq+/D0TepA7ySTlMj/UMlqzOdESgsxr6CCK6ALex4osoXR3g32YtKSPxuqYP
5klz45ZM30bgmTRBAda4hggZcNsmBHChUGP7Hyh9ilOwPm2BR4m+LGJv8/gzBUhDttySqrJYG+wP
q1kNYAF/SXc3CK/CFjDgSsf27wnWynP0XSQe6qyua1TCnHV/HBtmiik8/JbfikO6Bpvp4b+E6laT
8Cb15WSGvMARzr7K4Ssl+wDy6T+8PxfgiCWnzdb8McenRyimLbOEx8Byqi0l1zu8ujLGdzfIHpOm
Fsr3QGzTkRCUIF+ZfE36A1UIcratnbrzR1nHbulMNfKMEkPFcLs7pwBEYVjyun08Fx1ySVwlUgfS
VqWGOlVys2rB457tqHQAottTmt/kXEicAlbgGzTlJZHI5SpdTlEIX0Uj5o5IY9siXnesmAYJuTqp
AzdM6yQdBG6W2V5wMsqBLlSOoFbEdUPvtTeBm7kRudxTZ9HIf+ke19WT8Ag+2NAN0xnwwTzb0ICJ
LnaqUjLLvqlAhgM4yVMGw/Pr2OO50nBW0mMwxT6ZU+/e4IIaHcFjpLd/ZVIFT7MwjAg+Ymu69c+4
rzS3/95uPboTF0JkXMDeyYB7sWu81h91pJqOB72O/i3T7BLJ1tpeEls/Lw9dHQRC44P+DgIBfy9s
VzL7g9O4v7q40GaSwvx8pEDp/8LmAmus28M18acu7BQfbr3MC6+W4S48ICMrIFXUTPBrO8P4/aZB
a+qdNiKIjwPUqNM1vmGxaTUAi2L8gqO6HIpyMl1udyR/ZXN6y2DG47mjrbe6MmmT631Q7ytQdFDb
0hUK1ABWysYKI++sHt1d8AUE/7AVV+I+EcTfU5FFjqAeeMilF8J7XglkquKpGntRgtL2fnqnaXwE
Z4SAIluIOPLcyca7olJ6DkXEor/aZWJwFoe10Se/bExetWukGDX0NGGKBpk+CV8P10S2/yKHLAhp
lbzZz0wY/YHLJfRL/Dh6/PgJdn1M+ktqL+XEPh0Fh4H9LprmoIwG2vA+lF7fw/V/3yk8A56Xfvxt
MhmHwAl3dAmH0igsU1JlTvU63to5LAvIWRunFA5P5fhw2BW8KncUIFd+e16tjmYin9LZQptjVZ+R
FRiDsLRz8YvYUQ5YcWC3I/5ipYHyKwtiaqFlzk+zltH2CwOR0f/chjdGUFNhiOTtTgdKF9KmzaMy
eetzOPGWUREFIWPgzsiWNbFg1wGSRnYWB4C6QUWUt/kvxZczLZme4Uq5jbOSf1V2/JwABYl0CYOg
t51zQieoiQnykGykvr4/1RZQCmu1g1cbQy779hwXxHCOPgXlaOoGMtctQd9VZZD69QwGvfJMpR7w
vfsD9xrm5YVTTYhIO2gjYD/OLH9txTiF3mHRsftCst/+E9yi3ewiyinPu+GvXNjOiHh/Hx9XD8yZ
p8ZGCR4a4PDszQTtC5tsFGeTVIYzs7UDyzf+mqCpaTndbZ6kgT+p9C02MvaAr59Dv3bvZjMfJ2MD
SY73sjQN2GOvOFPP6fj0Q9Ji88KwjAA5ALN5y98HvZao4WuNOU6rT51kxmmDgE9l2UeNBxCVKa4M
ZII7murBN21BfzmOZJb6KkKvLhKbygKLoxS/6q1hOQBGHsZpbzodx34gBN17IraDHNOfvQuNFENQ
0MC9NxoQ1w3Fis+FdyHxTMCQObEK1BBftr7nkSKOakJPYWLgiEDZFJP2J9+82wUKNFT3Lt2EMjSt
p8RBoYtSmplyW6svosMTj5WhPEyhg9eYTk2YMusCQwFrSUeFo8Ucg+esPngSlmx6kfmQUw/PjjyO
6olZSM6F3Ya06DxFFDVdgOV05n2H6DNHqEGob/Gs0s4Xc1HgSW7vVlBZLIF0ql/CwXNRRUz5agM8
GOygyx40zQsECmeUt1KDwMKXFYjMAeCUKBDKBuopld4ft0U7mdRO0LyNxcmthYs5lm7WdE9ctOLb
krcybak6cqO1y60CJBY7nFFJrrezQuV4gYHnkEky5ae+sQEkHEoSKxRynUdaYsdq52Af4Q1jKd7j
tWoZ0SNHuv8Asq7J9MczoiB23oYPkIo3NO+Lnvk/LPmeCyO0fSAtjPRdmxvBTvb46SqIBcI4yW+W
HASCD1MNxpptDkyKPEGZYVTCfMURpddY3iH7B2PWd7+CBSZ0Z9h0N/NYvAGvns6kfMyb85kdCCek
eSsln3gQZbPCbVw6kZNPQW/UNhethCfD6XcaAAAt+cDHYyAuJBqw1E6LHlwqoH+T6IcwFJ1xNCoX
vLYvH7CyovyogUQRCWKCKeUXohd7nVmm8And3dnTWMckNdUUftrGWLs4eartgJ4qNDmHdEnIhhoh
32MLvxl0B8PhZBmSBcvDDu67ZaCVF/OhpWF0qyvUP3iEcHGdf/50H5ZwvA5QJe1oLURlu9lPEsTz
k1mTNymQVzwoEb6r8HOme1xTQnArCUvIZ2XskZlOHA9D0ohl3m43pjQ/A8LGo9gQSjNIYRmdYf75
NugJhpgGNKkSdOTKxaZK4kEgd3WbfCyRLUSER8WBWzY1Tnb4frhrXy/cGH1J2HNQwXhf/nPNNT35
OmytEGN/urDkHk+R9iZOH8HUCZrVrWLoIkidOoAFGnXOLl3bg0WmZM+zUICTFjZzeCfwn5N3NB20
x1X0/y9gKQwpyh2xXXO+r40dF4ufSuUoHTAR2in7ORlOFeS0/1HR8IsciPBO5P++Sx6iHE+rJka4
OsUrJgJzv4hcH5qGCSAtSpPzSU/LcRbEjDM6XW7DB8ywpoKTyTTeh8VaIa2KfDLjZMUi6gY7aV0u
swT0URMlmX+ToWExMxfnSYxSPYjWaGhO/bZq9AAe6M2AsERxSgs3lVEiTe+g9uiriAo4gcCne+97
9BKzya21OyAukNpPdq0JXSvn7hRFd2wzWYYZgebcvI6xL+bNsV9eOLhHKFopMjdbDuPuLfvtBi8/
I0W0hYrxT9iOxdonOVs5mjkyXzGkFnM4N33383v3AWREW32nkgPUbaiKCG+V3fT1dtvq/6RMQFv+
dGfaSR8vcU2ImUoW9LxDkb0qeupO02Q027bcEqRcz29tmZpyz6sjxG2taYxRNLl8ommEAXBlGS0A
IQh9cOy7X8HSL0eIR2fOG3HS0E+SgyguC8yKSSSf6bYsHgc+8DbuC0foPqO3vtDe/KfPitZvU8Sn
/p2bGc4am/QGJdBlWFa4UrE/GpGnfD8By2Ok9L1o6W3oTE24H1zxpGvVtUdq+Z8LqgbUFP3UPOlK
8wmReqxkonnwLJqcsq5akGnOdqjEDMX/jb3UXKumHFpuBPPMTNb7hX3fLOg1aVYiegi/l2/iLO0+
zYn5QMuHduZwmh90zCdFHGwHtWKxsAY/4r94+a63R04rm6IY6s99ybkd2K1V/NsfhrRKwvgIAAgE
LaV1YTZOyyx3zTxe8aiVcB7uPplboHIdLd1xGi063wYwVQntvE8UOpJDLMZidGatHAjmJeA8k8zD
9aogxJrQi8Z1vMrKHoR4xiAbRWHzyuyAbeKHKXaJMuikpP1buG1AR+zgVq2ii/t4xHxb3q2v9ts1
DoMLq8NPsr5IDj/l5//z2JJOBjmUZEUiBBfNDGZQUt7F5vrhWguluFvCgYSdayVAYJY9hfMYDAhQ
7nGxdxyCWc2P0w/QmEC1N8gMgNQmknyRiTE9JJAxafoX490vPfsdRTH+y28ehWrDdASH33Be5uUd
PW+BVBQoR+ayuD1jO+AhNGPYQFdH+mvv29wJr4NygPMVw1e4CHKH5UGDy58kLCQgs7T1RpMxAb0n
9c8tky76otdE1NvanC7jd3s0ZByWEsK5D3xToHnkHC89uD+KLagNA9TKKaF8xaoAAt40nAlY8xyN
nmXyE/JxImeulvP7+Gg5bN1U0mgExG6tzfhrxHCMClwJ/KpPe2zI2xHp9OvxhXq0jEnDvS26aEYF
HvEtJFMdYg7pkyv9FXtAcfo3Dr6w7QYOdJKZl3OF4wR91KsH1SOicVb4L/eg6Nu6gr0Q8xIagh/K
7Uh7P5G31AxC1HKVLBS8EidWHjGFNVuDjcS9dOiHSTNsRyspeyVZku+kOctutrXFaHVPpPlISWuB
C+SlL44xtfK/oUfWv5m1dTluzVqkmhNcBhzA7RJqF5E7eEpgWM4iLWkaD6KmzMooQ3UwE16Hdn/P
fBQUB9XWFcHegdfwDLI2eGBzNGsDlOdHkRcUqMrWpFh2KD8BY6bnGH0wpuZ7UxgAlsjOHxrOKr1Y
NcwSmYkTy44Ljmk3JJCBwrE3bE0fP++37pvtV8oj9Qw6Xf+8GfcOl82rhYklM8c1ngfdJxNmG/34
NwfdB5O5YI4wL/phxjh25i+I5t992pI1rGW87MKRZK7XgctwuLfwYXA4RZieb+ueY7u1H7CuEKYz
cEaxAv3sLO8Vmpafist/ZoMls9DtS1YVduiOHrnKK+ZJPVdbHZcQNsnenTOiozb99CVz6BQJUiaV
Uv2Z9wcJQ5z5ExhSAv406tY0WwaQo5vDElQtPuqRSRx8QGcQCZHWL0oNit9osjs46c0Ihe9zPLeP
Trmhpal04pVSNIk6hY5uSoMxqurPLMlAjMUFkF+SmVvnu/7418ZJnxzTQS/LpvLW3R+lqzfEhBJS
FyWMmRKby1I2FpuVxt/qVdLRoOZL6t43thxaGxOY7xGAQXcj8u6yatH/YMCbOkBvU9pdvC+MSFW6
t7tM3zMsNObLMQILY+1Xn/CU5LzKxH5YEX7Q76kRhqh7QVF5MVCGDXkxF2V+hMKdrzM2VURjJdzP
ErovmOh7BLhBiZS1FU65/1L7DPtJvIxLWmytgppOvZ+fY7bRHHHlR2zliCbvglEtJdFfbqxs/QVh
MljTXe9Oy42s3B/Q02NW3QI0Xo0ysZYM/CMDdQVoqIqAerXe/B2Nf9+cBi5aGHONjb6jqBe4/d5o
VjiXz7+j2g703IwKXgYvrLGIzOv+BfCL9MNtAWnXaEGFgWkQSzxd5jLxZfzLXFUOgHdxZm0my9h2
ICX3Ihqr58Zw318TKdlHjEzI/wDTfxtUgjiSYmtPrP0/E9VHyrFqnAj1DxhAdZJy/etZNnMclB6b
mBDQk45Y0OtmDFz8LdhwA4aXO5SiFBF/eNUI3niU98kSahORZvD9OFW/LX7sN9MdyDZvzUx5c3Or
GeHNinuKS+BvOz2SeGiq7NyehXfT+fRXjhcZlyMbUxARGdMa+P2yLovtG2S88clwzZ5LrqSMjowf
D+Bghmcm8VHwvsZmSbz+3E4KkRhAm+Z/3npoB+eaoeYsk6heYTPh6TuNVmlPAzM9RpkZMZ5RVpxv
WW13RDOB7+ZWZJlpvfNa8QS6QJxPkHw1E1yMXAAm+1qPg0ztrQx4fvKoLaUJ8S3ccT2pVrKLUf3d
noSr97x4/SkvLoRcAZ37tAENZFhL8b55jmJNrd43L/d9kgCIgWi6edWMezM922ZHOk0cxtuqdHeO
Iz6VQrkG8WZmWtxkXgw8o1fpMbk1GYLCfqXuqGOtdvg9FrglNf2V5hX7897EvZyhVsQsL2Ocpbsp
WVmVYF43ieL9npANrP7hN1MIGOteSM4qwiAUbztaugMPh58qZE02Uknnp31OPmJvIIA/ZLXykGmx
3n4AXsStf0rWqVjrFU1qooxaS7Z5FyZ7GWOdNekFYCSRIb3z0jL/yYMQXjX42TR2W/iL3syJZMSz
JrUfm7twFz0xF2X1kw4H2TVufeVB90iwdc7PTJU8xyWULVLe+7r7H3ywGlknx7Svq2ev7c4tUndd
oG63AfmfWExyIdLAKEent7jx17O+Cq5IvFENXv0hJvHPL8doQXpqsqzbmwQbFoRIlJs1imTF/ST9
yO8elWdG/UEiys3kp3jgq+n8rTEsFg1OnsyZ63pMPZN4XZA+p8sl7WFhbaLdfmeYExzJjPjewhbX
hNlBoVhF3Qoa1rdkWEm8VA1SOg6WHMnJQ8gHds7vdrXhWqvxLb6YhNY1Wc3NEEgnvrkCE73o9Fdb
lPr/CflwAO+WG/7BaRe1AKJ9IeUx23v04F/Etw8SIUGicSGWkNqB0YnmJ15KuFH7uOC9ZnDqbp+4
LkdIOkeqXspuuvVrWnikOuLELNGgF3rycmzu6lVDyvKXY33NkEBysHioSRoMLROlZ2vA6zOO7rl2
ROZoJetDj1VDebDu7yuUQANcfuDSMpKXX2eGXCR6W3r75B4SsVO0iwxC//RJpu9rkINNKxdaeIlI
C2IjlugtsgCW2z2qu/r6Gb57CDeVTOED0mNnuRbgenfZ2Eg5CsWhFWAL65oVna+UHXrg+3CUPaqW
IzN+zK+0Jlmezwd+jUMVyHgwTZPYeiSTaGPz1Ssf3TZT7yI+shy94iHx0yXd9Qreur6mvehzmN9B
CMny5iW+gDI8Bpd6RYmhajiE+FYysXpmSECK5payz9809n+27w13opO0QUnF+NCHvaN9ZjpbcOKI
lHOVgVtB5OhFwuHatMXif1FA239zBbOBPKuaLC/9IYq4eJhDsHJQ89zt/mlU751ymeyARz0bWHUE
EDceY6+EkiJRQ1/8TtY5RhGcvPl8LLsdPhEQRPqUssRs6EcYyU2tb627OXHhU2IHIDgsIIXfzU63
QjigFw0sOyXp8YjBq3i7PBNQyymMgH+v3qOpwQKk2u/diuy5m9eKGHe4hGbRUAaSX8syPsomOdX6
u11o4GVILVPn5JsrKlincSivI+gnEcZupTVC3pmKIdAqXYdtB54990gixTyTagX1lM9eqeHj/Rwi
rgezba4KBOSl6mtLOHvl+B4eP8XTEfizsj7BvWyBashoUhLM0HvzUqLv8mMFvzvV4PldSDFsJsPL
o0bWaXIOsa33TAv2+SnAxgyReELw6uA/iP67VS67JFUM5qIZrGHwnQApxlIpEqOLymykkAzUvLRb
3Dvk4KosLjq8bFfvGaS58WMmP4XtB+3SnxTilETRq32TNdJCNIPqbqKACNUqmFNR0RfEYe/q6i0d
wep4ejShGSYeTpstXW/KZj7DcfHLU1PjBROthEsuIzaBlV6FY5jopef8ApeBLiKzDLGE0KCPzKFZ
Eti6idto5Zd0P9nozuYAwuAYLAcO0acXUXBrmw/uV848uWbuJjSlLN8wucZijCJB9Z8qKzH+Wfg4
RWB9PBczMzh/gkuvrkrFJ0diQRLfeWwzmg+YiQpBZYu24qjb/8e6ugZiSe/YcOHzA8Hcwu3Xu48+
5o6EzW2Q0bN19olM2vDyxixElx7Sf1cOh5UOU+HXfI0voy3wnctu3enzp3X9sJSFoqhLYxTykpOp
qxLyjY+iDahsL2JW7YDaaPK/NGv8nK1el3rE5YU9xWzZ7w66p6LjGyaOVqjpntjwgQ5gI5eRNS8O
wBM2FVfJ7EjKr+Hon8wWjgOPB+L9oPCDpQYE+sx7XvJOYm8d0thUREOGdpMb0PmKENvjRDXwptH1
pVPiOM+3kP0X1GMcLw24rFqBs9E1wrH36V4qLzmL8LcEjvjFzWpVL+WmLHah36doMRurZCH3YMgk
I6LOMXuPgkXjcB0NG6Y/HDw71Mzq80issxZaYgBY9ppF3ouyFwMlVaIAoptn6o3ur+m03JbyiaaJ
nixoNGRiysla03Vf2oEagg+VYHNFnEne9UyU6QSsIYTm7hByH4G3f0qrW+VBL2NQ+yMjDnw2sNFb
CZ/koJkEH1+lWWJ9mey1NpGHrtjh81ICczR+w6w8Opbyj/Y3PNU2/wEAA9DaJv7TebeyfsLtx2Vq
wrlCZtg7gR8cpjxIMivLIlypbCO47GCjsVa9cfxXR4i8t6bYSlaNhLIuzPeTOQzwzINZBSn50r4+
thxtEn3UBxNBw1Iizw9krqMiRJnj2IklcTL8QnUvdLSvV+v941pqYatxP3pm4IVzmJmC2L2/4NWh
A2oqc33lYUgEgighEOI4u29efAVwIzOkSbLgWqCcVUuhU5wvVVAGFB0pM8S60giOXe2vqlzKJJMz
slp3XhfrI0tHYRYRPLPEXLghaRDGFZPeDoa8foAyX+TDFJpHPLrTl/C04LnUPMr04UhT5np6jIZ4
DozIp5jpXDVLdBZqsLVBk6R26gWAyWva9oQiZ4+92NwgsB5v+JI4EGEMK3A0ytFTLqsGEuwbC5v/
SdoLFQP/WDTkl9JLiJan0aJT3mo2+Np+XqYDomlJiBiXmMxkTIasp4VlRu5HH5powu/INi2xmUHL
CsGF+QB8sqP1fK+ncIzls4uyY5nK/RWVgw8LdYeynPl3QNL7jYOM8LT1QVNMlqINKevgWruCCgVi
d0uVnGI+V/UHvk2k5i91NH6ECeimqokuNMeQbrnnqhdmNvJGyOQ08uDBm5Q4lsm5LU+3oaKvFGVv
26Q9TacfDzm/9rspNjL1ZoQ9p9qDePZ9pIduz3f/+9QM35JILW3k5go6nk941kLzBfcBoUvxhL6/
SSy3VYf2JIxkxDTR2qeaayuIIj0lJJEe91rT6um2yRS/9qGjODTWJzKHHSn1NtbMUnxvvc5zo3Bw
Rm/HLQX1PIUDGHR+QUNyDNiZqsXSDbswhJhOFHEcXrhblOekrj4CT1f3/iIHVWd7lCcplTaaQNO/
1zTK0Ql5Bu9tgxLTppw2v2yL//swQ01eAOzhdFv0BqAwWHQrhq4+WznuVaMV5nx9VwcZLBNjljgI
yto9U6cO+qeYCV9u0eYwBzg4DNiQ5qcQezqdIo+0x/frPTOb0KA2+0/ATJhlfTnzDG766lHVG0Ys
lvmBljPuTXyiY8d40fwsnoDTM90es4iQFiL2+zab5ihPhdaLzuKLNFchCzYPVhrQ0xACwc8bcS0a
KQ9EZv/aLjSxOpLKF8DvANBOKzDrEt87bU4Zsx9LyVVOU8yBcpFYvuEX4XAumHyREuBhw2T9gUJi
Q2n+sZ1jwSRN2cXIsuyPpqgg4q21lVIfR2olgOkRuWsPfqSGEFoMa9ZPNsu2bC1kBT59N68HdWno
I1m4TCpqfyXJSmlDqwH1ElU7m0a/aCyKPFFtq0CCd7/EoujwwjMLcPj4ZUVX0VxmYRSeIAH1B88a
6BCAn3QujZE6tAYvmzOMp0ZSSDpVAk23ue5j9Ha6Xqd7jtgL9kMqApkIc48Quq+qyNsJ4YYyjCIL
Tjgtb8PDewZvojPSgsYzp1h1NIRGEXUB3jufHUV8MTqF2B9FXLFoVnUpouChe/oiIBf2cjr4vNd1
MZWFbOVclpYP1fdVy/CYKoTp96gpcCZt3SjHj8rkMBFOWsannuFMf0rAHm7hkHY46lDCPyME0xZI
pPW7NYJalT7kHgX9PEFopVy/SxtXRYMDFIwc0UYxs5fC5YgcpUH0X2NAwvgZacsnruCOU0docH2c
7YS0UurerFT5TLvJlJGhq6SGjsc/QHefGK7miMyjS5e1SUqphaGBl8ytieWfwp5t/GGZZEMPuk/f
vYlxwx4wBRhXxxOfA8nIMoA5ncBusJ/aBakgvVoUtqiJrPVLibrWAbDiA35m0qY5O/3bMBQyYp1M
KUXq0VCrcpZIzj1ljObUDK9EdcVZAgnyCpcpLDf0qS0Hw68f2nshZ7XM4DbRmP6SijDSdYB7Mmm5
WNIJf5TwLcqZUlVZbo3zvGlq57Ufds06Lvoo1E2fA02ZN7fL6ENM6jK2TuszU96WvibdKlELIW5v
/9E4Bc+29F6ns8DVIWTOzxFpJG5K0IAribmvCi/B1HGnfHe/1tJI0163YbTe6Anq50CkfLaIqH6J
P8U/S8/3wnqX208eXNR0pq7FFzH2qVgtTjSHClr4TQaMs7qqP0r0S2gfKZrevWXhKUW0RHPuq1gL
WCMS2ZB57hvJusndUiM+xjC9oIXhpqo21KVTdP8LmheirU4vsQKZWtG5Ht/Z5cC8ExXVR0P8+6Er
ewIcsvc1fRM2j5AwCy9Oa4rClZcf7hwXMsp9jtWEaZmCBW/gCW2yRlx34pEcdBGJZD0GK9t02C+h
JjovmXpA84sgY2JWMFlFnP0RbwO/1fNP40f86YjvmCeEn2pGMdp1qFHDYtbZP/2LZXVPIm9yqk5R
1XclotQ3/4gOCdhNI0DbynGI+SxfdHbv/Pl1HTrFz0JzjWNJC8Kbx1VFMb4VfuLDam/Cyanh40zx
XezlvxFfE0lzIldI9BFk46TI353A9ekFzBlA2Rw1Dlii7XeZClBA2TJcfPYinaJtPk1awTzm3PFU
pR8ILhv7WmE85wvMhcs0zMWF+SpAeJ9vI37rY8RJfC0MFiL9JS2T3ly3o58W3hWAnL7zZWAm7Uqe
dFIOlbv5zK6d3/8B2+xw8mMZl6ahV3bDpxrRyEAZkUwVuyUtSsSaBbGwNcAH8y2dOvd1fmGv5UL+
uZKtL79L/31/z/rA81U7vs+aOL25HDR10h4m+MEimkmlfhnnO3QSGqkvs5U7b+BC4SYDsrSvSWM0
v1BkeEixvhN84MYEVZH/h3XhbfqBeecOaH5s8BEutn/YRN2CHsZt+55w+lo2N8eePsPaeIZeHd5o
3gq74dgmqIuE53JuymHZMer5PX00pfZtvffamSlLGukDctt2H6oD9N62eQ9+LElqsHz9yZF4uUR3
dqPmZvuoeSkT/XqIjh04T8qe+x1OXkI/KWWsA71EPBgc4+uZ6JI6kxXTRO3ICDT6KeNMwD5L2RAx
CSxmziQ+VQ4zxKDA+GB2idhKAPwklkP2RJ+S13Rv5CmIHZI6jpPkRT9ikJoO3tMyogm+gvpcbMKb
PUySQ2KE2ERm5NIQhdQmOq/gMRoi+OdwOoMXmpEIIjzSFjk0hlxIoo9onsi4ttPMbBVm5p5llVuO
CqMNFvDwwe7ntqWz8UNpbx47d7m8SOuppbfNyv8cgCjlbie9f19TycOX+fcVfj68ox0PtEN7lerw
OJZSpnAAxCxoUlr2PKqspALsVX44JxlIvEMpk5xaSE+RYVLCByZK+033pglU7IL1rdvWG4Kw79l2
S6qrQZyXKVV2d2IrCdszRtPQ9JDu+wUNecKpFAF3a6pbsT7Z6JbJJ4ianQPjquWZKqtU7hLo0MkN
sv2SDzNGMzGprS/1EzJYX7L+6td2wR0iH4WtBGCKX3JK7JWGho3ga6inC41jPmjBsb09rx+4p89R
I6Mv9bIOm6bQc1+7j5AieZNV7MRiHosCCbBq/Sa0AMxRkpSdvResnSmX1L6MvXlDnZozfG8Z/MNH
kudPv3YVui/DOUb0/5LMhnsxn28GWYuXyGbK1u2TgX+KO1IXm9twh0tat6GXRPDFPGKcVYgrhX1T
uluWHYfJCOcXUsSjYlw6Tp15ddU59LdSsLvDLJJPTscJAmOTJof5uiNzIHjUT+pG6KaSIIOLBKhF
q8sZC5zmjf5zVNWmvKcbpeFOowXPLjLEfWVMNj/uPjT8gy4rygx2ntFYSjs14ooaE0eTHAAF39Ne
yToMqAUKs9FZGwSdNCVq1qoT4RffWmRg0sP7VjFAPs2ubl80a2GN3d4gbpPjOyeeKss11iL4v1mI
FKgLDpg+2CMrSK50h2gbpe3/HRnEJwUqJlBd2CO3VkM/qyNKOKeA80ujkGbmoyIH18bTmmguPTxx
RP0dSvqaPhmb4ZsKyoy0yQrElarLoTBDJT3D1xqws5fYeBqEt6ofbcs/DrVdHFTX+IWxidHvlKlw
OTFFIyJXMoYfrr1+G3Uc38tUx+fMzdSj8tdl9jKpDMSnmmH0E+ChdcoyhSFGtsMHitycnjwTs02c
h6M6IbuAx6+YiHmXeKN6gvp1UzTB3UWd1QVjJQ9EFw3NaxlOuK4ocFjd+i9z4V6W0qWu5ppfQcxz
Yv6QinmrshHU62xgqg6qEdMl6HBJRKFxu3vgRUxpr9ncj73mt3Y2qdUuSqovUxbg4qlYad/P5jdv
ZnM2AJqpzHAXRMPUH0HhgpA+DBKEjohBbrKk/Tb50hb9Aojnmn2pttWBtA3cRTvg+EoYrn9FwvR7
AYsllN2UbAOnBiDbLh1rm4R87yEfMeGZFXZQOX4nAXh8KlVqYqRfYYGu4SitO2sANcGhfuweCj0l
3mlJAJ6+GektvvAK9+vzwbQJQXjibi+cPlPOpcP4uHPUlGAozCbQVFfYYZ7B+hJPG2rNeJbtP7SS
DRCd2gmZCIE2vMDQA+wRrFHq8aOwZyMFOOXn5IXocuYs93pXpJJXjN8qEPDKHd9XFlLxZoxp2WE2
QS8GuQ1wp4vlrnWWjQqmEXv+k/TtvkBC5YXqwbGnq9haq5AVcqD0euud1SIl1jAAwm4VV29DxE9f
oGs6NagI4BNEXDmqvmaU0z2BbrMGMQy6uAB5SWDy6gWloFZFZ9UlvRnv18psgqq7+lQhOFYkj5UU
FiwpfydYVDNMnISCMBLbceO0tdlS4AelUs0IJq0Gn9hakdVP4YnKDP6RvxQXS4FObXbvu02jcsv1
KqNH4ZAAzWyksuS+0xp3hC3V3ldwBfefhsK8qnmEJP0JY597oWS2sSosLwRWb1ZYizWn91qas622
TADzTh0aHXPCNyEaTXR5XvCpBwT+mUlACEbVmp/mNMHXTLmIBG6lfSV1OQqziticKYKCprwroWVH
cxH1rDKpqJm/dQ0QXx3xTstmZVn3FE1RM1rRPPRlJtvVeuPTjZws4kICPRztDxBRJwLgzBYSJW/s
/uXLCSRGEzyBUeKK/tpA79SXz4AwMKmY2plhDvAU/02EYs0JMTbSEYN8D7nqJHXFYkJoGUuS8tz+
QlGslWrvtris0iam/C/dh8jS/bIONyfAi64vt9yQlTEkGw9w3vy5UeWJ7JVTzWbs9uHO74PThNEd
iRlNrmOF+tSU95kLsirdJauT3gnh2e9SFhDJntt5mnRcQlrC+d62q8RiP5SEsntLgsEaBGJsgcyC
7cp3P4Sl3rkBmYSuUAkOsD3MYsAzJfyurqTxr5brgFRvOuxCLhY1gsfX4LlcPD7iFi/tGfdQaxW4
BpeKysyyL22MlCiKpUIkQ5BGDYUA749Igfd4un0E6N0LH21TgEFkySVipRPi/ZNRfp+BrwFJlaKq
A/qVkyHaAiV1dj2XoTL/AS48TR6HZfxM9kbW1XrXCbqt7yQZaNC0WkehSSHkBpYTRYtNPHkatKna
ZF3nALfNu03KnHUurO/OCbgxQ5r6cbVcCKinDiooRiLp4uFcEsoxtzlhhQJzk6ZsmPk8aFT/y9YK
Mtr/eS/aMz9miHN+v+D8OU9pPpKQoSRSWoEEZSlkP++QpJbZM53/KDmi6LDukkt9TvhXdbEVoEYl
fS4nXUonN2r2EjXsCB383UTHdBphg3fAkBUQaGgTGY4iCLrNweB+gJk78q+U2fcRLsuhZwnAOoSS
bmRfVMcSRMeBDlgdeRcaWaujWGJf6RsOMX87TXBIVrITdHWEYBxioykUKeut0GihbNIOSbf8vY6j
uYXtUxiRm8KaV8a07wG5NZmwTFx3dYCpnCDyfGmdffScBpxCjgs0LDgMOr/8XpzSoumbGCW734GL
0FvuohxgStvJuLcAbP++eTd9M5UC/2eB8TNBgYBcqLJ6DNd47VPwD4Cnvi9SGbSkF1AJYDiJasTT
3tHMODTzX9WsFonngo80S3EYDuzbjtvF2YYsZK+gs2cPYuonj58LUdrce5WS7yd3O7xFXRs3uEp3
wc5hSO/k0vUw6e+LiZYfM0KLzIBct58lv52UbBqJOTJK8X3HDS+sJPOSNd8urcvWaDQcpQCMIlEW
Wb9EiljQkDEjAx5btglIldcd4BVMoZF+IRum8C5efDq2hjsrB5ac9knl+Yx1occE6A1TNwzm/sUd
yo/MgA2f5uPAkptdBhVbt0jxv2yFdJsHXmtDcMrvLcP3L7mECBA/jH18utWDQVsC/eGBKllRhMsF
0aAJiUtW05ynrN4XF23EmBIIeMxXhaUwtZCn0d/mS+CoDfbAvpBbIhpcZfoOy5zmvamigAwf4HPJ
FTpnIsMS6HzYt33KDKWVsWv1UP64unGmET8lnOaEsHsCXgtxwyu+agYGj4vti2+rkHvBHp66xjo8
SAx05X4NnkzohFUim75gaWD8lI8SW9vxPJxEktSXux6oFRSkEsRLta1tik2EgmolvYmFD/Z5U9D/
99V+je51S9LX8K53dyeSdFZKEhrMZJxsVmfdh24yf+QKOIie/xnneLKHfonAJDXH2nCnzn6CZKmf
Gb2Y6w59R8ohaxI4sh7Z46AT3BLBTWUeG0aPKYjA7nHYl4Fd/T9STTlBeVW3NFZO7EB1WwZJ10e0
NKxdGrWwbTRe0lpK4f3EjRpsGcCxwsxLwNTzOik4Mn8IYvIGOfyxpoHUMP5Gy3JFu3WyUN5FGM9b
iw3oXMLKBz3whty8onkwlRhQ4fWOyTulcVJ397RwK/MasPcYxk9HNTEEqyxPCVPI65rjwAyZXpSf
eyvLXUGCoc6Taqjh2k7Ii/MFG3IKtHFseaI9EjPeXjhNhZxsvdH1gV1vuJTFMBx/tf297JjK5LCi
c5no25c12b5LyQT0zGY9LoE11lktdyQyqSWiZr7DenFnJ9bmNEDTh/cxzt/5L0gSRTEjNejRQlvb
L+VcmiZJnLxuOke8fLOeJo649v3ciMJ0r2dlthrXOyY2S44kTEVBgMRb0zmYLDHynHWpA+zrq87F
yzskqwihwUPsgJvKPkeD/gLWCOWp0/e3DoRhU2tGw+4jo1v8pvykuQRTjV3LT8ME4wk9gAPhkqvF
8nxBUTupYyuAf2liv2x0Oa/EKflDCmSnZh6d51Pv3xxERDPb7/qxsPAp81j+3T4GyhM6WUblcVOL
1FuxgToxIA8vAAMVqjlZI7hTgEvALFpeWKvvTzSB1uN6gqHXuxNgR/5qXAlmHk4a6D07tR3B59D5
IuEVaOHeP6iKfWkz5sEQbJprMzsiujtTNbYIacaylpCzfPpvCEc+I1XwmZHkYXKal/t9WjeBEPo5
k5G8QA018CbntfqGqy03fPaT6H36HJIfUKIOkY6EZH56+ps4EtEecYjgjepr1WzRIxGqAFPoCQN2
E6W4EiS9EHQqLjyPzodIr1WBmh0ZK3mkWgNuw83e7YaTYDrzS2x1vzYIpDe2dlBwzlE9WHWTCpG6
aHp3bRyKYpB380QqN5K7MdbUanJHeFnzoWn8z2BPexB5wylr/tq2kU1IhU63JIgyEMCE/VFV2R+N
CC/klrozArflseH5H7arkwrF+2e0PXIZoxQcDWtffsZkgk9ZwPOj6t32Fj3rVGfyhlka178rxa2a
aSIQawhSiapOTcxRdOYP7EfeTLPIJ+gjIL0R40A6T+PG/9yUD9tf0EfJNVv2BB5Qz/6sSDL7nXtd
LYrEVSaa1Z5nqvlK4J5AsS9zweHYOR94bmI7+1+sUK3cjJa2Z63XXumU9Kw6JZaKKg1bhrUKT554
LOn7DlmhcM5DsG88ievLHpcwH8ioDYkt+2w0wp+tRShGTHv+j0DULxOy3qIsiO/LSIxSpLzlbsqF
Ah9gdxOqyU7Olq3HK2t4G0XEkKI9VzLhwsgWLyMPraFQ+uglKKVDt6oD8brM7OzsGuJQGpSDyHfY
gLd+5eZ4TT6bpH0BzEmkk3Hn/FcsM0b/IAyLdF2YTBMNF8/G3x22ksVOiq9R3BkK4wXKYPSPGKLt
BuoOu1NrvgMNoz35fhAzCyrUxqY350s73BSj1q/0XmubBwO8LWY21IHpBrrZEScP/3p50pKEG6Uw
HeTd7Ptu/xxg5KL+/qvre94LeMfz39Uz2nHtsa+HihB2mW36i8D3gaS8Ljo7EXzM3qB/MqgGrps9
EqRIo+RRObEqhpwD7tunBFWtZ/en/kwmX+M73LxyANJ0y3NYlmZGv6W5++m96YLqR+dkrJmyEfQa
ybfmZBMAJr7T8JipGqgL+f0WXacPddffh/WH6DFJCNMsayseI45MjCnPNOyrJpAax8j1cdZVA+pr
rwc//4Yq8tk+H6lC94tDfRd3DUEE42PlFlT4oFLTYV7vtZ5zmY36tsy0YvEUIzPd6TeIJUqbouSF
KaJpKFsl+s/Y/mOAYSzdhUwWu4vKqWWYyHfdDABfqDj6rCXdiH/q8pbQoTeU0liX5ETzbcRlXPq1
JJowhnpSewEDIg5EWiyP92bUXjTvtA09SySYzjHpZLyWgUqlsZnPi1aw62YCJR5WXfk5blGory0P
7bTvEjGzlxtUvc6b7+jgx/sdEoAhJj72lVa6rmJlCNGKCyBQ8Uhigmj0deRG5175ByrpK1gW9lR5
GKFMI9SFDoudS+6VIR1axdDH8eQFDrKWYtcgFG0wvwmgUpmR2gNsrQuXeGsrqwX5hD3khsrIExIr
9zMmQ4jUZCM4WZWlJlVtEHNATk03hi21HyZ6xn9/ijyydSEeTODvFAkCLKE6NuFC/TqqnYpmLWyh
i2tozn5L03Rc8FnbouEW4BJnBB++9smJ1T49+XnPMmuWtrp1hu72Xa5asVnqwR8xQ34v6/YHAoti
5rUJ2rQTD7ACk0u/4SFSODfij6pTRl4K+HxyHiUpGkvucITd+DJy8tQbfKpoPlE3KS5jw77drmsZ
hIfHuzw3MWiWkex9+t/Wtej+R086Y8uoo4OB2SBFKS9+k8+4Un1zSrXoFhFflfbfnldcAuVSmPLJ
nOQR9a/qhAEEuH/sGbo751Mbs2mIC+n048niWmB1tmDi1EbgSngsNKK6V+YiFjH/5LDyrVp7DANa
tUhbr6KTgk/H7ytzdAvdzgUSgsO76gkdXbcQcOoEd2XzHy4WbK0yWdl7jy8IDgSLdHt+UwAGes9S
VN4AQUoLSIVjCNIOsDCC+bv4reClxULzl6tP+FeLkfa9YXWmmtieeCGFls2tVr7MalUqDuqJ9O3v
Z1obysHsL3PbXO7lJOeIKoRS4XHD7KhPJ8LvKUxSSh/s8bbq4k9dQSlHFaUMt5NUX3czzh4FSnhO
SaRDui3XHeNtmrS74nrw1etJqNJ6GUsgvCxMwYkqthCRnM17hNIikomI/pPkOhiuHOLLriwVzjHl
lsv+TqdQDTdZd1MCxMj4ebKXD8552aJy6wAIR9f38l9jBTcWe0XAaMA4bjI7EL/U0BK7ixeAE8tl
pV3EYxawXS3o8+0N7mlwLr/EE1gbUcNPNw/pd41b5NWa7G4K9eAHVEl1AlbsqhC+jdtF5gxTkjeG
jTBqiO5iDPnaQXXMiIaj9Anbx1nvkUQQUMYF5TY7gb6ImlI8WVwSggMD8kVn6h1eBEG/F+w3VgBt
1Bq+H9HnVZtEXFCm960h4z4L97raptDQ24QQxtGiOEMYgkbXei4MDiZ/UcgR1BUrFeQ6A5tF7Fiz
hCMC+WgMAYIjCCc5GvDBqpvoXiZ7OLXrrZM/BEa7Jeez+gqKDNp2zSEYFZF0GBbQLclYMDvEbqHE
T/Rre8kGrk+TYwZYCdgqIzCB2m/otfdcij/YWFG4/lbXIGDCVjtndNRdVSKBeEyZUe1NjsCQG/xk
lFvqolMEOnNvD+RBNMg6VpVcUKYsS2KAY3qu4ampaeRtxpqym4SF+jYN69yAC4/7U+q37V+/rgyQ
T0kDv5ZBDmPpY6DR0n0fyOn0hKxyA67dD/JjcaG0bcc8TN5wYJ2TA9UB0tTAxBvsbe45T5mc9FpM
PjYU3kCE3zKtD3PAD3WLBA9G80aZyjckfy+IkGXJI8IB82/ddTrXD+/qgdASnFP3jrZyOAE48lCO
U9Myf+KZ1OyFU4Ysco+stRFuMUOG468aXKFhcoDu2mzWohBtm/5Rs3Y7E6hRqcHlzc6yP2nqucRo
oadcLI3HmuO3wf9rCQS06hb888V0mwaDfLzj7EiZbvV+2MTwHHEfaeiNBWFiZ8fFkNbDpz4A7Mp9
tVjoRGTyAs6rdNJKPC30wsazQnxU2qbEwFjc01J2t+OLwXOrioaYAfhMYbenzzLXCmrbHIq0IGDC
sbnswlHAyfVQPw9GbLuZUSAKJD3nvqlAPDubVp9RwnE/G41yIjFP0xnKWND543dNJ4wbv60EKQ9P
+aMvHzk0Jpx7qniMdvXSJbKlABzGUHlEJ2Pg1z9dHAk6iUZS2jDvHxmgB6n8y6gfD5CyGu4G6ZwZ
E4TsIQenM7Skvi8+tm4x8QFS8boGjM6UHoqrg76bqQhhwSjCeLZzmrRstJ5whcvboSifbZ8gPsUa
0xVqFFFYoQZ0MhdttX52mCSCwbPOj7snB6A+oHTfkZEHDfh4PJsVKfrW5JxxpNuU3a/gzBkQwmyW
oLlx9ceg87VkEuRPZYf8Wp7sqItNAfVjvU2J+M9/sM7Vxs2H54BFWOdy1pvdcdirNGwVbEBnKYZx
B3yP/gkXRdkbTd2swJdptipN1uAYX1ruB0jXpQ8p9s6WnkBJ83kOt1vVSYDCF+veLx0J23cpMJuo
1KQridIc1zj5rP0T66wZS7GNkKw6eDcm/TD/Ftd2bI6j1/BJzGmu1Sux98PtyzFVZS9mX2sMmK5d
h90Z3f1KGDexA/BnKoh9eG5uM0WOgHvkIdT2pi6X038EBYD7k4rW6m8K6MKfqhZn4DeMdPnsAvMo
K3buw1vYc/EjcCmyX/r+9iISh/yTSkv3234cMEqV3yE8TCVToy2CRsafjb8xCcn015tIacfySBXO
KUq7z2xyFw0xhgFqKkTpKjWJGZOHK4fmHSHLsh8wc6t1dE5f5igX5UibAUIheT3FGttce8p8jarY
B3rNMsTJcqWxb6Wb0M6JfEI/jdKb2yB0NBsyfAU8wZP2BGqsTcVW6yfkVT7Z2IHfOYQTV6/Ni9zj
4SKo97+RAYjUtm8wY2AcHvqSGrYKgfdtkjAoZMKIHOKoBBkQyH0MWZul56us9AJ6vGn6iavqod+9
abXmaQHHw2zUp1u5gJ1jIEoTq5b5TPnMXx6oi4qfoqQlKe4FGU7x0GkrxwOEWNzDQfx5hEPAQx6u
f/u/t8c4MLkWHELxib465/9LO3e99HU8vL5l2ijaUWnMgG6VpqoCL+YQkG4Aqd+7ZygrKOYanmtI
W4IFDEzLBx3av4J7S2ohZlARoQVzxd3htRYJ4wr5Y4fhssx3VOxiqSTWgWFiB53U6cSSHukQ4g5H
moGVgU9CL++HaIt3wY7WgPVs0ITHBoZrKl+0ZsQIGAUIAa+PIM+YzTe64UCjMm5e8JzMu0gPA98E
PqoJ0myJLJRNqGl66KG57EEQV0dHn46BpRE6lLJXiVPno+PmgyPsaIb+OeKiPK8Tp7BYA2iIJ93i
GjXdEHcusQXvw3B9HPw1mjB9d3OrNC5Q4DopnUM2zPFc9GLTRQ0aXnG5XJa+P8Wh7lxztXduwXkE
yubNuVeB9IbvEPbpeiPwdS6/KfgbJdLObD4RBPzgRJfRO6T/+nJyeXSkXChCPjDFH+DaFGzI+cnB
FAH66PgmbHj50PcsFRCJKdLfqH9TFye0AK4XQ2EYxP2U7Mg8yNvhA5La4+xlsz2sL6TTU7V2utyf
k/6x6XHdBDHwMuuVBa/pVoq/Tpu3OHLYGe1rHp/tlZWJKaTJp1g/6rcwxB1+wTBKZMW9uaePxWSp
rDf2kf9Hvd+emshPH6/teOq2TajKTvmrA3q4VIeX1OWWHs2gHqNnpujs3cDNqBvVZ2OuTNBUxXUM
NsybzGjbtWHrPXbc57xA2/RJMHw1fe48a6BYhcH6H5keMkGqHcwOZOywF1XjhUW8z8czlTxjyMSl
saNMDKAbTj+AIbzPCViRlyWJ0Ny15gb+3+yJEXw9syNiCnEKybW6nN4nc0nILjwb+HLXEA1r7x+I
pjIugYfOVqlsAW1iCYg844zd0FydWcxhy/IGCAqGRuU9C3nl1QVkK+UeHuMHcLVYBWxo4LsktF31
85lF6QuFO8gwhsmmY9l3X0KdshXCqKj/DTQ2zb7X6wetlYRNM1cvbjW/pUbdm7qocySyxg1iOous
+zwV1VLFdJ/VMvVqsyVancmk+WGOKiZoMTklzm7ICH6pBiqyLsrQek9UG5VV0/ysHsNf5fCN91go
C8safD1aAo4xQ4hQSTEph/OaDFa8zHZmuUM3Pkg9t4dc+/+4xZZxKrSnOMOvHPA6tnMtkKlmSNIf
18Cfj0scfRVSU5HlmRJ8FJfdNkOG4wVPQmXTA7zPrjgygTfibI7H+Rh6AkWk0HWh6U3Q0UlJqBsa
mx6N4ya4scp1zhNbCDg6jAcJSU1pvNe267K5ChUlyxtAA98fPjZSIgHdjPDQulxEJNvODVVTgpNp
8c8FVIN3uUZ03TVC+4gVAaEiTbUvmMe99wYczFGrxhlSuBTL181EstuQGC8sR4QXlyBNvSNoTOh+
GS/11mNfYDPKJMZ0cxffVlUg7cfzUkJk8FbOnup+LeOtu9w859nT1VDJMKoXMhRNw//V1ogM/7J7
JnunM15h7C1qWDdqx4w6DMGdR8d7CYUi/ZF2yjNPHi3ci10f26ynEYZ/ZtmLPPHVKm3UQfdfn4gZ
u1E3GNhpu9vTTBoL0x2V5GmngymBEfk5n86y2MW3SoOZXOmq/XyKMVe04bLpGGMKPtHNLw8Hc0Ql
zB0HfctX3jDzgdV0gvzt+ndEQZDnnooGe2nEiYDU1a8JCIUdS+FVuISnrYSabx4FAEL6o0o+4xCa
DB+LgLSwwO8E+r+S0hIZdW+l2W4gpR0Hqz2cuLb1iOZn2y4nkuW+Y4If0/tITZb4GymYiBvvJEoG
6WuBzAT+aw8Ucszc/IpW0uBSwq3scdtimQP5twR78MR6VojOpUvg7WZ9FSLSV7P4nY5imYZxaz6Y
4ozdcdY2MO/Mks3v8TWmMWCKaPMnNn5f5QS+unJTHnwKkevAtYcuKsJlKuZiONWzHcsYOViKjHCb
Jh6k4hUA4WwB45ydt4kIYSXCioLdWbnr20NJkfSEdHM69SUFyACW325wPIT8jGY6/OvVsdYh/XDC
Sz9r41GXkic+6JASVnTCOFJiqYZSS2GNwq99spM+EH0cAms7DYbXHUdkMStXvMiDOZfR6QBtgNco
r9ARMO/qgKO0L5Or956z2b2O1Cx+iAvKPqhmYvU04oMjH5iFSdaH8GR617A0yAdS67ujC2EO8bu+
LF3iw5iPZSiSjs9ofXqrT2m0Bi8CyP+8p5KCyJuQWfVU/b8xiBuwJtssQlbOPDvyjxgKkDAAtK2N
Cr75lHEmU007L4w4WusZYOSGg8wmezx4VQ1KA53otwpOuohDS2tG/Zxfi54HDSsOvlyp438jAh2w
1ju+W+SvHe/qOhT1OZ6dDoCjOtMS66qiT6j5OJBNSyPKp7tLwZRGtcY1evqlUaCizq9j2O0sE0aF
hmyfS7YI4WliCf0RW8nBpmQuIfyY7LAl5vEPnuiPh5BQNH3RmZLmNH5vk9VGxq+DD50kUVeYNFlX
ALHhvmEV7T3yVq4vxjKSgfrHJo2GzKiLYtsaIeFWw589OfcMs/S765Ghsif9PbX7/pS2+v2QEftu
rA9Dw+V5zUge4UwJD1z+BSjXBpg8vny3U55KEu2XS/6nBf+yzR5GJJ0HwgWKADCpJ7aAKwF5lAfH
/wG3/ZPhTjS24ntXG01kpSavAo2Am/z0RWI8IcXK6ZpHPQp1UAq8373z2bISelNzvej8AlEWFV/W
BnnnFiD3umlVLXgnEUSzqmo09PZ9FDfugIBnfAFuPQQZLX2V+eu8t6tGswSLzpqq2DtLULOgihwR
jmkV+xyrOpEfaXkO32S+jBt+ENEmhs2frHokTsSJ5lNDfe/m0RrPzUvr2PRmxPG7w0zsdQlhI/L9
ZQwc67nf8MdSVI33jO/2ZlNE4KYMRFiwWiQhFi6S5e816wUYe5m3/X6zEhw8aXUXlgrqXVTjK5yO
bKCmFrtsxF3nuLYqK2fldxHo6OCxzNRLKUyNjBejBRADp8yuts+7vLiKq2Z2D13/asmAACEThZW2
RxD0lUvZZbelHlSMLXQ3qU0tpLZsJyYNRPSa33w4uQTGF/lMleJQ6xyrBmoNxb657paW3Eofzgni
cGGpKxUOaHNRrA7V0rryNLKdHxVE/QCVduiKeh72yBwAEWSa2TTJydAR+mWrcn0j9ehe3FpDail5
omnT4ZI8ajhyF5sY7LEjtO09wTrCAn49vP04NxXHpYn0BlOH4OwXe8MvDgO9Av+5gykZUnRYoFJQ
ZoNpQc4tVZ9Wh2WtTeZHLJ+eE5aAvYbmysuvlxGU8gYLWBUfxzqWuyr5bxQXac5vtdi4+1cDkqx/
TiA64Y/ScHPkJGqXW94NqBI9IkNo4LbhWpa4PVlCVe2r1cn2lA8Dz+DitUnGLyDhE2FrKhHck50H
5NHuUtorFgqTQPdKpZwK69bn/4xxqIO632HPtr7bgztOaeE5OTOmCT3WpJv+s7I2hrs20e7p/kWm
OT4+/NcBToFtEsfvgSWeDPR5lwH9zeLdTVJy7G7kVvr2WGDNcUDYLt60zPPM/b+/1aAVSadXfL9y
2vxFDpoW+mAMoT0FsyvYWqheeI4Oze3pvjzLJj9ZQO8l71c7t2WSLEMNTaT+ibBm4zql5CjDi5Cq
8IrepPTUBlNF3/OmAb1BBs256+xjV/BggTzsZTMw5qIGzSt3b2ZFR5DJn+ONyq97ujV4YRKz8/p3
a7pLJwm7QLAgvewpDbl7/BfZKKxyXlH4euzJ3WRU21RU0EcDuI7GLsXAKOjX0zKxk6ypnUq7EFfu
9IUU45zl9oles3KhN8I8sM7Xnxvujt2/7Ut1cQJkGRa46EIvE4jP4qaZt1dxen+mCfe072kivWbg
8SUJ7Vj8DbGIfYcS3shj7a2dzl6/qc589n22jMYtzHySeLSu5l+YQaW4AudBH/1J9wiHRAT9tSWn
IGuZ0R2mHdHhgpxSFJSN83ziKu8Zje6pApBJ7A1JMWT7zjf5JrvKemKMiOJ+MQrLVfrnDCQ+pPNi
MSug5y54/8bhUxjrdmij/VkTmkL92rwKqHdHeO1CpRujJZKS5kFDvsjB4pSVT4wbETqjUr0nRVmA
GOqnDZr53eL8W9YWUKY6PedQ8bZueqm0b/BorO9p8Fb2GsZ19i1zdaPERCf4SQqJ0ZNNQMVD2v+T
miZspywOPpD/sr61maqaBEeFDbmMdalZ5sNsfC9LABLo9SRzWc4kAa+7NnVJAgNz0lmO7iY59vLu
iLPEaxIrEXJRophXCVvtD4EiHhWLin2lG4I/WG3tEy7kH8EW0YikAZkP4Iospsl6eiYsg0urq2fT
P9g+IlQExcT+PjipvGF+czgS/9erbtRdoHLOUqWT/jOcnFfnJcjikP4T3xYFxf6ai7jA5FtvvTTd
IcXAY+We5ctPjEqh2tp97BSgM3Li4zoVp5tGlweaJctkLE01+nqfdPqQlBjIP3Eel80nvvHIeF+u
T+NBSGKb8loXnJPti4JRCDZsn+0i02murn9kYVCEgHlS/CnAVOgwuF6qJeiRELtpbg9dlduW1k7B
YHYla9Qu+Pkgnuhg5W+ckTX3DuTmskJrlAYwqkkywXpJCbSBxPw+k11uSiUfzCOB/JYcsrhqWchb
p5bp+0XBQm/Z3FtXzXN7C7n1OeF0unvPlsaq5b53NYFJww6vBzSWwmOxoIGNT2WEGeSkfypOm6Zi
P1oKjKNeZeq3XzsqYvKXBUSRkZG4GffFqJ5LtQvKz4Ij3ZUxukm+Ojs6DUqOD3CESnEmQI5aGIGb
97RgqPWZRHhXH6fp5/E8LZlu346uC5z7nhBi4JLsW8CPLzeduSkWf3lVfW5NO3EB/tTiVmJR12cI
9kVCuw7lRufCOUgAuIWwws1cJiivC1D70DF7BM9R3pj25/ltAH0DF7nJJfuiM6jbZz8J4LRTM5p+
6ZXlx/6IlV6xN6afkTyBoSc7lYw4WyUL1xTuy6wLNFtUgTZHWGmow9Qk7PdSc5AC+2RbI0wdgq6R
F430ckOI41St70Id02EU5/ROyEXxxsvKORUfnFi6kQMXv57x1UCsrcTCdvn/x9CvgAE17q8LOy1j
Ne7H+DtRo1LkV6LYRk5Ig2l0e+jpg398FMauTmsHEZrDUMnhk7TEYH7yV5aPjwl4bzKybwDj2uZq
l1Ohv9pMaZdzg1ceMr7ArURZNyC1bnoXYyXBzn+SzlB9Y2+ARnPwdrLgbiG9LKZ9eT4Ng7gPixKM
X6B2nlP4NGhiJGs76y+bB6QOl0DRrpVUt7j1jSbWDtV8zuylem40ekkgG/N05aVdqTCPQOTuYH0f
Eet2iCSLToZ/vZ1L5H8c0se5dkr4qIxk5ij2Mfl+rjfS4xiJmySMKDhcDqQa/XD/F+Rg9ss4J3yf
cmkRW3qjPbzG3Kn4cah4dWDY7m28OmTGIo0/FUT223ozAcmRGF3ZNdZQDeePUrUYv7kI/YPfPy7A
4qUAUq4RK21WgfGnL9M9B48IN+mXXhMD3rObnFpjbvEs0wUsaG6cJ5yM137dtVn5O/3Lx5Sq53rE
WMeLU8ZY/svVJkWWEY88PV1uqkkHuvRC1v2Oce6davxq6dXOqw1pBWHbxxly9ObL/fpWNhIceTJb
fnVzPPLfM9MlQTwiy4oHSLWCCFwlQ1fyFYuTvFSIgnTqZ7nMeNNxRXxDATWzJa/fAxOr2FwPwcvm
0zjNFfGiM4RHS7UjGymEq3Etge2Zelhk2MMYWZjCxOJyNGcfrAnLr95KiroCZBuDKeU6IuR3MQfT
2pDu0+JIe7afwMrF0ZLtajNiwY3jj66ZMxDg8Mrys/Hk+rrS1TTKagIYcYNSxKwVf6rIKKCjpXmL
jiZmelCOZD0FZNAd+gpFfc9Yg4/FHZJRLv9LnU0Car6Jzj7+JHOv0hCnwZvPYyEVaTuqjnKQACMe
d+UpGcHoke/R0dRBSFIPVoASAa1jhTaYGkej3zUIFOyogNHQtz7ob5Rf37NzC58AzjGS5dvsh/o1
9+3wHYG+dmvtoxRMYZ/6DCJWfsvYq2Pb63oMCtvFSIdOsgLsQP3BH2uWpX32wYJHSxMvqVwLVKkr
uxnADaj4YF/HuPz4q9zoS3IEVr8UJQ8u3XxcUR+opkN02UGycoB6QF3Z2hGuhyAbF3JRha5khsl3
VCiBsUSn7vV0i3eGxhBE87qW7lf6Q1emlyOOmRm9KX8ttZH7wdVcarhwPO2rRW6ir2mz7S9omPLR
sDPsOVGYvx1xAi/Nk9zytUUDUXsSyMhmT+wsMFEmCazxwo/JNUVYzYG+gAw2Z+6joVzSOg/sXCDY
S1o2DQuSOFQoS1W0VCCUAFhoKO0xuwSQYxh5ERIexsXTRO7dQnOLB00QMilAC4+IZU6JteS33e84
5B97wuTzVMmiy7FF+LK1NXno+jl2MR7thr0nBPBu+jVTNkq0l2KuefMo3FbdmQO2PemgPpDwPa3Q
TvuCBJFgsyErEThV4tXuNibZYSoK3lmalV91I1MoX3IetCsdR6ElaHvTKrf/pMCAw1/9eh6mKVQU
zTr9m1O1v7s3paTkrNNeD50qzw5ErzMpIVnJXMvnGz4gWuP1cAGeNX2kRU0F2709w33eL0Jqi6xS
kOY6jDhU2gUbE3JqAygcV+6+qhaqvMKt/1NPjmOt1xEjWNnOMrE6LnbKkMmvpilKu0idCYcjWYAt
8az21T52hdXEHjPwWeEXRn0HECqgW3K8RObIvqfhTg6A7+zeScD8FdExDs5qJC5OFyuP7PqajPRx
j4rqzKFx12GBTKbXuMf5pmL2ya0/w2q5IyBQH7zmHBfK4PDmXFhgWtXcHuVT5gqZ4MCdnArjMxSE
08tsD+6OKjGNnid0u0CNI27x00scWJCN98nnxvETzVmtu8I71KduyxaEIjUT5TFFUbD8fjgVRRzf
+kHN9Y/A7v+gsR1iN9pQhrQVCG1MLdQiRbPxnMsMIhRbDg5jTVZuH5PyU856e0NO4yYHfsKNSvdP
n7UFrBlwPztWdM9H7W0BOk+l4n8qgGSpKrOCoJv3LNoda7qjXfU/uWSx3NQ8QRAsAMZmyXz1Wa6f
uIsdO5t3/pGJyst0KfikASaRFXIGYim+0p3Lfl8DS0GPsW40J3Lgq0EOMD7nIbMIRKvM6Z2kdXC9
xSObUjef/K0MI/Q/3DBmJUTnOk3XMsXmmViycUfJh4kJ22Ee/hqQxWkxv8kRgPrrdSkkHwqhIdBq
XPcJjMH0EMASq5rmZEdWAnMyCRsQzrQKDjpXVInXWIQ83uTuaFpLFZrt/lVRnEMEQjlFf9rLQT/c
FsiNrzY03N1RFpZ8SelPtxPZGW6jJQsrqTJbgvRdhkd9+LTY1fQ4VUX7LYJAzjPCgDInJycdCl1W
0GGpEtpLFTgsFYCIFJhrSwl8MariUiUzL0wA45juCWUCBmbRZsjDKnGzJGBHDxrHJeRrvYV44JAQ
yJKvoY247qry/YzmB5y5yZoOKBDFKbpSHwz4VCXVHoir/gc5wX6SPK5NUPU0wwpFELsGD66HjZy5
QALt0hLIywZFyJm79xGHEbiQZa5Acne+WRtQkJgxkE6o1roYxHTKqm8LVPAu2MnSDZOcZUPtrVhE
1YKdhoBTNDAmqswqfwFV5Sj0rkjw20DcipTbMgWblI+WHCa03sX3kZ/uIQ47Sn9AB2e3h/P0tO6B
y38ktjmLEqkzlaBHgJH6b/f0Go4rCvZ3Gp/KUBPBD6pSoxN2+V5A0RA6ts/RiIKHsPgupdNt9BXZ
kheytBDDmFhyGfJnbeUi34GZnjRnw8x1H+pMd+aVWO8u9491V6FKd0hL1Rakkmt59hYvTNOvgrSq
jyJ1GFvSuWe5KChr3hdjs0Ij0mAUKE9idPO/DCMOOMcHGzGf1Emyz7Klgt5KVgllYrYL7unSDgRc
oF3x3bY1WL7dhR7JfjZnPOAj42vz2b9l4dDOlXXx8nMRADckGDKR0JitZJB2VFs9M91Mduobzkxa
sm6oFBsseT6ucQNab0sCgTIfCusadDTel+xvXCm4r5E8cFSyPhf1N+9aKdd/mC4ilgHXz3tEniuQ
DCNz/0byc96ehuRyppf9FmNjeDeBhtwZgQBQsze03YEUniDNJ6sv9BJmlkbV4cYsY5IaYGc+V7GA
rxo135k1Gu2FBrS/4dW0J6y06e5LoFiEE7sNWMafOZ5WJNDxZZ3q4VJee0LrXWUpWQg2UltkP399
EPoeBvY6Xc3HTw2W1tI6kJskJnurvRGn1jydQtbCdczTzWS0R78LayVw1BUsKumDeF5jLScr/FD1
22klSPN16bSSQGwpeAA3u/q2tLgvXXjJJL+8Fb+z9VTQH/KLqiLQ5kBYaKKU2eelTSkU+5rYmnmo
TQFmnkIF/WaBBhILmAnC3JRIsl6zeZ/rSq38HC7LgKsqkBhChBLA6TgpZme1lZDqZgxolJzDg3iw
OtNzRB3qLMJoYxFi1l15ZayO3H/7+sTjF0jfvOlv/6zT1e0fZ4Uo2KiGRMpObqQPwPfw/LMp+TW7
fJMpBy94MEsrNGKmXNoF8ZhMcPNjYpdjpEu+d8haOIpPwZLVL6D0/Zfihof0KckGeusomy3lg7bB
PCVEXpNhneNQf1UJJb08K3dMyuR5PqF0VNqwDV8u2DvIAUih1guJmha8Y8pDkCndNc3DVwtSBkJB
Tz2PfFdYLAqJKNajgR+DAdQQWuYUCB+UHq17nt0/wAw8eLrR6nRerQCJNeCRc1U+krKb02v4x1Lf
fEG0lff4L3lJLpVdZUoP+bi+q0lKYdCXK8lcO3/tu2bTlDyPhiVCSagLTJa6OsEQeNzEo7EnFg/u
iHDgLo02uCTb5sFAUHuEpvh3fWm5SfRngUJYUjFSBb/OvITeDNSG3RE9aW+81yltLJcELlnMcCpW
FNwakWGsIJLMBRwH94S3/t71F0yB763XDwke97g5CNbKZAkQji4kcGtNdgtC+Wt22pEOGdRQU4F6
d5MoFp6FCYsRDiYVlwyI4e5XLxsecJ3S344A2GhNhgJLugLt0beZbR8OT/kWzX/9xmo0ulDJy64D
oQlbDZONJlIy8YG5f9qCHlQnKO7Vd35mZGfyq1ymvSgJFYD7QvjtfrcvDv7OgT5p/vrI7JuU5gZJ
j1CDgpsmPqaGdqu3/a25R/FyNS5l8rv/Mjq0RUp3hwbP9jn00witu3g4lJvGFdt54r9wlC20Vqx+
F3Z9Er07md5Pn5wKDmRtmmotJxbm7syZNyXzfdF73c0XTph2H8SV5K3pXaKfUFbLlgOnjEwWwF4R
1BPHhrAd0XDJpb7xnaUBB00Wwk1sSAu09dBNBssVCJGm5Q2nKTvjIr+R6yMtSvQwUVkRhILS7vUh
CyIdOe6AJl9LBQXR0plb8Z3DhZwdHksNlZ84l+ED+vqd5VSmGcWQAnisKhRIiaODDkJwwBqRSW15
oLopUS50afAbiN9/tBLs2sBRe5dbXXmFF4laIM0N9WvTs/GyIaijpyIDKMgoYSv0E4ve3lqncFSk
RKr+6Zpf+kz6ffqa+znmwhmuED1DjDmauoAqz47rc1xTFLfdRXc0kNye1lWhdXN6NzG8jvLmgyDm
0HovJvEjYv9brGuMVxxGc8/xWgluAuKWWQwdB66t2CISdtMSkke89QBDGXuPwa5YRc8jXjseMoN+
JsfUAWdcsWdcYukFj1uCE/LB2rRcdfOf12SWOGBMtLR9xJ7fbJ/LpgjoB7KfTP2+c7aLP/Zp/bzE
A2Govy5nTx2NhnbFTwQtMLfbehga5eGZn2auQWxkZNygUIKuj6f9CSwh/K6HPxnxWDu5XouSkZW8
o8bfuX0uGJ2Uc4eODFPnzxQJQdBQSog+RK7rTq4WT2WdbaBww6w0UaVPQvbnRhdl0IVN2Hc+LGJ0
N5pwV5yWE7EILqznSre5op9ses8V+OI0iw7kfM/b/TQJ99+DjS7j6zLZJyzapVZrverqXjohUrF3
cUd3Icu85DiucWurn5sqlEq8zYV1Sn2Pkyp8RUxL1TRUAPtWcGU7Ziib2uqRW3VhjZ5Ug/ZGxAWD
WZNRjW3pkOs1vYaRO45RAT5vErBuq5otYtFTXzhvI00/klsQKzQE3KFMWiRUH388qG/jAnusNpa/
mGCE9/H97kgirdaL9qIZcCd0AScr1QuGS0C4sby09mniJjVzupE/hS6Y37n5Of3i9NDxtlYmREgg
mUKa6pynhWyUKYXY0+a55HaoLkUvixdXfLLI/BL7sa4PXmYSz4ihkR2oKeRQ2zjEXMmd0ycyFuJA
Y66jfLkB3iOzwcxroGe3hrWLTmVc4sVpp7zG8u9pLLTrNEdgQbflbfaZCpQ9ss8uhEyZOnvKliQn
C98SdQTZUaJCXdi38vxKV3SiKc8CFj6CpCePCUS0u2DYKsr+2j7HrDju2PaOeW3JMSv5iYagYyin
fC2gtnvt2AFB1r9E+SdTSa6jxvHWScgaR3OYMD6+OtxcP/pifNAeOXJX5dI7DTWN14ymN8rshW66
9nw1mBX/GQYzlB8zpwJfvhR6XznP48dA95n7LB1cz0HYvFm0iLBvJRuJqbq/5haHnuYC7GiYymmf
qzzO3GnXa6V3TooWoE2uHBUOJ2C1oKwm2e/i6SC54zAu+UCeNPqMmTwRYMclfXC5Or7ne3sXbf8H
cbSU6pYzT4EhU0GWPSU3wskrzC7xzp8Egbj2VcsncFiWEXlK1aClSi8KsT7sXDItCHbfy24oU3Hv
6X6GFYY9OIwHeMkphxPy4Z+SwEJNsf3ILz6LZX+lIubwvdWfVhhCO88EvxpBaTUDt/5KQ2wEdTLi
oAug6WwQ7DuxGNY3xd6TCX5hu3cb63OkgCt5GauJdTRg53RsutHgOD0G1mM61vxc9pjFCMl5VxLJ
3G5UbRlE3DqZTSizskP3IzmUY+OP0B0fomO+817LqJHm0qTubtYAbphXExG+SktY3CEJdL8jJU8s
aQoBk4Rl+rwJSWJCK9TEzCEmBtg9Lkww8eHrzZmFJ4fDmKTf7qqnK6ZFk/xQz9OsUP2W3qGrrz7i
2Zg9rV32D0UWmqVS6MgT3K8NFUsEMBSxbbc6o1u9RXou53mU2YD0pYqE8TGkqMDCqZpv4JCwOUao
167ZNyqGAr6snS5wnPW0hmywKkn4UYmP++MVuLMCgFUS2JYM42/Rc8iWbf4LF13hmExjq5t3QZwg
UbbKSyEdzGnwAlFR7o9qEOt3g+YjOz9Jwo3/FdzxZc6WWZOcPC//7p9B5WzQkoqi5XiKU/vGq3QI
J8F1NA8jZSC/iW/ozHuqDZYZtEC7bHBSiMf5jShBvpVAgjHf9fBiQFfy7oPlycs/zdwiXjaQOHic
JHZ0FhGh6KwqCUHLEKX03dguqMXWuGQoEyKTMcTJdJvG+tyK65oLMDB24KgLigwZaWKjqY72z4Eq
7I1tBiCT9S1TO9RKn+xpWKL8aMB+hNwHfYhE2bebTJ+dsmSMfkB/jlO6PYrbw9Oc3/o7fQ3TANRQ
1Iz1vQJnnp1MoGYDeUv2sjRsST9f2RWiqiDL1/eVAQH/WDFqx4+bKENhUcNYE0HuIo5ePtKd5Oog
kz9LbL/zRWQSrK3KtRDn+8FQWCtHQfGn/QlCKeWqvLY/ym4NZBpPTSiPZTmZh2XJ8/pWgTkl6G6o
fNWqmmDjIATN6nHyxoIVj8saDD04xyFGkQGGdYt3IO5Urx5w559d3YMmMLR0YgzY8Z5mzCCsA74h
YI0+v92G9gM5xxMwGG2iJZYWhI5FgfrA3bcHKAXUvMgNWfyczOwshIjocryybYAFbPDJj1XS7cmY
9njGt2g3+0J6jtoGcnFfyqdWly8VDWJaexcAJNU4x9sPhGYw7cSVYFyEutXbjyM0geC5SgYkrmji
UoR1/hlOXEFBXKlIkfQaw3wJVDivMWXAM6tx4wSFtnjOWLcK6OUpYzXPHnJilW8x76aAoY7KFvNi
1sbK6HoEFkiNwuInAm/jtricESL5zo2moiMPXqS6prN7mdB8CuAuxgQbQMnnXw/MODuvVNKFlHJM
UN7MVOuqqmQboSjrb64lBzs8smr4fE74qgV13Y7eJmsEfuaL/05HpioFHAqM/k/b6nxZwLlEZWQk
tmhIElW6QeB5iGQINeqSwWRwQ5ulaRwaoOGDkaAA3ycd8olvjEx3nIfumJkKE6L03DeMXetrRpz5
4hg8WKDegn/4Rgiic04DvtaD1m8cCX9n90MjlhKbrIQqh76gsGum9udxHteM4Vam9dxAXKTn0ywV
UGvVbiBLRGcVcd8v4dtfM/3GhogMfJhR1E5hbSPBmpEuMgYciK0jceF6oWOPHzsAlz3/aHyM1OO8
b7NJxNbAnaUO5m36Dj7+xdfwVDtVuUnSfqxLqNkW3g2aQV2XSB8UwfCXXESo4OIlL4Xs9hirxeMm
AGPp7AaDkNMurSNkT0CZOCwNxQariGsNzAhwPPupSyEaWWLpp5ukry7NYlZoow0PCWojoxaH+vbr
LMExoe55mVH9ywkIIa+r7bINW04Zmh2Bh54zgYiPS9ZyOBidYJAAmJqXZRUK5Eu3asnH+IncVsFG
A3ANYGzvZ3tUDOcdTqrvZvLY3B7oI+JnK9wPShHfzeJnlXenc1s6KWRh3ZfGX2qgZ1Uz0cGuPxq4
D5PiDDCKyUkddTayAOZezqJj0a/bbzWM/N4Qgwv0qyny6d1OjMdX18YPKZl0xN5F+Z7D5SW1G41Y
V8DJUnbhvjYi9Vr1cxmOitqGGdvvSGV8nhakb9q+fEOXdgE0kpxCqapaYSckye39cezEEfAWNGub
20r9QTvPSI5zgHU+bm9MDsR/TMaorHUgAZ5UzApeWWUPUcaa0wVkR/JDTbSLu606IlNwcgpARX7P
kGOlqIbCtxF/QLjNivPOyYfJig6WRO1Mq8KbIEAO+xvqdZAk2W5yCWF1ZQ6GZaMELSPcOqU359Ht
RrXcasxe4zi+gdJl8BIZyq/iiY6v6d+megYOx58IIKLIV7Sh2oxBzOHAqDvKbmD9iNE5uFYIr9CT
N2aMQvjwfp/kK4tnVyuIIW3mtv6gdTdWZi1Q2kfnq3DsrOAv8FqbKZ1RRptgsr5ykEz2TLSTbYDx
nuq0svEdHaiHYsptMjfHD+LuHzvTW2osdHa/7p3bmmp9c4W+1/p0c0b6PltFTVxLuPwkC7hmWDqr
9mciu/llNfBnc4p4vdSP4KOGeYSL47yu5B7WDYu+bt2Bb33YyWeC+J9KrwbhMrm9CDuDKqrDZH5o
3McHKVmijVmmvpNk3SZfuefoac7WjMnMEDjraha9JR+z/aW9PLC61LWX2DtCjIMmR8FoNSSLyUKn
4l9N9RdoCYfXh28SvVlCNpV3CWIn7HweVDgnlBWGUcdTkvUdJ5M58EVIaRXiX3rcAj2OLksWMGHP
iwMXghW9M9N9ET7OOm0J00mC5cy8V0pJDp3HQJJChNsulbB9hwYQnMWaNLOXxOG4rMf8Rn++lF/k
8gj5aMtnuXdkDZOURlTtQVZYoqPDBF5xSiz+Uin5PcFtHk+jydxlGcUlqO09BhC+TMciz5L4+ktk
OrZLUBt6Aq+9tBDrxokWKk7EquSBIxw/rcCYUwbO3JKg3KVXmxFqctRE1OoCAbhN6ALZU+VHI3GW
s/vMO92F9WzS45aRfzZbUO6quOmmyLtwVF0xLhgVoH5uO3lso38pCf7gsTAyVrrf/Krg8VKa9Fc0
il3mvutzoRU+P05JWSUF15Wy1+KBBpS+GRTtUSy1ThwBOCAXV08Tzg5i4JfnpXETRDsierJAxR8t
zlM7PqyEu4ra4HY271m7/NJIbsJ3bWYNyRhRa6H0UXLmCVrMYK/irSe9VOgl3O3Fe/aYQdxCcdCh
mFwxjjJppgQ425mBXh1ubpAePy8dcYQUaGpjYItkUeZrZcfLqPpQKa/2TDRHqyoNo4a5R0kgzqXv
M5SKAQ7mbU6NxERNXkY9CS6rGDdkc4Vo+5XlGJjts+ocrny2I0VFPZNNrDgVHML+1zIGE6p/Azll
jvcGDFLG1CVHOtwRPpXSJa8IAzNups2SVHqzTDwx9Ql7fAyl/iix+bFpCvyfSlabb0z2kTywesFb
QUoYXTWGmehSPaWhtO8wM/hejoggBOlIpcbnb3GdKJs1Msg//QBI0TOjdgvYubv5o/fMfziHTE2W
lc3EHoQ6jjJk8e5lLPzvq9ls6WBfE9c99IIL08Vy44n6ex/e+CTbhIeT1/915pXoWyM6x4yZ6xWb
3Xd4I+wy14SrdnkLoichdhC1AQTVj7FWyb9XP+4u2rGEo0vrx+9lyiD00wqczOsgib3kd2ylpCj9
VKrMB38QW3xYKR+5XijVU7x9QCoHWZtioRj9My44VQ9d2u+k3dTiepFNsnZTAvXc9PZj41bPSGMY
+SAaaFs/4iSkxz5GXag0+iioQaEmNcme2xwnseMbEC/N2t9+ZdsVGdceJEaz35psMhZsBSRskcN1
8hliaWfb2J+fbJNPPAtRWi+x4lXk5gW8oKQ4AWSzPzl9dRR6G2zWXtW6Lvo3wMljolbwYKmZII+l
3z0z2AH6Zgvp3ELwOtbp231CNlOt2bdEcQ0/dm+jBS1Ymmnh/y4uE8BYPM77NDrI2sXLsvd8yeW5
33nRSKE2oN/+dabJtu3DNbnjYlbphq0WjP/E22iHx1oDb1kx2nP3Ia7TXwiXgeTusjaLj4xycv4B
tbpX80hyCnmlysQuPlyIBzWr6mdtLfU6FZjvix/jqlEUk4iSN61iQH09c7HA8ldU25nj3joIRQ5/
9gsHhHb63mTcFPMxA1AyqaWzam1qOxsWco39vRJHsEtTIXua6j4v5OLzlbfov2V8XdVb16Pu8e2c
KXceSc1K+/rr7O0UvfHqWkqJgfFtjmdTEUnyeAx/kj7uhCt+AqPHpghodonWwRIxal0BhIVw3/yX
hzfT9+lwzaE6eNTFyyk20vYB4ktqWV3MA3UqX+ahWSqUnkSshb6ylcQsyd9QjOFOUu9rfTMaogfb
NqiZk4XWmikTOcuEst8CjgBx68WmWZ+pUdlzTP0FL02qoUNGuYRbwHFb2MtrZhcUE0XSbXLqvSiW
z2yOG/6wVQ8MAJqm3MUJBAf0nhVteiw9/OEziOfAaGxodxFwC3M0OW052Dx4OGEJPvF87pnt9kn3
oP0MdmwO5fX+cusAu6f2Xx2FrLbycB6ErTLy8DHHghS+Moq6csNQ6nEjARbjRZFpYxY2zs8lZH1z
k50e/THd6NIVIYKzM9gWMO2s594EvkTZBkC21urHylHEAVce7CIGtSPEckxV5VPavDpehAKu8lqI
dlScKrDFAYN3canI77JEGjuLDYG+w5JB6qsKHPQFddoGWimqeLIR53g2q02oGNsbPVaJwtjIQdjO
zXH7mmt6e8bsPxrglk4gVVdl/pJ56gkwInLxzOjle9LedrQ6O3lKv0S8hfOICXcoTRhlYPIssXet
VFLmzQr25QlMfrnFde4wZR6CKadNSJq13ynk+sYdGOVmE92thydzxojMyhwUqDv723RukLXbAqIK
swJUsxgOvOCHNfYJElYBgCN2Yj9q4w124ntB3/uDFPPhjaLqMJmf+VKtGIunhBUt8AJ+XsxgywT8
sYgKCdjb+pEZEOO0S6FFjn+XxLhnhUMEyEU9X9cYA/gT+4LkvdqjEH+MjWUvTOGUUSWKl7GXMeIa
JssyN5ZKDzhwLApjfsqHN1sURmWdg3qXXMgUmXVpQ7o5piqMDs/8ozLzCtlQMKN7b4lS/fogvqCb
hO4I5TEQb+lddgUtwOUW1YA2uU34Jb7Ov7uNPkj7xlbmv52xtWsiJFCbxmdScxLR+bepGN5SjTgu
JbHOwIJzPjcV+L4NsSrE+/mWylsvMg2pIyZ4G8DFB8lfQdAP8gm9WnWCUmww+6P9ywBVo45axLM+
H8bAa4i2e4JnORW+vb6x463NX5R8Wv1AEh3rchzi2+mmZQBUHuPCzavxjNYcezdVJzBFRNXXooqN
eOQKBwiYledHQDqxof2jUhiekS/dbEsQQ/zbNxzTuI/UXAdjPS8QHjb/x4nXH6VCSpQ8aoSUMbAp
bAOEPX0wCuPhsRPqtnoNHE67DCmM+6R1WqdweXmFUBM3YLZAct5wpWJyF1idNYJsr6jEow1OYX16
uUEJPNIpR6rNINzmKAUOK8Z+McCY6UOVOW3XP736gq252k3ur+t3V81myxjByvLY8dYu0PWxI2k2
1h35l5hl/I0+3Z/anmut36nL7sKpdYwmkrJRv5cu+8KaSDTWWbT0l24AK+ApQRLKYH1y1AN6i/MJ
237trO2wkXcYdunxjOi69NfcpB4i/eLI8Lea9f7zFAG+QIbJQBg+7m1uDvwhhCzSkMWU/+AbnZD5
j8/jHfohttlZQ8g5uOGzsWirMvDTt1lcfLG+odvhvjFINQibhD3KE+DxQd07zMNbBw89GVAMYc28
asgrv3zodtT8I0HR0tYMa5OSXpNvfSyVMn/x/GFEibIAp2t7e6LGtFuNFGvzZnN2WhYlVyqvsma6
CEn0EOKl8OLVYIdLKnC1xCeA+ZZo4p1hXr7n70q4d/naNtdeFysnuKJUsaZAv/Pty9x6WATERS+t
slNYxyfJaZiW9cISt0mtj2TKMuYqXJLsSDVqjsGrd/iwx+YqeUjnksa9ElGdrb5pDJWobF/fXzvB
l2aRKWiFKcrC5dOYODpCArcTRWKNgb/F1tNN/O7Yg4qbZptQbkv4FMx8vDe+DYNbngaMvFR2aXji
wiAF6bIb7D/RfdOd1ZZIa8lpF0EKbFcTwhCWAVpnJgV0NaNk8t5Ji6/2UiVrT9vCZSh/YfzqQjzl
9CBwYYi2Nlzdo+XpVJWulhoJkSZIaHJ+e15sGkEuv8wzKG9fQlMTU93HYzHIbwmUXPiaLN+s77ej
v3Y/7vtWI5kZSae3sxFYMggv/1nBI3ePt2O1BwnKfwifNxvj8LLuSYwSPlGkOxnWLWvNFMCgDthg
Ay1CAK7SAHrMAxq4MGemmpRzonl/FaOzIULPaR4uN+Ld/P+weqLZHdKZ0+YFyBO7K6dWanEbA/d5
/uCYpjIkVXOI2OPcwY9Wo4K3ukdqQVjyhND7zfoAB1N9vBwYMvJtjR6B63vy4deZXl1NTTPMbEcI
qM9KF9ibKP6/tRVFe0p+MDSdaTtlpEafn4jX4jBKpdcEVxD3AP73D8jQPH03h7SYLJGMSZEcGahh
5duZBdenSOXPELCv75Q0rKVmvuvw5RXC5W2AAELyr7xT/l4bftW+w3p5HqZXDAZgF8BbFVRkEJuO
lZo4MDEjuH9W3tiMhc/pvjTwUJ4SQA1gT+3mLkSP0qtroV20ye1vjUS0U74VK/QIqDbbd7yJnlpl
NcGULJUfSoWvG5WRKNYGVsENE3ntJF1/tJydEPS6jlZRpqthNQhsqQZuItXyARJnzFGqw4ByiAFc
gqKtlIGVL/EkOURABSBRG4lZCrjvwv5iWbBUgCK5DplX1r27xdxtw/md+wY6hxCUe+XsDwX1d/Ep
SX7lW2taPrRYSuqbe9afZUJOefBd5q1JjyC+qt8VziL0I8wFyJ8ATUli1ozdZMcoo+v/ke7a8EY1
UFKoEnUIE9xfVAFaDzbvxFlN2fKh2ZcwEyFM7gKz3oRxhV0W1QS7ngxbasXAy2OcCLcfDTk7oj+F
T3PRjPHVW/UacuQgasWE5fyFIBO9tzgNDobv9AuddT1qt10CsytSAeeldES5AvWuRDxHTulPcMwU
iegPdp4+rAxMWAZa9EBf4yrscoQpaX3PlZwS3RtQWum6ArkZrCOCjfu1SGnJDfgXfN7GoZIqq5eP
pHkIOeTfaGaAth/J2LM1Ez9C5j+ftcMmh4+YrY+grW2JANEeKw57j4WQIxOSRQ8dm4W3/jWkQNC0
H0Nlwvtt2wgN2NTfPSXZDQvxkbvIFQLD5WHaTEgsYHocvQZQmRWWP6tUhkt0yTJlSSoddqBigUQ2
G1O250pqlsQ7KsNH+v3zXPGOYLwNijA7bShkBUXMCVdvfehkNKl6P0Ozh0XAQDJPhBbMQGRg1LdE
YyCyB17irUSmK9t2WzPvT0HxJ1Da8KaGry1yZcJcv+/qAfj+2DEBuGfDM1S/gyMQ2sZSqRku9R/i
A0qZ9CXI7onOR+Ahmnb6kkQEpi8Ybfg1qHSt3Yl7BDCh+KKhL8FkpfNgbI84vFpK1JCbObdvbIK2
Gf26LjgcaFX3WL0kKSyrl6USx0p1zOZMBRorSnQnhyn+orGFZX5n+pxl/oao3thIpe7fxirGnZI+
OdW3puuFovlxCiCo6tOk/KgcnYg3fgj+lu0KLoHwB1qS3g8z8wdjTcF0m8lYaIZ+1taSHTvl3nIV
8z0l0vLgEewpgsRDf7czoZQuECBqiURYuMpfHWp/AENEpQ36HZ7e3LJVH61wdKOjhDxf4pTPklpr
QdLAKhFJ8oldTy7dr6ySkH69bhC8O2yq7gq0GuEZ2oVstsBkmZKU6wQYcK1WsZlEfU0+JPdF7HVr
dmJfKPolPWiGk9JKMJMYwyNZf9SF6Z+F2LlWRhtxMkNF2Ube1LWIlpTvMk2irOuVti/SV0Lq5YjC
tPD2Rq0UshaZTijA+FLCAjofw6XnUQLt81r/SUXWN8ho6VAYCAK8wM9DDCfBCePrSUanltdFADkU
mKGhcOwNyhuXikMXBLw7+0D9AQ4IulcSAFXQR+KxRwTln3paIIs83yJ6NvoK1KFg/2EwEap2rwNB
I2qM0FueanxeTpvrMt0B42A96WuxlT6ljQlAgGuyIy8kUELw9+0839ESnMPw9h1giZsjV+itOamr
Y6BX/VFhwUEJs9yf+buCu1yKqGZRJWr/0p30JQHqRyvcwlFWVUn12CAWi2Iy15ZsLEf4iKxZEte6
TWASgBdYikLmFPWj94gLM49MpM9gu+2d7ciQGXMoQLa/4RnWTKDhTbHPrK/kHRqQfIPUXX4Coz58
uqz1y2sQfAhW2SAXrCLt2mfoXN9kG4LWa6tCAtaAwSEQYS0dTFNwaCLIHq1b8fPBYwA4FFhlhnUn
3j1qiFgYc4m/7z5ePd9JPjoz3HVmIux1aSqfEnaZh3fI/XhUpLjWAXiysAVswDq5dwo2Bqhz5PF0
ZmT1U5QqYH915KqV53P1ZyA0NvM+iXj+q5CBAfWcHaBhhKGywoQOxkRKmD6GXW4yEQGT7/SdFX+9
lPOmtTecbngBHB2Ha6MAMKNmdMkqY7B24yFJzEy0JU6uq+n/kqftaMAdVWIqA36P9aRUYZO7dQlW
0S1MnkTWwCuuD9NgG328RbtFAbpAI+4Jky1Wqana20gA35W2y13/kyIn4M+T0DT2KmzpfQ/L4zSj
8jo3E0ykvzgvyQGjJSJrk1VAlTntBE017AJmfjdVLjbTPLwZS0gbPrWBrG3O/KQwNuYh2iwBQ9F1
Ij+pmGIsQoO4h1w7PRZaYDKRz28xi2Ptd2N1y3b4OWfjm2R1Vy7LBKU1CxZ53doM6pk/eyGPlIaX
DAjlndlQtmNLym8y9v3KpwGG8wOhRNAH+7pzQii5Tmm+tOR1i6oTHhV8mNRIYy3EGwW8Ez5nzJDc
byArSjbbs/m/wWPYwIQHt0Lo6dnMq5i5f7Vi6Qhpnacf2IW4ho09PTp/7flrDPHAfezK/73I638d
9Hd/S5NfUzbRoSiQBNav/NbkWasYawlkwFVJpHSqvsKLHm/nWvu3UCA/CjO1Or7G9NK3NhtGpgi3
9IuoyU6YQhpYJllkRr8WrVbOGcjk7abrfD12cW0rlsaogPMhxLIybJOr6fD+YPuUuSMTiVpZnD+g
9ECCjFlWrIKu/yAHkFc/bOUd+KenC377kOSN1z64sC2f38f8Im7LtCeKZiEfSRxb+9fkzYjqC98j
CrqtlvZLvDrNIvM06OiA97TOfyktyj9JSL1laOaLEiWB38F8raB+PdLEdwPllmQVU+OFxnLtjFhL
S8VQzqKY7d3aDWRC0tglNH8CqhedvU6WDvcRPTkJ0hRXHZVrfAG/YZUK8bpFtBViumMvVMo/KKvI
dHQXMr6XjhOLNVjJE8eVJiA+ciPgDnX+h8rhgu23rAVZ1skSCcbzAy3jXv+4wJpqw5X/E9YA/oKi
aaXIWu6bbvkOO+K5GxO+olAq68MSEYnpJhzLCbcwEg2LlW10FuWjcoj3EVaiWCS8RSbkGkxd39VF
4pnOw2hQLSmynXF/E0ErY5iU53vtjXiPLvFfDHYkv0uBlZRGjMOKORWtX3IcGa9g9tFehXQ/8D0J
aMBM4/Hw4FXMEhZNwKZ7/YgE9kz4U+Gb1zyf5YhAWK4E/IdsegLPIDKeSHiaeYhlffmTh+XhMC58
w8cKhfmRV6IVWJbGN2Lhhh8EBqjclanZcL/9A3MVYAetyDZS5F4oRXgH2Oj1Y17rFGXyyFc+ko4m
k1N+pAk6Q/BKnHVxxY8nr51TF4kJoOEV+uDNHACOdfogrTwOEhM7RXMR2dCz54dfZ/2FwhZFs9bq
SKdCkMoXqirWfEQ9yWJPlAGpH00xWaY6W7cHuDsz8+Iewxp7+iGRbMynFI2UJRPpBJ/qa65uNfrc
2ymLVyMPz8o5d+jlUIwKnSEdGNjJysqoESJmrZJ/MVp8hOYWxtO5CHEgFqGFXxZL4jFGR7sh+4LQ
xS1gnhOYESHcyaUSlgLzTW903TgerDYcIwace1eaa6ctldDLcmGz7vxkGSNfFBwbB7hY/GD71IUV
SQYJA3xk6y1sz8am7PEWsJmrJ34Bs+ek851eRNvpEvAhVYMDeFdCSnm6DRE3jjC5OdRp3n3fL8L4
lUMLtdJ34MmtVG74UP1cTFYAWE1S/Sh7NJBMFw6vgtNGPfgGfdTg5Mv949kj4ScKP/xoqTrepyRH
UWzwn56rFwoQ3CrHFrQ2wqQayRut10/lmI2E6AiXIxIL1+70Go3bD72ECDoJgVuUr99urp6yn/QC
+GBcDvRfraXxJshkYkigIQkSNe2CwvwxZ9sFV06jLyTa0xmo9ctATvkYbVSuE2cEFHZILwXaldOD
lWxznC15wTACQ/UzyJc2YEhnMt1LgKbQDjxNPAETyAGg5TEX7QFCw98QV8bIg3HlOCGdulFCGTA7
sEXpmKBvxsP8gFV9gpMZr13q6NakI8N6wZSZhjcOrJqW3d9TSiMYo8aS1QFK/s3eYfiZvk60vJlG
6+OQyb00G786gJkTXZlfUgikVDTPHRDkcO+cP5kUVZ9yLlDWBFIS4HSBOX5qws++Cjh4d4L1LTcW
KbDy1ekVRpW2Jzrq6QrDxe1+MX1ME+ce1nzYTE+xURunzdVPd4W/f+Qwsvi1gPufarLKXeFCXG+E
Rp3jImP2YdEM+NnBIaqGOi2nRi2IykpZvVz3MaQxPmW1GTqae1FWsORzQF9ireMAJdynRO7HAo01
yZpa+YtsOJ3VHL2v5nIygVOAZoA91mwusmxTMmcMURD+PrKWALm/GJgRanblEs8d4s/dWG4S2BuE
52oPKgEls97aNvii8rY/7YpgOgXWTVxSxM6bM1k2b/GHJUaCHMJcTlelC4mFu2gUbjELWaD/nsPn
S1KEuAcFnF6zIwTgiTFlvzrJb1rnoS7eYr+NZGKLx2we+pabwgtcLJUq3xakmGmMJ48ij6VEkOB/
jvSwQV8rkzRWrS7/J6VcxQkG5hc/DPwdUPBaO8BK9z+MbTEmfPTIgha6mq7TlskGNKRdXCdAG3Vr
jwOKPgYPS486teK9jPgh82ZuxIU4w7JO/pgygMJDrQjODfMY/ySC1VRIvhyk7eV6KjzLt5XfNNBJ
NWNAyqsenezU30etGMm01HtuOwZmJX/Y8IHBuaBs7vq5WJfhkwL+mOl1jh4uhcy3GfUjzeAs3YRC
RzCpUYdL/k/yjAPfuZbUKujDKhG8AxMMJFDXOAmhtQhjNaf63rjrNLmgsRZVwAyIoZGLl4l+0QXJ
6emNp+O6vrjHkkvlgeNt/lT3NQjN/C6IX/tITKNJ/eQrVJ93+yZ1f39l8PeT4UEjFJhMcF43JqRU
+kYNglz/phgGu61pkwCe1fPSiJ3XNQiUhe2ykdb/1ZfmRIPfydvILE23n3lNdjz23If6VwbdXLyQ
0C51AjFvVVwERWs6ntt2Bp1H29bV/CknB9Mt6T8ejkPtAd90dLqlsEGYw02eTykHcNTNS/kXEreC
HatyBmlDga5ixVTNPVY/7WmDGrQPKEyX+a4g1/ZptX8upPlzhFLbe1Yv374/gUCz30bg/Vjvn3eu
nQpVywQ64UvvzQ+FX1jHdjDvCz31TiderZfARDHERgnSsjIbm/dOvV6HC9aJqgpNl+AWzBSks6Wy
6YSdR/phwJViIeZ8mJuwnBMV5JKy+vX151JsjUsOEjY6Ro3EyDRMP/Hg8hah2syvmpn3dmPudSc7
HK8mx4H3a9W//pm38aNVlnP52QUkgaD345VfsSSXCcZIOUWVDh7AJmg3iiQPDsbvOWkPzQmEspYe
jJwP1THEtcjPh9nEMvpMqdyj6JlZcA47LbvJfjl7UnhHh/EzhI/eDmcGYYQLvZiOxf13Jo45biaR
vyGHICYSOGb73362CbIEhIkeLnIABgda772nWBGD0tfp/Eu8oCZQR5pbDrBJP8ZcH7FQHKe39lX6
nEvDxRcA+E1Ey3DiTRdCDn46kc2CPyNWCHVD9fk6Y8j6Tc798GOIY1KvaeZAsTQcwFDqtngAJ5s6
80TKV8LdCkFopw5A0+JmupTyDnltOihRcZt5tUJzidYJ559VlXgcfpFMTp28La9hs7qyyWtFWEzP
+Fcu78Ex35M3Hi6r9/6LW1EdziGex4TpQ6VJ8g56iPXOBuqDKoHBD2XOdej8iLG6jCKAU35xnURT
fQuFZUflQSK+8gY8Lakq7xIb0SCNdsZFeNqbcOJ4OFmGIlFhT8bZm601hvKf2EuY/r9sZoQ6fP+q
2VmYtNcAqjr4w52cnnLZV3LsfZFs/lFimQOyKVL2lk2xGrAM1/bNXu0wDAw8ZjMlSOwCYH9GT/GF
MJWhYiP1BT7SFTMUR+a4Tbnl4WBM9UnSnbfYZ84GdySTEb4oyGd9srTScCqpZq3Hfz+PLq7W6ckR
cBulZQz+B7Xiu7whSdb/yCUFJkpj7l+ClizkNTW2sqIvD0l3/NSF4MBKMkT+KOiasm5zjbGTk/JZ
F8n5UFn5cG5XJ3yt8wdD42IcJ9sQDmt8N0cCFLYS8F3FUGX+bUXrqTy0f13qiGHSF39UU+2PBeeb
UVwdG2kdolEW5bPfCQjq8CE/t5I2L4/99SWOHa9aXbxyI9xQjkCYul5pV7okLqMVhnx25FskTByj
Fkpy8+5EHgqbruqlZq0+eaVq7bfwsNPlGwdKo4zHYEg/lBw80j730jFDsxqyWJqzElZh7kqyCKfA
+nysKz3e3hf3JD5Clk/w8xCQOe+3u3JYfosB0aQL6QtsOJNeZFgbpZ86B1BYtx/Efon8B39sCXmN
rtlC8OeW+lhVA7Z5yL10C6s0zKkdREjUESylbyy7uRxK/ggM9s9HYdg8sGmyhS7aaVINYUNLdohF
DxDqgZOgEazM4c4s3moBYbW+r/kT2uS8nhWHo5wVgsDsM/2FBHoKDNLArngxB9CQ5ksJwWQz2BB/
Y9W5foOF9bs8EI7Q+i6yqgbgs7WB1fEIdgGVDt8hRho/LEaDGLo+BGT1Le9tTvyhzn6eM1cXw4Ue
cooOGQ+P0bDYYjff171xTfIy2wVP6qc/EOlZ0o8i2/16iDbD5pzrEdmfjr+mFZYF5TIzKCZsWiA+
7W9wVbMH2vTH+uzKiboxqiwvAUHhAJ5Jl6q3RoWluRgSEUrlze273u00V6SeCr3YHpqRsWKsbAMx
QQxWGrCB6GISN4eI4hx1G9dgZjTgH83HbAoI5qA9GH1PZyXVU66rUTCm9MbwaN70lNcvWFDLkLph
bePqQFALO8ILB+C03mYodsSeMEa1OCPSIrs9hQSQkjobRqZzoRkLRhg5TBu165PHcHWdnSgfAFIb
CMzSR9I8xRUGSlKmVN32dSNmq3IgASRZMumCEdiEMAfj5XRjas7atlZ0i3/TVVQPzXIFqmwX94rI
a9IWEjl+jCFqsNC8bM6y2MiwkDhR+TIWzDrk9B7DDoHrh0K5Hpsj0oCEDbn9ODyHVU+sEK+ZuQqD
xehWAcg9Q8ckEItQAev2EZI+FRwxYLzBTnGS7qjdu072RAzAR8auFujnpwlzztRepwjRy4pZ9bLG
X2RvC+FcuIFyKgYXXCGTGfok0ZcSivymfQgqtR5iDosibhOdjTEYKAsRmJOHG63FOqLQDtAZ+ZWW
Uh8oRagMVhcNHuMJLZFvQC/s/PglSusEtusaU28ZUplIS882h58UuisUXad7rLsE4G361XeGZugh
VvhcF+flvGUb84DxgU9bHOTHqsag7g+LZ6bWzjgAr7uxXAIc4rCn9QMKl2RFAgNgUpmrbsEZhvCS
PFNqxjax0CI/mTR+EliWFapQ52NUJO9bxfpJHNIO3jxvQQYE2cX/TX+czOk6D/odb2mOwThhYs2X
XQwFnVNrK91iCRMj50/neny4EUYG3KRNzpFHQYLN8Kqpfu2JYW171X9RdIc7utTC8j4O7w8SSZzd
uIDXyv7qgqivwaJOj4pPjbYzH+Spime/6liyymMBte+WXu7wkOjLoHh2pAAaW+Q6wXmHDsIwL8Au
P4/JmMd13g3/o4E9f+44pPojlswQZAFz54slTEg4g/orh6U+/ZQCTm5pTdjndDHfEiMx8DxtpBGU
dZ4QVsiK+UzOAa3uN8sDnraYqzVcgwTcVGdKwQXaIp8ocGFV7pLUV2Mn/C6f0+w6ZibhVCfKcCLM
XyBfKOrOFXH3KtGQwn4FwYB4QTIm4NRfGYqFismni65W3/POOw0d4zSLdtprqdTh5RINAY+FBycv
E4jQLuB0pvjRTFjwVS6o3x9MvJqxxc6fDxv3IivUj7XLDW2a4RvjG14yNmAx0FV/hQPvZObKiht2
qZPDIa/VEhkq3N3IZ+D1S9gRZODUOtEHw1iwfJSEb/yej873ulok/wMK/otez5Z3u1Zhlur2ol7u
1GzqPIn77SLEWZIMtz8yU6ZfOQUaL138DfT/qsTcYo6BqvQ5Mx+QZI4L5IgnV7FffhQuw6cDvisf
BXAau+oKWprmr8w/fC6BTpqf2o+4mS4TzCMFx74rP/Xw7BLHPTfv7zr2BPKsVbuTnKUF/srnslti
zD4gPyg5XFE5QTlVZGJxpmS3l+gvi3dwv4Pozzl/Ddfx5MUcWG3VbpdUuTiFQvnElVyNmODPKZC5
2rUVr8I6Yi7VmHFUGZGQ6WPcnmBp1eUaflTfU4u6TWvLVinYruTRvw4F7nJ76nFyLFkSxOSd3imX
EXkIc0kOCzYDfM2SFRzg5wwKh/Js2fCuNBm6QP3KxG5AqQUpu9OPEc1S+TDt1P1bESvOkOkEA0S/
WAgajiEN0uMi0GGAUDksJdev+XUiu1YkYV4re74RsnkfeKegiFK87MfJ/dwzoPuY4W/juDDMSdaY
dnDgQbqKfSu/dBUeFwqWtACO2sz78JaJi2XfmAErvbywn1P/sJluJeIjNYmYAd35reCwn5WXBaQX
pt6kx0ezC6t6QnDVrVY7DJQofd1pWaEngICd071G3Iz6wuYPpDYFcFncjruYVXpOYKSMdN8vPjtN
WbA2fFQ55zUD/LVjzCAcNBHyEZty65NyDm1sxsbNHMKOO2lln9AA2chCJLx+zlYtb7UYBumDmw1o
WKsaNp4xbERpBEGt5YQD6ehn0GJmM4pQmwpFtqR2pGFsPe4wqMCZzqmxPuD+FUJZTyQG53F4DDHv
SOv3wRJgOoL/rWshJ9NDNA3fBB5SKWEc1S6X6NXLHuzl/Y676Pj5PRH0YHvlnhSN34KBcGR5WnVI
rGbmCAC4PxloVw+YTWE+pn7AyHg2Q6Q4iSIDAHMDuSpyh+bLcmEQ50JwbLkKIa0IYBrXgV5DTVIY
URgIWuf1NotMwt9pHeIcVClgfuEERuhobYNo9Cg4CBbyfseQ4XJ6KjAuWpTpQtZazGGICbiz8LmA
266nD/zF1FMjbpxY3Pt61fvI2UBUmoYniIwaRlz3c9D1pQC9A0GiarjIWUlahQCp0+P//2/kD2C9
MrW7+63pMjKgByqEQ3wdp90Zn2DOsxqftEQ3K3C5AzAb/ynfLqB3rLrFCYR8x4QrunWF3WYNUa1I
zZzPhuolDJ1+CbaOe/yjDJDYkdYUH0hCNAFTkX6ymDQStynaftmSD/5m5NeGDCm3q2YXJgiFtv3h
JZkWId42wtua0yEe/9Cf3A97BeEd3YqjRkMkz88GZUaxCFPQhingMcB1frY3kES/KfrRL087sS9Y
iCkPlwioNl3HQ/icTfHGZ4jpuqX007rG6ao7zkNvMcW3/B2APFLQt+u2HMMSbGYrxI5dva9un9A5
bQAMVfPbqw8ow8urw9R10nRlDNiXpY28ZeNr6zeqfdUWRE8wxvsHEL+F3ONEVg1te8ACQpRCMTeP
1BbvYVv+DGJEYp8+zaWnctHrjzxy39hPpSKconJtA6xF/aoJyw/N/rXA6IcbMCn4vqN7pqTGVof8
OTJSH6v7s9foy85oaasvQN2ijdLVHBuznh9UCgfo/Vybsqvik6cncDF05IO7ZU2bHvRPZ0pllSef
4iiYb3YWXa28gRnDhTjZYah0qifR4k3FREHPSfrWaJZf0o7EXzq7HrQmIFrwuxMqNOUveNPcxkwT
r3UmwLyfGJJ/r5g5J6MiCwFpLpAagpN2CIRxXJdc7yRZ7WNC48KgusFfUdTwXlQmKtx2XDpKd2lV
ChmNJtjnJEMVSIXl67bVj417t/RYPS6mCAUECK+Z4oedR1dIL0Stp2jlhsFv8U/ZKZDnpT49B6IX
2SQsUi51HpArIbjLJGEk36Lj9fj3Y4iyLF3XqgWiqeXeTtBdDRBgluSOXzZ+SkugBjJP5b47HVrZ
JTYB8IHYLaxKUcKUMAf8wkPmffRwqshK6f/ju27bLSdzYTyoB1uz3mkoz/i+1hgebZI+fJbxnLjM
HHMCUjI3RkLb6cWuXfmajap+z7XvumZ81Ir8xHv4HSamrEDad+VnE7e8jpGlbn0wxkOeJXaFgy3S
7PkRNrb+tcWfTcnKVcG+Mzl+f3fbSiD5Kjb3z8o/1qqdZw5MLvjWSVW+XW7vkImaQalCyGPe8Dr6
sUM3FlhIuItvgw8VUfRm1G+zTgJJtDSMMxG6iMXl/JqByhmNaikL67r2eP08WeN+FDELuF8eg4cH
EBotaECJp5CoDtMx/Hy8Aweiunxy9zs3YrCi3yJgjvBxLgG5s+772wqEiqyjuX92BujNGysUgtuO
xLzDR4f4d+g8J3V35LcsZZElohn7P4yX63uf3PzcAudTJu2t1fzYnSiZY8Tg5bHJK+uzFhPctE7V
4a6E85lFz4TmobvlBNvOllQNOsVU1oNwh1GSY6iuk6FHJYYrXjldfb76c/IZhSwO42EkiidbG6O5
7J4shc9cXXtk7PfJ9WdUprSlz/pPAcdKReMJJY9Qz3v3LkiVqERUax0UDLe7J+TlmjvdckO7KQ07
YR+EBx+WBn47lUl1AMyXC2zMh8Gscrs+HZf06Ry0ItuDqEJ23MCPOrRJDI2e1hcqx8OZr3YWorgy
569qVx3hfTNhdzwdWpXUlD01JIzWAJStNXr7P8p7TbPNUb701rTbwnN9OI8fge8SCxx+F/fkERQ0
a4RUmnpUW1tCcStz/xqnQuQ2FGZaxcdwstM8gNmpoTADxo1mlkLzJhV2xuHVjNhDhuQjhY063sJt
DHfcbdALSXdmkl0JrIVlgo7FTLV6ZH9mMoGWD/96ks0myAav+qNBH+zQ9pVZE0J4Tk0VeKYr29uY
3B6omzLFtkBez6gXucxiWdYV+8798TqY2OgsK/5AXAzBuC3LF2MsLKRAa5kucTXpKVGLALGibnQj
WC8+cLGqDK5L74iAWu6n0cHmVRVmpNCC9HYL0ccpAuc3UOHDS86Zz7nY6XuUNaK4fWWojw5QZ+Z4
olngiUfx9VHPzK9uELx9me+SQikPlvrBFL2djI4i4rqx4MVY3yLmQEKv7c9gGnAUiRjICaM28fM9
b50fxnVwcIAN31bHiNHjDTFUm7LXmlN3H4sDDNpsQR55D6pQApq8/pOnECwHYhciFGOpQk6jPLQ0
FZogF0TlYyWg3Ktvkkb55JyRgJWGBRiJPjeTQjNWDhhIdaDXukdFPwfJ6x9Sp+DvRS2qYegJx5sT
lFgAV3ygPDNjyAFHkjgOVkyFATtiTrz1XvndyqwiUfLOBPNGiJUq2WWRxvpSTc5B7yWNZoL9Tv/V
sOeJm78Fvf7iLnNe2nEj+2D70SAe164eMjCZ8d/VJWVtHS7aHsyNjIOacNJaAzPQlwdqy4lLenRO
bFtFEsleY/OD5iC6y0KnRBcnokDbQHz9J9SRhRY/O6NquTgIv656yJASs7vd4qFF9ZSRqxZAET06
Rcnp8PY/2BLJ8gGcUSfxIj5g9FUdKg+q9NdjeES0flGuVB1V9LEEZzLdygIMwPY7/2hJxSOrcAoC
1t4zL17HKjOlq6VVYJPv6Pqi9x+UA/xVNVpgHpl6ThWiIIttjFPhjnfTTPRh0o2Qnqx4dGxUqtQF
w6tOCJZFmsfXoToP68F6vPA7W8RdWJ7B9bc4ptJ0mqAkUd7smyhommtoqJnpVEEtDSZ/fSmWMWVH
EprAXI+RtiLyRLwC4lbIkUO52fApG5YMKxjZgbXwaRTIYOPjYIhwzj9yKG7iE3RR5J1DwLEP1+y2
0k3d5tQ+YmOn91p0/iV3ybEWTlONFoG8JZ1XqraOl1lC13xsPHnFUyfLtHbNw7C6DmZVS759b7Vp
4WHL+nVWFLloNe/BdDztOKAAfzQWym/mP7skJb/qgO6oCtx9shcs8gtnpgTAbm6gEj+jkot05Jb9
aVxtv1mATDgPtTWnh7JT1TGfJR8kpnyHK6I5qIE4CxOZuWT7IoE7pQnb2JdQzA+6gihNzAkIIO5z
a29p8/TS0S+NkxttyaOwYID9Xp4xYcx/x0X/X0Sp9LrFofNjHQZoC3otekecF5gF5v0IMKcnDxFq
SO7G2BmB6gp8t6Du4ZzkCHs6fd70cqq/XrdzodQZ9c27zSKSYwLvUIFIXyYg50y6ON+vWVjWK2My
TKFDFLkogyQGl5ELpQLb55nEBBkf5MhvyC+jVx4ZyXzxba1xmHQ4Pj+IoFtwlwaAIlK9ruUBfEvu
VdmV3kriFjkeF5hVivvyqJ/WfsqrzYZzFlMGLOhrJAllkERgWHIVPn4oxwSnW9zHL8FgMwZ0VOQ4
kEjsQ6aWk6TUk0nOM+BuZ3C6scgM2RgY/krDrUuRphYEqCkgKmZmN+qERqaCGTqjjSovJ8e4xY+4
vNoEECYSBinHH6SS7ZWfFqZKPNqsO7GO89dSehjoAoxt1rM+M5XUmX8oi67YrKkoabmmuYKDOD1U
SSCUn8aUF52FS0lSa4aM1HZoc4ktL5xdcw/0KrOiYnmYm/QW5iJqAagD8/wgiqykCnhGwi7CJ9XB
FfSJS/trxbuAAglLTMlMdKX0R0PZ8HVtksRC9srST07Rb2R1Z23kpCmlzLqX3vHROZ/f0D86a4ai
cf66J3DXUNV4+mewfm9Y4WmBj80wYeJpF+OnBxl9gZAv8RbmuGYr8lPJZehmAvHpv8id4Sr3ntog
u7cuEkqtggSeSwJk7wIT+NBEugTk/B2XbwAL4DE4nVURKro0mHWWix1wReenaLoAqOKG1W4Lt7c/
EEdoCqAA/r+tLs6/Jaf8P4nWgrYLjtFDW1SLPc2T+4rGrcxWOEuILZBFAId/LLY1ZsK0K1J8T+fu
VTJ+B5tRWsTxghXQpndcftSExuPiBvqUYriJdHajzkMutsmyGAF5qPcQ069a2Q9xtXkYN8ecSua9
FUjCl8fBHVMa4isObtdWEE9aFJ4Vh4McMJhhqi/2sLtb8++xYaujjKDMrbuKX+MnizJoxVz/xsgy
I8wO1znSXWUoG/2pr85CR51Am4oxlc1LkGIUYzVi5TUKJfUm11kEHEDo4cOAEt+Ma1+UlVvyz075
+zqcBI0RaX1A12u3F4RKum0XGrsNDXKKD1gGlSxwQ/cdE+4eIppbkQLO+d484QBiM2fzqQxeZ1Bx
undZ/fcHGpnnO7aYAcBXYfp2zocTQJ8LnxNwx/8Gk0F5Lk6bZp26RN/IrQb9zZKzs7vHeD5203Hv
mzXSxhYbH7oVoQY0vR1H0Vh2OQ9GEMYCZIw1yU9FpTSsMYHTLW0k9cpsgs5/x6m+0f3mWcPD/oYp
WkOOAmrhK/jTrSl80XqqElkGMocaxxiZtKSzZp2SyDBBAwRKk1LZ7fshIQzQUefydBksnkteu59i
0RQsWYQw1bF9tL3WI9e3jyx4QEQOj7hYdoqrPeX2x10Jews1yM55HBJsL9VB76kFsgNCPUnKq0nM
Hy4zL5RMPlpqmk0Tq2cxJJkvAObiqsE/iadWbRi266LVjloAzcEbG080TE7vdChVRNDkKgdVq0vu
2of6PVPB+jm1//JVGmbF0hzjzfFvfDKBjGQvsr7O8SYkO53vya3BVzy/gdNnN0UMN8gxwUzi2CiR
xiTNXNgsJ5tsk84o7EGzFo1MatJBx0OlGCj9TlKRuWqr2qWGLadagUdY7NZ/qoA8t5SRx55W9OYc
ZI5cWcieSW8mVaEQQbWXs9GRWlrn+4yaeCYvXVYkuKPdVFWnF+RE7Hwc3/zA+4TacDcL6kxfKgqA
3AnNoRE2i08ZQgpVS9IK4Cv9UtrXR1UTtGjYj2JprmXVVVbM6/6B7xwU4IewbKXFfDaQ9My2YSQ2
zzDpOu3/ToKLGyrnmOg0a2Q+rj/3ylqm5DBrblkQV6oYxVR1jD0ICbukRy6p92asny94QZvlrAzB
lQUzs4/Ki5OYbbPfFpEH3vUzKJn6mx+rOK8hRTfbm10rck9mMHyGlbt4Ukf1+bX+/DDrudUzz/sg
fULP9tq65SoKhKgAZMK5pDvPQUKRmNx1UuPgM25TcQwTdCIiR0DGMm9Al95IJTxe8prh+6SzVj++
+MSlJEI0rTwXdpGn3lDGQXEWpRreddPpbIxXt8eXyyWx7Igmdy6CEqzzam9ebErTZxzOjz6mz9MO
gLzf9cg8jsyyQNnYhEj7f/Y0MRy6hjT2wpL/f5ifDA0ODVRw4dW1v6SL4JBQoHoJeCX8iNycA/gr
okprfDaG7Csthmwpi4nUOqZinW7lYJHMqPPCqy5vL6biq+XKsoQ+fqZlMBu6FKCbaLQS2nth8dwM
8b5yqG4QxZ8AayZJW3vHhW/1tSx6DRsJFGtCm9NQaKmn0jsuiqZ901EkLw0iQvzNOsCBSNakRak7
mOihCiSu3oyIFn0eGGAVc+VNCfCqb99HVs5FzBi3x+skXnC01V6VCHVxazR7319E1GdjmLRG/2b2
rgg8aMILuxICevnFE6yMa+VCHesVpuJSQgXZCkGR0633Mw6Mm3t4A4E/ucAKvU3kj965VGP67Y/0
EOXHgr8qdJd34OfFqBafSGOZ65TwQGf7Vacgbl+SLRK7w+VyJ4mYzDSwRzXPSvMsBq/ydJoY/HUx
tP//6ZD6wP3jZV2qeEI94ax4WyJtfJx3Aro2BCCYbyBf82WJXy3NUMXZk98/QucOrD9SBlG7p+G9
6/3UJrOCpoRcCGs2ToBr5JOjvCfnNF+VaOYm+maf5XIuh7NBbQdfCt6A9fJYHxvQzChqlnTDahnx
X1Xrt/dV5IE1JXC1juAqtNy2sJ/ELy2H0SE3DAjR+yh17B2Y786pAQC8KuLKQvFMk9033dc9recl
deEdz2iSN6qWasCrtNsyG7v2wNzb4oZEy7OWX1n+xi/+/zlzUPI4fN3EgGrQmjVf7Tr6x1c93i5j
0C0l8lW1OV2GLOQQpaaf9e/pWDqTprCmK/s+lZBU8oPUT4kdGO0rgZafdzxiJG5KzRKek5QRB1pV
Ur8vujt4IYR16xCNyt8iUyN33SHWVfQISJJIb93CzoZ9pWi3++0YtLH4UdodM0WHjKvl9QSIKMe9
+FjZknpwS9Fe1TCn0KpEc/+aD1ghBm+Ytj6O9PMIvh39E70HcEtLBiCqfGj+PYEK6bhcDOB2fxA/
nm6rzTb5OHHs8/BZJIZyYmef1aMrwJBbX3yCMVeQiW07DdFE6XND6Jc+6JUkrpAUtVdlBJnl1/eW
kv3EFpEOycUmlbL5/oDiN3R+i55MYT7kTjAQzc/cVllbNyC1T216xGcrls8Pzbjk4xw3/wzFBe8k
6oyd7b1DzZXkA70JsIigPdW/8LTB/hjQs68OdXhNaVudd3WyFPKQOD4Ru4xNf9b6BTRvxfplWO+6
UyKQyvPpV1r/zz3YOLRHn1louVNRffdbto32KDz9ZS/YAxMVgNiIhVJuygooiQMkeTM5Ohcf3C/Z
3MyIg39h+u19H0529gcdvWiF9eO9B5yAANfr1AT6QzG4Kr78+Gv/BRraElgn6CUSFIfH1hejY/r8
gCtwWWSn1VWKrSE+4qedJz7UrHenmMxPFNlfTm9vQdHJqH1vHlLr0NNZgb7vyp0hnjsSGrHMcj4J
2UW/gUtMNHqAkVIKhvw4B9O70qTyJnLgdDAtfOcPvti5b0c8JuCF8JytlOOE2PA9K3PF6FS8+h8B
ctwTQzTJdRaaDwVAoCpi7bzRKc3RKxBdZtJ3Sl90OprSCLqAqsWfDT7Rt1cfgGCBhvGzvb8Lz3eZ
x+lPVebJZNxFy1KLp2cNxWOrwJNTqvq/UheUw3h5fnEDcHIgfEmYl/lQAZ6SAEeOTbb2Pg9X1tVT
dP/pFUNWECuoUtu/35kCTb7TG+m5CENugjV/54CMe20Dfmp0GaH+1CPsjGqrDjoHjr4bSzdiXIV0
0VtORAhCxyr25sGc72n1VaYOZFAlTHXm/d2G72pSL3Gfuf0XextkDhTVPLurIvZLh7AwSsYEV/jR
s1IVMj1JZlAnRa5g5Y9VAoDOPT0+ZN3TOD91VOYKnblPcyyylkBelocRSK5eKVqoUPEJ1Gkm/WfM
+v7ddSbRJgY0703ey+POb6TGx8qUasYDIxNm61O2+YLHkBpdmY4WYWedGA/5yT0AlGHpBDcWL1bn
sHyijpCS60zr/pm3fBnIl5IQ6cEjytJLm/oV38QdrXv3S3y7VXmPqtO8Z9/mxfGvnVo2e4f6p/KU
FqkfMffwZhwFECWwkrLwRl0XRbJkEz++EWOh7thEEaFv0AsEGtIAAOA04sgIBGNSBQGWynf1oKAy
JHvZ8TI0UGqRZg4/3B0FzIEwk7lUZ1d8i0DbGcPXLbcJovp785ydY8cojBwg+C9eLCC9KLgVTHqS
t4t8q6j6cyHJhxaEbKvtb8kDvyJzbvPeeXaFjNgV9nw8yw1FVekg2q0dBTbnZwmYwiUwnXhIbM7U
VAZSshoZyUEyOarNlv5zy37bkfFV6IWlpGvJ1+9pRBqZz+Hm6EGL8B9+qV2wXqTdxJofgao0Qh/M
HYUYfYVIbRgANHnMLGLq09cZDrc4KaTBN8SYoeJx4t/Z80e5Wd2HI51+BODIqgppBzVEPnTi65w2
KfGC0gt0RSEyW3+qaaILKgkE4D0ZBppCJtbfOLWids/3AAaT6z4iCtCIE7f1LE85SKqZlnjT4ugv
v05hwes7RrnUWetoCwW9UEGu61N5PCLICHzbuF+UosCX6HuyIMRZe/eTnxPSUiPcTim6trstwdFe
kEGCfhgoCVnRonCYUmMkJTH+w4rWsj/QlqRV1o83BpfYr/v2GH9Ood9lj45AQTiJ+jSvRzOj07VR
th5tYqqhNv3sEMqpzLc/TE+O0RJG2ofBoWtl7R7k1H29rjPPSoXhPVAjgsKwyjh0dUSqIhlYYrt1
uoImQm0SSwHDEWjqVvI2KMwPJmLl0xRpWJfmh99NSF7J1nlY0KzPZTxD/eDT2B+JsNlUXfJMmSwH
2rALUnbm7x+uxEGz7rpoOW+0/AQGoPy4ZBSKqWDod7+R/A7CyxsNH8iIbNOcKx3Dwzb2t/OKxONT
H8Eo04AiX0WwfCtm+C7D/LCQcvugGtxUKq4vvQ5fAgPEUVMH1OsZ8EROJfVauOk/+C15iJP3xVNL
b9/Abm7QUkG0hpc4WIJx6Kl0s0oGaqJxd37q9RexRpeepGmWzB1hJAz9KKDjbYVn934DjSs8EG1X
I84P336vOYt1AIkKm5Wy8/6G8waT4+LuDiCv7VFHRQNTXHakvCSWmrm0UOht6v0p64QEahf3oYPV
oYx1lGUTRchV/8brhYUSNA3ALWyHfSxYXJ2TUvUo1KdoN55KQYTRAY1GKUmXeSdKv2gKaXpsqS2o
Z6FO9yoI22NS+6WLT2H9KcSqHI78lTCSY+YFMY9y1am8E3XdA3wmOWRuFyLxkD4alLfZgihFvpTl
rj00ZainGDXAU0rvlTiyzMiVG8VJPvyE836Sk2MfVrJI/ncVoz9VV7gIqjYrLt7nUZGBgbAmaIfe
IL9T80ka9622KxWJ+emOPCIMHlUGAZe+SKDhXbWoJKELp8sGrV9WQIsdNCa7wl/XfE8FfjeuX5hj
9fIVAuQom3ZxAbdTwVl8DYWhefFoNz7fTG9r+e8OM2aJc+aiX0QV7KnFSWUj88++hAHm+ZYig5aP
kIfobZP5Fl0BQK8UPxDB/2SMz/JXhGLZOVYLeX+pKUgEDjwxx3pduBJhqeqpkdi3A0mSKydwceIs
oy55BzNxHZrsEj/55PQaGZFo/FGXkDuiLU/zOmGC/4HVqh0IW9jFp+Ta+xGqsDYDQw6w+vM2NAfH
dD97vKKngUyKZ+qdf/h+UR2oy0IzS8KIUo1GYkyRJVZgHKjN7JZAMfaooeXcZkvp2VWC2vUuT4CT
2PVjJNRMtGjFz1l13r83cxjVFgLQ+/HYpgF6qJQeuYro0w+n25X0dqzFd3HzEqTJjBwdaHHLv/eY
XNBrH1QAiE1LaJOlEEhJEW2zPwjv6qnudi+3IaJuKf/KllYEbTMWafHoLNUKi5Gwr1sOq3poyh9g
Lq4/exl7aM7jDTQBH7pVV+MH05syJOtziPrZqD3RZZiTu8ijaNdvwljyhom3CQ/9II6TKV/LPy7B
DMCSrUyqbxlEYDjMmpEP/vbQ8cCcr4CIhDzBOes5txIsssWsTTO8r2KQR7BvV7lhgysuLawvFAQz
WES7KSndzn0g8Pl2NO9WuP014FQgk2AjqFpmTui2kicEpGzyk+EyVLHl3ZwpbkBpTeoIDq2T3oyL
MCEaESPEfRU/akQpCSxDHK0Amm4poHT8LUhEoJBZ8mnqfOR1XRwaRNisWXpRBgTypMY1YWibgX1D
mUCiNBidKYgBUe15iIKOpcKeiUQRquqZV/4dnlRoakGAtVXCttx39+1rD1Cj/Fq+qrh3BGqtu5OT
eh2SLvt4WDodc9mJbqq2anyrsRbW3KfinXbMymGd03yWQHA+fmxV5cNrFJwYdTi/KUQCZ5A3Bvnt
XdgvsitUkCnAO4uMNyAEuh6B+F2oAX2F+Wz5/mKND07+iQpjqS517k91YgSd8CMNhNFN451J2CYK
tyO67gVCYJ3MepeAPysGmmj4gsdD5HXx9DzfDagIU2kweyuNKvctQ8FB6UzEJ6BYOGLNqvll2OhT
+kSjq9GG0biwPAfzP/MOBmbHtJLMd3VYhTl8gvfIgF2rW8cQiFGlWhhMEIeOvcmCDFaVGV0aAR47
NdCw7ahd6WEr7700G/QQmjIcqk3lSUfy7j4+1y6ZV6Peby0cL4qhaz7u90O1/nggP/bo7uhGsYBO
UrsG9RgZHYH5NpK9zd2pX9cG+DgW34UcR5xSWlGpAdnicZC4dfiCsv3gvCxil78RR/ANx7nY2Eve
ikK4izOQtbsBzoej8avwPtxwbdU8DTCeY3ZfNKFc7xSHSR+ONiRPLxQkN/E+Dn4tvayu3It4wuTe
Zo0BevB90f9+4CAiaKCs/QVTaLIqpxeRIeSQ0luyBmtFNurXf2aZgWhoikmyIqJIWla8DrYPiiuF
Mfrn1hZCbH7aP75qaPEfY6vzTaC2Rnw1pjoofxONgTEOKUyS1E8SWp5lpkJaaPYVOosxsSh71yeC
PDJ83By1iXbtKSB245TNdVSMahu8KEKW4GASZo4+1/TBTlFctPcvCpKxvk86oLJmWsIyVaS9dx/j
hCcdkj4Crr23/Qq4zv+hqYjSM+eA8pYKwEY3RaVbUkdXToPjAm/iIhGph+IwimUIVhFkcRHUumUU
Wxq4UsB0mR3ePsPd3rn6sYSOiH4egATa62gvSuzgmuF8WL+apWRQ1ggOSpsy4gbjxld/MNWGZKvQ
haSSWLhNsTxAXRhNSgXihqgPZRzi9adMvECKPuLi2AjJVhA01nLb/fVqoexEqx26SRC51FaKKIAS
k/Y6pqraErrm8GzIyJbA1edJ+5vSVf73CJpD+6xIKFf7jnQDZmLySVlKo84TCrU0KBzHA9xHCFzY
R7EC6fdvlHf0BJuVVmb41AJTQWpolzSyCRLbnuVoKcVLPE0RKbIAlZXpPEnBPmtpPr4EqHUDiV+0
UtKrPZzgZjg4MzTrcWap2sgRmQDpNN2pndC/KeEOx8sUjQY6FaNrZXu6yPFLB8HULq9HP7+yr7px
DmYdUV1f1wYKUrdH2qDFBBgXsffleUsq8iB93LXoJgN6wvB4kZIvJttg2J+voqrkg05x/Qej0Cdl
T4/HNFTWRx4q813VL6/oBRrMKFAcBbpt2XpSw6xZRQ/8ORKh7LWTP3O2WHKVX8fUQBKVMQbVP+7b
6rR5pn3N8a725ntoY4OSfxt8VYrDkJhDwKWw/RqHiAv6UiENMwPZVlK9q3C/6NXBs55hyyUlPgV4
yqKhl/diUSGaiOvX185X9GS7AhgUU/83zZMLYy37fy4RaVD5ah8V+uXNY3SxfnQhIZZpAY599XYK
dIwdnidTlHv9o6QLRTvy+GQkNW/7WtVJtoomvHtEZBYhduAzfbn3GqDAx/zHav1m2odLVb/LJIJL
6E19jARZQTTSjvewTcDPFWDd/aguP/gNixmpXy0V3g0TmLtMlleKlM5Dc7/s5PD8yMMWPPzeNKXd
fhl3GgM7WN99ETSLsFPvQ6ekTY+964VoXp3WmezZUgecvmZTfd1S/cdeAUVBaFAZdUQM6Xe0Ony7
ZWodOYnM76kUrZcfmt7lczRuNpdRuS/pkqfMFmZoj1Wfkcl60RZTk6eC9+wWvhPX5Tw/CWlYcr8A
gfGRw75O66nmp1JTvcORs8YBz/psR3OlX3bNCFWdCWOGvgdXZVrL6AZXErN/qXQeMa/9dsuoKfpT
1fsrOTtw0CPfeenmeD04oonmsWAKr+fkx8sR75TEQxvWJlIkxghOJqcFIAtnZ1oyAmWOJGdNmzeU
W/0PBcgZhHWixxLTI5js/fOHv7B4mzGokk5aAnvXnOKinYcZcKXKrNA9bipFmKwOVDCzFYGYorE7
Od3+BJ3JNh2u9jnm0CvmmcmOKbuzzrjRyJQ9PcGCfZYk/Z51AvTe1yEN4zJ+M8gTSA4oi7fk5eCM
zGeDbGakS6APeFa4pHqoVJIQbLTYi0+DsGJPwJUsvvw65f/s50qVf466IGhS0nDMaAYLYDrPwUva
TEPfGG7bBKyzeOXxgHvRxoJrwCYax8/p9i0whIqc1DKxQMqpcQencHGutEnHb7SnsCoF/RzIc4ZU
HsFwM9Z/GreRSoeTNW7Rk1wxIg37K5yzFkXSIMKsRqibAC7TKuxw07eXuSeIKuthKSiOPXfRkpsm
tGp2zC3aN4QTtwQQp+SqYbgdqTimxfpn9XGrxbQ4X2N+18LtmwMXp5gxb8z5lOlTFBC/a6dUggse
HsQhlAQlcI9zMxl56OniksN3/NlXZzDmGrxq++su7eVa4Jsj5T9elM7YusfwtDuuL4vXcsblbh1T
+g0okdpVNbjKllpilOyczqMhTeqoPjwEgSFbGAmnE0zYqR6rfLSrXYsnfOtYgMuUIMGdeMhtlwb7
Rq+m1CfSWYNCKBCV/Ze9hNlbY+P37xOMvcr2vKLXI5F71IF7f78XcHlRyekc74iA2KoHT0NMDy74
0bO+yb+w0Tq9jhIkknb/tSkXZ1gaeJ1xmZr/7hwOg3zQViR87SlEGUH46niNa/aol8h7UF9/ys6E
I7WaQ/W0huKMO+jfrsTgYKd4Kl5neuQenX1Mft/W6suCqRXbeSCTx4bcBMOncdYRCWMziazWhUxt
MIzdMCep2YcwqwPTCWzx/01HlM+X14XnTuOu9GCNbO3KnR8a+yTgDk46BvmxSuQOTQIegy7G2RQb
qnFvwv73mznyxVfRzJj1YxAUqDutUVsdeHk0EPrFRx2P0mO522eA8ZI7n8r85YCTwqWbs7Kg3qIt
uCueaV2EtVW+2JvorFtGohf6QQ+2jR7PEbht94jrtgzu0szxnxmlGZmr9BDY2ue/NfadsQMVVG3o
/8aK72NS8TnwhfokAVJ06wbfCfBA84FfTSHR9FkSXmvQy4n5ccXxLljb/Po4Yd/LMX8ctPRaS62h
QrqNbM0nlfe83zZZQ0qZ98+VhiefaINEwh0CfPwUaTQ0bKYjZC2ZfTI1z2IMNVI1/Uzjag4qNj22
gUvnRkSsqq/j57M8efwk3pgP01nzBgUc1u2N2gcLHO+XxI3hVUNcGHZqY30pi5YlRa6mjAcoBvRi
TCNTGNU5LDK9n/KML34vLUquZ+9yELFLWG+77/T7um/nlH3ejWC4CjJQdKAoUxwZ1LUFwvJGfvoe
Mhqd3d3GO/GWNKNeGtvb2nAzc1jf7LdMu0hj0mXxfoKbmwA88/l4IB79ynh4prWm8B2bHT0mFBxX
oEcD7fZzwHb/QgzajXU4gZT206W54CLBAc6Ji/WTU0rnCx0/5M/VNcuuREDF+q1GDfMHB4wQh5Wd
1bG/v36DbBgQQZV+mLXB5xy38A0/jbi3mizGGnAep28RFdj4Qa23I+XXQ0457ZdBMcRtLUoAChLo
U6A+ZaP4fssl6Ufgn5uRaicSnwCFLhApRLuG/PYEqD7WIqffj6DK3bMZa3HEHblFr4CbeKUyb+Sc
0BG2Ni7oa6eihgUyYQUeDn63e9oB38azp5rsxU3anmUqYYOo/VT40rCzSdabsP7vflphR/vrBr/z
76gKmYwE1FMsVoav8SIM9ouhliw4IwU6YnhbhWcc+J4s1CyrHAePUNoxcRYL09jiqrNTm1GocGDv
Hx7ugR0j+H+TYfBAu8hW0xJ1LDH+KOutmNWhU1pM/oie4EVstD/Yt7sZAKM+VN/i69K/ipnQFPtJ
pUyJr3BAlVen582JWJcWNWLnWNHP1vy2WVC7H1zGCAz/eJgugOzVa8ZYA1XVTjApboYFUmIPaakH
QSFMtl5J1JNIJis5Pfh2C8VMQh9/lxXdIUefmnt0xVrGZjzzBxVZDD/rJjUu0sqS7UhUbXdknvCV
pqCMLb09dgtMPVTs8uoU1ze6XzewGuEry5h54f5U+R9X0+byJoFuSIq3fwoMoVpu2lOrvMIx2ocR
1ehGVZ6XNbacQrPzuHL1uMCZVNDUr456CHAKDl8AKwWr37T/LLj6OQjoGS5jGtKoEWOBxjeKZXh9
YHj9q5JXmGQohqoe6v42ub7j9UKdL1x3fN2rgkZAAbR8GiorPo3616+IxQrg2IaNGjnWmwp3XHJa
P6IEauab9J5YR9REFDJi3fH2pnE+fRk7GKOlwq94Gv+j3++tcLwe60lucfvYd7WT+yV8B9uH3vn9
p9btnqw+iCniO5bSOmtMNCPePBK0cv4u7yPqqqsEk+CNWqKtCf8FzH0Ae8L0gfxH2Aszwx6/tj2t
jQIvFq/Vwv7oEBD+GhVazax6l4euTS27k7FQTpaIO6lWKsCi46tbaL5o1k7b8iZ4OUPahALxngdz
z/V+ynvsRS63c2L2KcGR9AUGSz3G71KFrD31F6v22zQoio2l+MEohRk/1QGsGgv4MRfwxtr/lU54
GZPUSLBTR3aRwIrjAUIJpoZxjk/ErXn10gnmGxMHlaKl6F2WLg3puDgVStzsSDbQvxsa+DlCOmO7
2glXLREXQo18L6MFweyPFPkzwO4aorteuiUkjdLMtZmzSLEOhLdnODC6lQEemSS/qwW9MaL3yhoS
i6EARcaEJJsCNH/6qkG716AE8lQBnhrFOSOLvBOxAdKnEqzFRxHc56wMvsFuCcUzAdR0FvXnziWi
HeadGC87Qv1TjHpksss8hdNPR7yvG7ReiSjCqzgjdUmhNIjmQ60nWmgsSUqRXIu9Ux392q51Oulg
ZxL3vTnWEcP0Tptejp6gHLOdw+24z8LCxTZ6GOE43J4zOzOV0akkiH1qi98oOZb0nHAttc6Ske1l
Ll0eBOhFnuL/GsqtXgpfUqxkt+EFWaPtSriDCMTElmO0SbnOJKzXvVUG2AVnNSmf+alayrDsrqXq
/C/EchkMpFhSdZzevq0dcfwZuaf9xFWvx0ANx96TVfw0OaURX49o77ZjZOXwMH+hOsH36lLBUXWU
M50T0rtUjD6bCpHD8tP+o1F2/TFATIdMpc70gBR7Ti5jewdDGFl9ggBf0tncIH9EqAWxcbA385CT
6e1ByetD0bi3gftvy80JhRUnlKok2bMQSAl7ft5oOXdIS4i17I+AVd3B7H57X3dHHlrEZoqkFVGg
nog8+hDJgBRk8OYjp9H3TLIHJREbix07mPFU7fsRRdxe7nHajD34pDJGjEG0ZUzRwUJK19EZC0X1
4CtBboKe1FGVoRl8PRvmQBr6G+t3OesUx/iYRsm3ZKB6Mw+wliyzSKDofQPrazRCG9286zWBB9Ee
Lzgp9Tj30Y9wlWjr49jLmkjoLQ4dmGCaI/gC7EXbZSQcHLJ5ygmZop975fOLnFuDcXloRzR4NXWM
9m66/Z0Kd54utqYGhHs4ckDwYlZXprnzTl2208Sqm06TOerGjICtQYG1N58ctVKzj1UYdaLtnlBZ
94o4/wZuhsO8jxFc2yQGRdj52ZYjZa44tSVb1POSguMzYFtUOvuFwLiHP2vhaaonJ3WmE94dPJsV
/6h/YdesLuf8pXZyL1UCrCTTWH6RqNQW95YbQNm7zxn3F3b7VjPGQ37IQqTo26I1cwfo1Rmqe6/b
BEqLfBnBKsRb49CWVgi6LF7xEAJJ5JtZL4gCq0EcJKSow1abyVeY6fTFyUzzVh/Rpm/CnuDbFgae
+H/hISTrXsGZ/h64yxc5a4fKR9rr4cekqiAXrQtfkWNMnoKIwZQYIJ3eA47l+dXDe25q8w4bnuu7
kZiF1sz3nost25iQZcuwKoeQvVrVhHZ/OXFwdir7TDAeiQOTeQislK6A3L2maQWlMhHt3MV8amHJ
DBW3EiYR9Rz77nhTvthYkedF7DmoN65qGcpIm+vYTq+u/0TXhOLlu6awd3uJWPkk9XcYosz2+1ou
4ip7ImUG18B6a3KkQBlpl+INXVitKlGTM1lqqaDzSJH69+IVLr2q0gYRT5M3ScFknqEiXRuhQP2T
KjuFthnnkmagf/kDMBxRw/DygyBXk4UgNJ/2oeusDnK7aVNHKwKxQ9hQkTqCgORgqJyGmfCjNcxx
VsjyCpMsie8wTo55fXvFdHajoIdH8dzDnkjf8En61bqwq0Uk15ZTj1+9Ru3y0kT1Ic5XAN3LRT3Q
k8oxhcHZaGen7qLmLOOFvYdGK/Y2WYlX0o/ol96yYu+rz7axhwJs9rEoXO9TjkE+Z/vhTQeVODR1
b9SLsY4n2qYM024blAQYA3jObjBccka9IT5o5Qvmp60PEBhCLadqrZg3Ftn3YW4ke9gV3Y7cT1RX
FPsWmMWJ3SIUVnjcAtg47Cc+xhsCqMKtEqqjlhNa215TcoWGDXaAw12X1GGha1zICZuyk72+kEiS
4Za/3O+yM36AQMgeBgZQ6Fejzs1mw4BL5ubp4YZAdt1Rygfxi8LhkOAnQnJwIbY82mF+K0G7o7Z8
NxvfHD78Vq8zhCu+SOtf+bGcOj1//tJbxFJxal+bieXA/gUVowwNLiZIzMtPfYCxWEh7iklvCRl3
k7uE3W6KAnE9pE++bhmqkevEVYEF+jt7ABxX8BcPHb4nxsvm4n4/O//lrXlaRubD5g4WYp7i6XhK
Mvb2J93rx3H5PRgjP75LznKcvYC5L9hSpI2c0kb5XSKzwCYkpBiVdt8tPQ8TiZwJZliD40RQaycY
7M8fkl9Cy3ANYizDZoEttV+igzgHRbMpfaN6NZ7+BO6Lf6DVP2e2k/9XjazPhPhvCYwoqCySmkpF
fN2eP+/JwcsIJy7dxi7W0tI8LanQQf17YrZOlUG3sI64a3Rq9LbCqBxoopo1ppDaxbVsI3T9Ztkf
7Mh5su1mutnI/4djzivSDwid1Qt3e7ox3GY55raVv1hQxtXsizckl5oPsLdJjOUu83kr/JS+ODVp
w4CihI7oRglCPX9vGShqYpCjCTaArr+BuICQm/2KxaK24JWN8yafA9HXufIxWWZ5TCiZGSNa4glu
N+uiapbsFe/KPXXi3OwAyK32dbPzADzaGQhG1X5FDfyzrlDidN22P2CyZ96nnIj0dfZ3Z74Ct5v5
TTE1vi4CIpESxjlH12rmWkfeAQuRvgajeqPyZq8hqCy5atLYJB1e3W2X2OUQPu4aJ9l/0rFNv8x7
8s8KwD3hPKmFK0LFvEFDlY5rKHngeRHih4yqqRMUQc6NbDT3H81e56FcS4lHtdL76zt5yLcGcl2h
cmB9r2KMSkDXk6L0Kv0L5B7JR2wrYqW+qGpyMtcABrcA9QeZAOLaARntHSaL08S42GZ70qcpWirY
zgTOWS/D3ovzkw+rX5h+gVTXRkDb6EIa+bXkcnlgK6Lr8QoaVJ0P1xNpWXnFt29/aowrW6f1jVej
AvA2EgngWQOvGB+mJQVCTMCxouVXf2KCG8Q2n56NLKV+Bjqeww/6tr4uK2asjZGwfw6YwFV7mYhj
+nsn7ogBfe0Du9f92JuB2H3wQdP70IJ0mc7s+BPkFQcYnzm0o1Ojz6zS7uSp9umtgkRIZorxexJ2
l1E0oNqQzlNI/dZuMvOjjaUiEevrO4mCJ8mD1TL/gHzD6Rvv1VU0ePut91EnzYf86xh5VlLLS9m7
OTQf6IbgIr3o7PwOV6AO9p5kHjAKwlo5YgvA+l8DE6DIwVEiU/dpM8Idt2H7WPFsx91T5QLdzSJ1
NiR1tQIc4DuUCVxtmNRmXJhEc5bQ9vqo8uTkpR8wrNwG1SPbUvIqu6r/XORQrqunREW6asaRe+tC
SQbs1ajwIm1flbFmwEKos4y2pQdZ9jkrroGIi8spC1xbTD3qkvValOsUDYNS0plDtjp6BV6AU77Q
exUcOScrNogqtaYLgFO/fWjDD6ZlUGqMVjhdckR3KBk5qYWUk65kAyrDwrH4Za6/g7Xjhsvf4GEL
+ux9puHuLneXxfobfAdR6l2Zxk1quCvgyPp2TfBRZBWHRk2/q5evinLlXsO+gdC8itii4kvPxj30
EB/gSvvGyAXhZ+B+Na3ZWTRmfwXOuqVzptLW8cfGBK5TWN1o/F26sImyGGwrSJEkqTB+ma4wgS1g
62jfFUBJPicHadENmYFl18Bjy9ZUU0Wt1QJeOKC2QiIEtTkJIVAY68X+BebsunANjbOeHkOGFgbC
zuhxeNUQmXZcH0Pjg7vNQIDcNdBmffBrueVl0jTCVWns+REx5Q5RNhvHAmGs33H2+7xYUXN5QY74
sHAdwj9dlMyYvT05Q081PQEy1Mm8E/y/OfIwDyCOqrC3OISmYBT57SPRv14rrtHUBx9cwi+4a0kY
x5F9AESB33CIwgebzqhY7BruKGCd1nYimiBnuzFuKEIHZFC6tLuVgU3gKP+Ijw8aZRpDzYwk1iUT
T94VvW4RLcwx6RAQoRFeSj4/cofwUanbhTF2jWiHJHMc/Pw9EEVNZZb/elxKkTSG1qTgNsr6/LpJ
93tEdgCulqfGGkVltg2Ry4ZygZ3UBS7X0Xq6VdAt12gMclyhsCMSMb4/i4nCvjVlDV3ouNUlwRbw
zGxGuIRA3p0vz2EkTv//GDoIR5ZvcOx/EJ6WM92+/9MRS0oWCXvlKLKFwqOH9+KYEA6ZHw4JG793
SZkdJCBcgFoMbNF2GsmR+7Q6+kZXuxgnp3Wd37jzSJSB9imm9WpT2Y7RKWpxV4HJyvnbu1ADG9o1
GMVzfGRhuQgqEiiAoYZ0xZ0PrjgCFo0Rcuvej8oGvSZFEIHMkO5UHoWQ7cdjgThvG73jmG4EF+6+
yWqehj4JJt6OizUaJ08Rq1lIORziRQgYljlUm91XFyKP/qGTmVOoDv9CN9qW86aP50Z306edYx3t
KAXFWJtg04+U62vSqS5wiKTj+5bMYy2Yzr8tcDLcsaTTcFMzWuBfUb9KR5UhWXMXusjr+d/KgTqL
6y8yMaxbvPJ5bAvVp1orXBHRwXbLhh9tWTWHkvGwlANqN8tcqus4Z2rOdoSld9OCl5HKg43L0aRY
TSgjwCvKzn4ri1fatxlsf8El62WZ/d4KyYvwBtTe63o3yvvIQipgTUMakrjbv5HHpekcDSkrYj1f
8jOPGN1iEk52vSUZeES7hgO5igOI4DFXa8M8VYqnzkm4pQtFaDIsKIwUXLvAiII6H1L8gwHhINX2
ruFjraBs+j6QRlJFd6ONi+ziZhjlUK04Us4LKfdbVLSzM9nFr4ZHNNBgJ9VwVDuE/+SpcppG3fKQ
kEOZB8MaKhZh9AYC1+Qp3/PjyaATXYl0gVg67OGyK3ymi7WwnX9kZlVCU2i95bWDnYdOg+cyFWkZ
7ZPghQ6nKIgrp0Obg7rR89jH+u3inVGHuv13a9nwDWv/bdXiMnbxbkevlzszWnzXaccAh5rK6WIY
THNT21DZ9+bFp9UPPZyKddVckYMNpe1IQcZre5s+vQ0fzM97uY1zK7wCzlfO1aNlof5BHx9BXYS0
K7OM8NourGOyNTzEHTRUYQxa6G5fh93Ib/q3ha4tPZFhZTlsovXsGU6BlwabL8ITqIkoMRF+83eC
jvbQMCX48eMklylWKyEREsrGpOEkg2rQ0rFJ0fOdbxN9I96e23XVu45gn2oLugCddvl1Q1q6eqDK
W+GDAeoTd+4KILvDNpnaZKtj3d100PkVUu3VM037NUPJahjs2NaKFktYqV51jiP56kupVdJGgyRJ
XvP2JYMZxnVfkb7v04RD+FU88HwFMKfBFLpp2hKe12z1iBCTHsQVl7eEROPwEUEWVs6SNlXSWHxA
wFOvgqaOTxaISoUfgOg1mQ/632fx9jRvNIOgRCBhS2bvaKVrV4gWtSG9yACFOX8UGrSXJl4vdbs1
XDAy17nJ7I1Gh3adniTwq9sg4jywlG7bEah56CPqc2rXPZYjVnou09A+BNdcoJ6rGMf59XaerUub
nAGpxrll3zv6/sVkN6b995eNydsT3C6U/SAApYec7O0B5eU0NJb0Ve0midwwtNtRFyAUbS5Gv/EE
Lg/TJzoHn3DfUwWRJ5v7QoAQPPbcZIg6wREQaMfZ1CQm89apljxiL8N7s2kidkLG5gSusjgGKg59
1uQGZoSOZ3pWO8AU/Pt+cXinJx7wPweQ3GCUm5x7Pcp6Dc3EN2CnmuEigmKCrsrko/qdodnYK+S6
CWVRsQI5e6EsFWYsLH8TrSjpkAuzGrfBTTXyPuK0JcTzym9GQl0iF6mRLVHteJ88ia+4ekUQCbZE
E/1fiNV5zFpRK0gEhYtgMqi1pZvsst244XhVPkLOWtZzH3VHkXNRgpOR5z5ZSPXPdh2WNqrrT6HI
Tw2dOBw43oHraGJ/WSVR66ZHEMnIGlmrAomOr7CPqCnepz33hVTnaQr30g0Nd//4WNcmhu8KWGuP
6HcwEfolqG8JAUGR1+ZQjFHWnzojuSpDPPc0dlSQXqYHkP4qsNbzGpMNHaFEP8fg2BQkqquT0c8q
XspOhlwQm8ITcZEBJSjqkRS8HKnR+7qfUJa2R7YxfUmmJBZuI7RuGrj5Zhks2O9G+9Hm//Vo5qoP
KGyBSnBxKtODBaxCnCGTHTi59vua4O068jKhqnae6CkNhskpvYGeOfULEeayyAyL5rcaML3fEQHO
MOPjgIkfWdXy4PV2BVT55nK7A7WxhiE9QbP+ZJ4X+EknBHmx1SraWaLeVFcjdxlraxDpChSZY+LL
AQwurWzmjetE7B6pj5WrWoQ41wDJqEa9IeblaKxO6EqSIgXbjm4NSSvAFaI03LiDlW8Yr7BSMPy4
ENS03znqiSQIrUapp41qsReL9A4KUE7WncagROyuxy57l8hbv3o5Peu6wp1J/X7ngndKzeze37NK
881CEIoBueMfACoxCzhCfpFLf+Z9Rxk/emF5ThP30EqlXgXx5WmnbFaCbfE5P2PgZdnWTfbarqBK
LkECasAvjKccXId1B5hfqBtBmaxSJID2wdWw/XGKqT/bbEV5e8fCy3Qxqi/BZ6hwla9RxRXkq3qg
rQ+sKjtr26BoDUZ4QglyBEfmfSBMJgsnQRkF10B0VFjJY8N8BZt1EQmM9cuIq0cuf83RFVU9Bc41
qGOc/vXz/gjrnzYWF0No27I/tZ5ivy1bvQ1Ypf4vhbHuopobphsAMu9cJzkoSBTgAtz0WhZOZxis
Fpp0Spha6M/vUep9KBUtaaDVp2hmDKpIjGj5+1olMcPZy3h8C76rfEDFdUOq35lXrgeYtoTNhhov
8m1mx58gS9w3fUP37JUe0yOSuMpRtg9DQti8jcs0EtLNMaz6uK5Kmaya9Zf3hdW6mmKQZDW7qkXL
+/MVg3SsOBpXKr7AhnssnhdAs2E1v/el050l5PIrbI5+C4NAptimWWHHEXz5Ojw9QXCbtf0xNLew
aBTdo9RMOevqBGmpBcieJmTQyGH412u/7zQP/YpQuH00LdVo3gwtLKxzkodOCfshPJJX9gK0zAQQ
3mYFRtu8FF6LXtZmVuTbxapI0GCTDgdy2k+Yil5ZgfHyp6RtosPl9lCTlJZ/eJF7YUZf3k0IyeXc
KvCkkvWXksR3Zr/NEjs8VTtDgiJdxAErrBSYPca+5d9siOCA6u+9+hgqazTgKjsq7VbwjXMLH2QP
Fzr16OMOf0TriFTew9siK4bF8UI8Es8cyih9ec72AmtnjIlSDIjIFbuEs55IRHAH+5E7JhqlgNwL
BLTfIBWEnNYJs7NgTv6Qvv2BbpHdO/4TvrpPnO2A/hZFAIUQjMSci2CjdiRm6uUFB+VTQJrROoQ2
qyG2rwzsmTmRrWkaEv2UewYHZ/N2xjYu6PACzTiIf2p/qODg2PAlklysR6KGBbkwrnD3J4Q2mYk7
Yp/O1d8OOTG41P/k1ySrKdw0braIUSzXJlLty8Tb4qAt2QPQiGxCtsfGMzEz//0jx5nAvb/kgIEL
P7uXUD2aIt+eH6L4XgMGGYFD2ORryyEFjMkFjoE1vDDUhBbFYDUsqcAZYJHAXz6bP14Mw22BCE4T
7E7xTB/F7qBui+vmwQO5Ikp79gznIpdIhq1Szm+URGXRKndAlNmxaDT+AdW24Z/GT66AXJE4is9G
BpN0EabsTJ/EOiRFCnjWcCFPJlZKG9tofvkkawEzGBw9a55dSQV6H7bQVkn8IfmS34DKpRcsmI7R
3sZPeQVbl+wD3DOSpTiqUADjreRBrdBAaXsGz0D9tVAla9pB5TKRmcZg+w+dRbCQ+gxtIRGOXdvJ
kcy4I2dxTf7xJfJIVFLHf4Ist9qgXCipzc32BLFhLme/NoYcgrBRgWwHKLGEaEOlXrfAjy5gR3Kh
o5XEDy5QV7B4I78//ayLZjEH43sH6qRgLpQWa8uKwGCmb2E4mpXvsBYIAqV3sGRmCLwRphNIRvmy
bbBNlZsajg0f/ef8FtnOC+hYXVTzLkVBRIcNT7a8TZAIPm2xvr6y72rUGJgWE03L/pEcKfvYC7Pm
UulakuQmjYtAPbv/Ru0NejNrYIkEnYs70x4BN80bsBdgvh8v1CPQeawW5ylNMajDIN7UkAs3cMnB
Uf9RuHE7OWhW3jSx2UlRc+R5Wi+bXnOZBZgjX2CnetdDe1p+3prcoeoyk5y2HyPV1kC4Cdu6ANbN
ca+Uih7W+NxPh+UZx8PdFduw8uNSl+IBUdfahVRo3Jof8kl9RgeC2r4WuLdYxjbXhwJhCP38KaiA
Viyaq2qNJKpXrnDrnardvrPhbMF+q/mfy7Fg8wmywlqBWChpCb1hm1atfcaL3lXjpTe0/PxIz4Ef
6ILJg5iZi66Jyw67VpCAnfq6Pi02e19pMh7BtGJj2q7KVI1eiLNIObZRPkK6T/0f6V7NydSiP46o
7iu6yfZPPpwe57wX5YxHwKAOK0czt1ioata2/xEHJUl4aPIOlW81k0FCAzBSXdrD3V26Y1qj/GSz
57yFTcRBhs4mcEbhq5OIS7inUrNi5AxAW5AmwA8wPN+DqGF+v9VAlb0aOQsxIySinifJ8ulI0ha+
EkhGWME1DitWOA4i0QWgkKVDxem+fiamIdwf8mgsB5mkfRZOkvqXpskq4YtSOrr9TyQ6QC47B9ca
v2BJONLUOeiERFciX+Rd8fDREdjF0a5HHz5q/Fm8D9ayWkG/r01oFzQ7He7qXq3sDTTHEiHF6yaG
Rmw37wGBHMiYJWYy8ufbmoLsGgFQ4ZK2b3R44ANHnkefgksziNtNF46BGLffLMqk0Bx410UzQiGX
Z5CWWoOTd5z15SF9owsVG/fPhhGmktDouF/KrwvOYKbhFdC2CG67w7vayx97oRj6uTr6Rn8R4PxZ
j51TKa4So1qLy++7JwW15QTJSsLKODkNWmSJnki6fTn57VjmVw9a4NrcdKfFrDxFXpgJ3wTMFKfB
1GWer9mcuWKZcqpYuuLgqTO55kiy6QKhmj8DH0bOX2yGV+uR1gAJ51GiZ8tlytTTm7qf8lX2tLQo
LydinveYCatfLhv45JxlhAxPZbXmcdfdGu9AaHKndho9sTXn9mOQnXFX2OtGsnflzsbAcAY0p7P+
Kh34s87WRZ3xJHZ05mZmeNkR3Db6iUYrQzpjvtAufJ8xDcMXJlmMNjLKB7FG5d2G/HhI9NBEowBB
65XXZ27H9z8K6QJEunVTwjcefHLk3TTixCODhhNtnGEMhnxt+gA5H4AgUclcAbqF/MIMA8E7lto8
HrjM80W4baDzslSlNURlXzvoRzKUstmX32oaOtviGRJwf8e2jhJH9dlvkCfcv47cRy0WqadbbWAn
U4wXwAXGKCeW5aev1S/Og9/CtYfD+KO91zrPhzE4Isk+3QoU0zwokQHvd4KKhamlaByPzJLjQGTl
29OQjg5PGrIJ5BWI4DWXjB7xaNuuJ3/pXIdPA48EBzQOs9vG1vbAlg8Eb8kKcNvRKeTpn1hwVQ2K
SasanjyPzJ0EQenMXq+lPZMAZ+LYi7fcLx7g9BOFuwfBwzpLiLL79AqkTxuQjlt+AV1oAig++Hos
HqwoBQQpjfaVQRvFuxf44Y3lsz2VXbUhzN/3RRO1oPmIDvosBKuovKEwBL9MhnwdLlSJjtYcupg2
AzFpZCAtT5+F00oyTw9CtWqk8GPavDqb/7eXMRLmnMDE068RC4MBdG0dgKIk6j1U/V0CIJVGJy9p
BvKa8IGTnytCYtT4VBubSlWiVQlqBITQ1QH6ImJnFXY0zf12mUlkBf5ZmZS/0iYa6jtVzJjswq06
eOPfbMqdNB7WsSRqgkRnEEFxtinqw26Fx6gE6hq+G02z8ydjK+4WYG67ZRn8Sl8KL77id8c9iror
AUkeyIBOzXtLJsRirM/DamZfLV/KKwCF6Zh/FKPtXlKpE5NYS1fO2+xqP88HieXuEHDSdbEr1kLa
pq+8JX9XjrxLiNUkRuuGTADZ62+sqUiMKyxYnJxKIZ8pyjgZxXKysx3uE0s5eleh5fpvcwCEXSdp
Q8eAnBpG8oyCjhRV/4gzP8IyM3QJJl+moTGC36H0GUhFJ0uUPh+2Y7t7j1d+07zj8mW7vjs9D+F/
hcAa9BkfV9KAylaL5pj2GBv1NJcKjx3IyouZoRHFc8/ZfD/5aQ1PwhRTzD+q0DLV/F9Vz7HEVM+b
YsAoNpZ0uNASa5rPiAUfu0ObJa0IU+5p59MHvNx+666rtQaEbhgAlQ+ML89ABQAGqYHYeSp/suMs
E49IbksC57HHxYfrSOoC5WqWqz8uHTSyoeHFFGaD+8CFeFb3tKjoesxxJQfWBdmxha/xbfrgNsKP
FvAPHilCdcfzpi9nqnlcf4jSOupSdvUQp+QHPAV72muduTQeBGF7c0IG2xxFdPVHzGwMf+RX+rEL
Fhr1sl4e/gxulU9kCPfe/7VlY7yoOgtFixp+nKsX5QMjt4qSS3YGfXbxWQfoIz9qZJPldrnfF3Ej
q3uIuu3ytjlL17ab71K43djeDs/QI8aWi3G7Aqs5Hhcs8jdyn+KSrfAaSYewcEBy0+pe7dqBu2lU
+X/ywt/WfagsbHZkE4Ax24ga7aqAuMCONyhA0X/+spCGJtXPBVJm+l2iGjQB1w/eppRPogyyK+Ve
KAWuHPdvc5j546QYLGKZ5BRkEwlvY6xqiiRQRfJBMQgKshCmGfYfKOhzS/C2nefP9aNVdUNgk+2m
bR3DWg7RbVCqm+pBwKZjUPM/uKPp+D2S8LE0vwAEe/mxYDL6Hc8lBx85nfVHOevzPeTXjip2+Fdf
c8FFYwSAVDMiWFMHmTrxKJ63Be3R/JEYd+LYBPLD4xbimrSIBuJfSEgalQw7VkraMDfHJLqgEfTa
Ml8zuXVWEPIAhFSvAm40d2O3yAVcUE/LQVO6ancf/+XxOpKrbHZjPc1hA2XGwGq3Tw6pOQZjFSMq
MBFbD2zcU4wHoso7nzLXHdd2WVz3R8YFIzWfiS1mNfa7sAxlX9kkdew4e1ZHmrjXLR5WUt2sXcVo
rJFU0SFu1c9FBsSSpyGfzoi8Q/mDJC504xYlRHKhbFAFrKw0R3TCR8GxOPOCwqDtub7rev/Ihtyh
t0r5QxPSsGWK+7NKMHtB8XKRFqTsqWBEznIO/DUbAvqr+Slb+AKFQczyYK6NLOnl0TgKnYfBk6D+
S/f6E0DQkTu1sh7M5wfcUTltVtnzpYmAo6n9CUHyzohKjLTXy4S2kBJQdLQ5Sw7B54Ua4ccqKvzd
JSHgthGL8TfWq050lSftylyJhBMcIS/b6sW1UWoYPFZhR1KlZf6pkarHx4XWv1qmbIPajuofJfUi
4SB0fFUuikjdH2EIB99tJRqTUgksV2jjhxx0NoSkiDE6jBaei7UxUES/wVkOEEsxfrB264ZFdMdl
Rbo4OVEkHqhnwiASkY/+kAyUB9nmFk8acbZqSUE36jtffeYbxg6CR/9KJj0fnRVy5Nr6J5UHdiob
gScEI1f4HVqD/Glcod7sJGPxS55MqiULd4dT5eMeiJJPnbDNEWy45znPZ3KZJTOol1w+lm7yTqtl
qd6MjHT4j64/CizVB/uiBTb8jgJ6GOzbLM/WTmsA0MzB6G5ijzDISWqA4nobgYgYNcN01kEz0ySu
lWHVY6fp1qYDBkovJg448EA/aWnDA9AFKAsqVT867Jz5sEHbMHj+FxAG9jUm147hjwLyatt2Z5Av
//Gcp0HvvFsR+yJqIsjLp77Rch8JXBggCFXKFkZfCKxfBwQAclXCMhYPQcQZmhG7PQqWfd5Roumr
SJMrZDE8hjcOHTqPzkStNLILWybM/kBTzNoQz8bp/x4G2rZpL8u2fikDSu2+ou+jozFQl65pW8Z7
zuDdTh225FFrd68480kUkTbBBXtXMlOeC1DOtkctWkVLC+tPQrysurZfLJpCPUn4qxvoZcwCf/oA
YUj0bCNprTcvFP4v5FoY/YLaPZDx33mqvyDydOP3fHEDR5ZDRp8m3hs2DaIUPupL01/xcnOh0K9h
m2+1FXhMleNrYlDRIzhOplf3ui54apdxBC98u/xI3Y1sIFLbLnJWYEV+HBUb0+E3kKMiuXl7Jlct
d2gtD1pVQS0zHDoeZGY7VjWLKbqDiAq+DVYkhMGOrHtJy6c0HXrY/WC+m+U5HjarM6nsB0H3RCfp
t7lcdN1oLTkcCBt2T7Ix6UevzLmwMuQ7Yw7wave91X8jezqGGu/+1MzouPBh+ofeis5gEowjkD9/
MgG6czhIhsmWSS3xn3ntjAtXoe5lbLg5wiFaNNv0zt2pMTaZtJo5SzqfEsRel9Vt32qleyFY1q3X
I/wbg6ZNv0xeOoQAmOsPYyBaVoozV89RHgti5eOaO75xwzIec32Klj5Q1lF9MowBsZ++Wi5B31ZE
Wvdgd/nGJNXgdWtyvTP4ov5VV4SZPat0AvAa//04E6poz1bmzOdcW7X0AHwEGRrZSd2VB91+AY4c
64eETEOeEZvTJzOIoXtlZ7TlIRvrbTmBjF6joThzP1/JmeFaQvQXYdQ0xmWGKBSsu7ZmWGf5X71B
iol1yUhL+CfMmPT8PtfzjwIdC63Ef/PLL3em+ifQ8dmD3Fk6kSQn21ubf6GftaVNRm7tk4LOUuHQ
NzjuD66kLXQ6jDOIqTa/CEHaJfP+7p6B5F1B5S4NKkxJA2xmdD7YWBsw5F9J+m3HOMMsaP4wt0zI
EpsgDaHi6PgcQpHKt9+SWXB8HCSCsy1cms4bQMgSDmo4k0xPTU3xlri87YYwtmC5ivxw7uxLmyi7
0FmMKd0SkW2ApXy825rID2fQB4MDVoFOQYokn6T0fD7HPliiQIf1gmvmdalFqTAJOl5TeGvTiv/T
Z5p6NY2FHXAUoHpRtQnV/6+rRebTxuBhuXm4+3VwO91J2ka64InYFnRzaTxRpKBys+bQYVMf507K
SEGymkja/JBZbjVogTaoUOpWoMiEbcEoQ/2VbE/xzelirxPPr3UlZqNpL1jROoalI6/ZYY0PAW/o
hyQcePqtv7WuWpJuaa+0deW/DzgnginXR7sy0vBR8L7XfKYxZd3V2rE2fsNi0Dx67inwexv+K7Uz
UDHZYDSdP6RnnkEr3iUNFILVzmS8Wl70AnEwA+d6QzuPJYvklvWhyFCi2nIcrdgueZ4jYMf4lDoe
uK/V9gJ7CcSPgP98hF2XlXSH6ff97XSHlbo5n4X8Aaz+pa04iqAUMfY8WERKbfbra6/Ktqt8D8R9
HybF+z4mFKF3o4GUMCXVNdRCbnOPdT+EPIjgT8qsJdHLiVqVXq7gDrz3vG9vSuUQ+c7NlGV4jghy
/hqzWbB0wz0/0cO3TXyNR8oSG9QsauHbOW6gCWpX3pgMqLtCdteknxuvaCKzjgsKhjZyYxty/Fv6
kPcdSTWWCRGYtiKXPYXUBXXZIc6kdKaDRM9DPJTB5xd67DI/4E9OP8iMpU1/zuJU3mKKl3QMn/Ga
4uD1rSpAP/4r0iQ0bvoyb7U9stCNe3FdMyiSTVRYRIMPJDpUVLlQQodHOyPW2S4+oVGzLMTLbRUQ
/V1rtBWmEtOOECuR8Trbh8xiErkoXfw8ZTnNJ1IMBVHJIbg9e0/hxq7/urYlXQ9qISv5kCFom7q4
pZ+OAIPZJWbCXGk2tvbT5zY7dueLYhxKkRlLEQW3PvB54f37s1R3w8PCkpJByQK8PMM1P660COIW
C8ItB07ZJyiyZeWzvA3ZGHVW5A6joLv+J78dN/KGnPlALQ5O59V9apq7/vgsmFbQHac8wbHrwJRW
KAJ8ZJJdwr5/78VDlSbE1dHM0g4vvbHNm3n/dvuDeEFzPedLUzvClmJ87Sx6jG/RWgPcDA5ym9GU
nY6FKWbUb03Do85WAIhfTC8zjM5U/Hgzkdd9qyDY/KoXrkbBzfB1m9n7BWUH8GaIrZTRZ1ZK9kpa
fTzDza0Vhmmj7zkFH95cS5o2gGJetYjYWeyMPLLWMbfxPDtWWESKUiJyP8hrHs9xi+uDaCBGjr7H
pFKQch6a1PkAW6hJ2v4De4OnmV/d1SO7y/uihbg1N4r+o7SnadU7UQpUiG0xyIKJPu5L7iJU2FIQ
Cg7nfJfCsivHT3hsdLafqgWI56Ab6ujvNo3G7mcx8Y/5pF56fS1zQS5fG5HApLRVEawzf7wsBCoa
jrRtka89mtVI4FYIVW/FFPYzg9JTAsRr2UJ9gGNImiOJ6Wf21bAHTP/g0NCJD4FC+8Sz2pSC+zqk
o/rs/VhN28LiPzHdX2rx9uGD286FX/SQ47kiyK/nAiVJgoCItpwcANpO5KLX/ptanbXaR3lY9G+M
3/g5KeSPAO8bId6bDUnJeA5FNpc/lqrY+Z4YlyvSWv9ctEKIxxb4f4/dBPLwpLVMVTlowY6FbEQg
YUdrLUlziJ9Bzpcm50biUNDEFZLhfKewx2p5UkyONZnFeoX7/81iFm8uUGlC8hmTMTKXoR0UaPZJ
9xtL/EUpFFAKGAG7HhE6w6t+NyxZ9OvgFMx9PxKK4BoudUN2HORC4NfIUdgI4jyTpvMoV9f0VVtP
OWoWefC7gA+8PJ9Qc2WFhPmet8pa9SHnA+55SfIp60VYS+mL6Tq9riseS/m2n5VrPskspp4uidpE
7h4EwTAE+YfYAJO7QO1Z2Kbs6fR+g/0H0VuFeEBCC3PMV9wg/JhU5Ol+gDRBZcCFdRtZRzKVsqMO
xhD1j6aNCpVj+pQ1N0MYUOT6hCyRcL1UP61+HNpxVDOIIAP6kZK2PoeO+sjD86LlpjUC9owOAkL4
rUAWB3oFTvEAheshIgrxXaz54XY6K/RAymrdmyMN8AWrij9XWyFDc0JKGK8ekPNndsxDcYbPB3pg
UBjXh+T0fVKTJg4HahERt0/51W2omxmE5nLwU+BMv8WpUU/PdhBLW+2yf02ByxAo5JxmHJgTk36T
u8SZzuSgVs0M/HfNAcM/PrH0+OB5qLWtXSCHVspqp60+fzAa73bg9p6awr28ehsUkWylnk1X4nx+
/IsHDwFwsUN12EiukCKEAmSFM0TYaWX3MOEdoDxAL8eKodUKLNWVioT3ROCamSgocp/c6+kOeyQW
AkvnYk8Y61LB6udq8KXiS4yR2clOkidZpdQGUsR5cUyxj5V8nKr3kvSD2LpTewhfUvokSMVLBgRC
U7SQaJ1R2M5OF8dgqLEkcx5V6oc5PQJ2HmW+x/1iPxLhtXTBqMAP2trYlydLI2bdM5xKVBZmHS6j
yfRKiUbDdjIGYhb02xkDTMXR8VLWKiMrojFtvdOJBIgWXgyJYhsdlvlpd5CT0R+xFhhuOblsqx3O
wyZbQSeNEMRyaHV2MUXuvF9281w5qhhYWS4urVqR72nSvLKablCC6RQY2Xu+pi+GZuTb5RU3thZ8
q434Zj8rNe0eBDHHcFfrFoO6F/6cBTpyrb4XJPPEifCkXA7rcghS2Yw1BkZmZkwuwcExl6wXf9Bg
BwbARet4L9R0Sqa9sNUgitmE57YsyWOyESg5uclq9B5r6S66bFQjVgfpAYtwQlS2hVfVYKUBuIdK
i8pgeajFhP6XCiu6nwtCJolYyvXpFGRYyyaG571Gavf/OhMUGx+FUzQiYYzGvOcmLR68/x0zWa/k
EcKiiTUaZ2jzJ2b9usLu8IuhXu0jHLwYi1Z1jyRqAAoTro95cqbswGnAUI80QP4YQBYK0vAqQd3r
RSbpVLMwvXqiLlKFxHzclE8nb8c4oRrfv4cREaLek4Hj5TBBGvd3k2TnZGxKDQAwZbvzCs8p8xFh
h8P2FqmmU50cEj0NFM68ypqbkBwsW37cHqUtAPLS8jy/bpmPdMfkRQeDGAp/3EieD/dtuUwROk6h
1FEE45II2GuhClHugKS6793UN0G6iAZ8XvzcwfWz5BDwjZ44spww9Ed1L/VsxNLowZcbXIi8L4iI
OhEqRcZDoVX81Gx8LFdt7UaHdkTV8KtLxApnacFfCRJ8UaHFhN5HM1xrsqdtYjAHyyN4SwezoVzu
v8Yn7MLM4HXdF4AUfI2KKKB36o5UAxa0eXt9pZ3qc5OdIfJdPa8sjw1BM6AV3DRkbNwIdkb6V4vZ
Ryx8QweW7u4g1YrKHo7hbv5MrHp/xANAOcOlFZTkZf8v4145K03ShzYn7NYufGkoPEISxY+KY5zy
OGUEUYD3F9Jwknr+n1lKdlvPf+l64cM0ActSzlq17WPHsIHHO9IxcggNCww2izzB9/VDl+HTgIXY
tLYUiz2O8+VO5L1j7WNo8S7M+p+zI8xhq9169rLXMPnU8l3zYuLxotzHqqtoW68kaCG8ypFiKPo6
86GAKAMF6ZkX0lN/WRD6k8X/c9QplPWnlmJQ1047/H8e8Zok50wIiRV3SyDzUwGPj12w7eAqxz/Y
v3/58x9AqKVIWYSOBXLNS9S+p0ytFNm6q2i9hnLfUN82bSBOYR67CbzGnZXBYApk55k6rrGS/+Zw
a8EDuyvrKR7WF2o/3V+hqho2HMNQpls3oVm37PFtxqIFsGVriLEWhDNeD4e9/jOFSKIMquNTQ59y
HqO4pDvlm76rvZuR4Zq5KQI8SMM5hUHwplioRv0vJJrN805ZDrCUJbOR7mJvdxByPzdyi1ScNxn2
N6giGJ0HNeYdXKO0ANN4BAgzGMh6NDyXqiMi4UcAKdhx/wg5nNfm7rPmVUEZC4LHV7u8uWQ4K7sT
BmgnHqyblbK/BEGP2xD1iY/EKPiJhE3ONBarb6zFMtzilFdiCFjBmGaCTVYgjIfs0n6O7u8wGRBy
8CR+M8W+xCjyBWq4INct2Pe8lbqAUQraD0o+HZ+h0Z1HrTGZkSZ5MGeke4bYHhZPYiUVzvv/P018
5YLzyWS+WBkZwbkVIZYgf/svgxd8GMEFXCh+LMFxfIInPFBTks8dfMztrgiy9PyB7cwal3KahMVq
JgosneamOAOTXdCd43ddrwefYxTp5BE4c4IH0H60jCoIxKHMxqy9NcncrphQnyJQuxZsVn2/m2pJ
/s7GXDJmeb/2Xen4KpNDQCuKJx5xJ6ruTp6FBs7zNU6AfX+MndMEcWBKWMEolSGrhgHszOCCldJY
l2NYp5C2ElGFSXM0teLbkTrZcvgr4JUiJ0tqjdq2kuh5L8FJAxTQQIXTFvaS9D6+TBKhW28D45U/
W2qq1T0jGHp9e33xT14gKdzjOcBYQAkCHmh4SvEvoCt/E5oeONuwRUIF7KWqzZU9ve24PLq798XW
Ke9NW0eIGxzd0tTjwroOtjxcq/2Avi6iboOccp/3jnx2bhixvQf/+0Z0q97rx3iOSx0ga/T1kLpS
kvl24LR5F10EQbJ04/JUhwwOexKzbVAwvx/smCpaAARhGcyF44PUG2gKJ0wdIOgVhI4FeIr3YYDk
0VLh0OKksIzeoiuaNv9gyMYZd3T4aWwQ77aN4ozqSOeamE1+xWx0YodKKBp0uaokKmKpQqmopOxH
r5XdL4Aly/6Vo5+rpsiLqMM5w8ImSVJ97TvR1qYzicJLW4cUjht6911gEy01q5642nFYieS2G05f
0y2w4JhSmvexmkOdF7/GbzaH5n139TevXXh5BlxDm8N1ErAVv95nkmi82wl549IBhAlNpLW1Aprf
ucXO4sy+5leWGBHwvBAxKHIdCzHX36m55Vh3ig5OxEczwdEIMBkWeZGAXH9YpLfxFY/mcBKKlbpE
f1LAc8MCNj4hmqlYb7ZbdtkFeBGwUHi3TqRlQoHOdVfqivJs4HlQb7IwnM60j8qkmUUkQzMT0O+M
YI0N/QgSfUMufGfk03afx8FKO2nZy7TtJu8lhTWJsLx5aSUTFcaeVFFaBvN0uwtIsg3RMkmWtZg4
lfHAf4QosTuvgvn4kccfCHpr9QsHo+rQsh1mKDMB5mhdZtF7/JdVpuBCQcT8dDInwwKEKbnFPRuP
HITGcB/UZMBSeVhMBm8AHMSHESLNCxlFBImSgarOgJkyGZzmgakTTPXOROntdLS26FcCPQmzWHZj
Tk6t7QflSL8dfRrQyFPoqZRcHhgbK0ql+YnHUP0LShvwjtQsuQXdt2ZTH/uoVf/evrAdscun2ooY
BaBrL1jEumbDMgY2l3mRIcPZzx8hp2v7K3EkGORvMesK4E14/ccONaWnw29tNIa4jWfnDfJYLRV8
vdEM0vfLNuNQQz+j8ozKPMgvc48YxnvccNYcAymQNP0LV3WNSWBypLu4Oezf/N7MCPRMcLDKzMOb
0q5heaxKpWE73UdBKUzuWXZWuN11isJVvsRPXLIYvdaCQzJZhZ1EEP+DRwgyAadWedksaSgMG2j3
krOIwYe0SMRE9anzOEhE146NNi4LmrSgXMNrcKsM6gvH0jx5EXeXDbi1vyD9UvluDeGrBEz8Q+D1
oE8Qm5vgoPUlhIzXM45XA+UZPkqL3zxxHWzeUQf0Sk1aTKV9Yw/8HTXhJS52KHH6Rw9CWpjvf+px
1ymA1hStJ0gCowCI+mA9wIN/bmxPL1HNioygSt4FSy3ID96oZASSomGwl3z3A8Oy7jsR7WfaDJaR
FOoa85J5IRu1trC6EAcIuzvUknP1XwrKojW7cL07hsxMmat/JS9pNPi4aTwYS9qC3SrVCpKylPs0
d0Xv8+mB8ppryPVVmYNW4s63IgfL+UyMJ6uAeZBqglLzUHRwS8aHrJ6iSJU21iYVJxOd1tk/RCix
pIbGp0LD5wES71KpBN0eAuVlhcXzFDnQ99ef/hs2MwoL/L8/i4k8OrHVx2Fyhfe92wT2lZjpyNdg
7UCAOGsBzC/g2q8XiMVT+fAo+ROKYiC9f8gDWch4g5t3f7plyCafuCQWY03RkKvG3QWia42/E8Cm
AIk8IV9vQeLMT77WplwOXB3yoPEhFVc+PuQIZzhTgnwXrfUxBhg6mYDYuaV/MBsBP019O/WAZ0mv
hQZlMN3gII5MRhjiBMFtwyCfDhpRo6i0EFKOgfNXufpRZCJAup+tdrBbcjiqKvZz3bUuiJdzA65W
g00HcQN6PBJ+RP6Gs3kCuDJClGBpzuNZ9WFFBGwFlC8JbjvGi61AQTJpX3TcVbJzDlIatBZgS7vU
4HLMSAurgs3k4ZCOUYoWDRv95yWbvhzbOSXPOKipu4+cqfs7dgmfMbwyOMx7jXsAXHk3mJ0HlCpV
BWVvBSTpz/Y/2F7E1TAUj05r8gpXa0tdaDcLe+co/VFvQAQwV6d8rDJ6z28S3wVg6DwQ9VySojvL
RcPr1Q52+FmDlwI+v/gti5fwDTO7UXbyRaXehNQldK+VtstslscW5fyer2vO3UqihVspPLwD6/EA
9M+olIwuKjt4+y5Q7vRGXzvi7YoxZO7P4RIZAIal/AEzywWg+gVa8bUd+5CxzeghyoWyfQolCuDg
gXJKUr1tEj6dwnf9M1ArQvXcD/OgqToVeJ0M8mMyiJu0TUORHr/aJfnExpGqoxdbNmZ4Dpku0Q+E
RYOXJyrGGlvsCHIMuNhmaFALGd61TyUGp11Jg3SK2igu6NZz5AXjMsOAicnMB2hNxRZaQToQyaO9
NXwtbXoEkhP/NB2NF2zOJNNYUq2c+kQks01P025RL6HfQBw6XbGGzz8uwA6EmTZUd0ugu9dQPSFe
aFAEQ0AhqgEnOJ4OfzR1tAF1INaz2rgYceokDYYyUKXVMv0Y1uJUd3qhrk5QTr8AoTkJFIRsgwcX
2+THZHOMdBsTCtpFy/PjSrk3PwmfXWi4QN21//caZb9qv3W+7ARhaZKq55yrNKLoYBjgEjX4J0P2
ZFLC+jnYFkqrKOKXL2HkYR/ruLdknGgblrH4qSC4z6/f520Jitc+5VydNg/OKfof0elKQE8mw1Wf
DxBbh8E8pEabOzgjw998UYZ5eSyS/osP11WbK4uUiM0RJIYadlrx+a0w7/Lr3p5mywaXq5Di+8Yc
ClkdcmXDslEgOReVq+9d2ZY61wx0e4gqECyXrrOOhwvy2mkilei94wHss8WGPbKbPA4Ag1xfLHMd
fKqn9U/5uBn1i1ggY88ZYw9RalSffEqabRqdH8/pnibV4wcTY82Pofx23Mwus5O2hai9wIuCcBTA
KsMU7hv16CYl46nEHk2R9sYPxiU6wrXCCpXT5peB3XPE+OfeuMrLhbs4eTGgPR5kdtUd511ZWJzU
OQ6lBF8ZBKuV59bCs7ihBhZS9L8LGORZ6M7/WbZ+OOJKYVObvPeIgFJfbfYzOWrM7WgTeKUeGzLX
5jHUDFemvDpjmRrCryIJaKaGlK4UJtklfDC6/u2HoWpOe2ktyMa8kxgEgf2QI1QqbYPnWSXIawRV
Ua1+A7tFu5qDap5aRe3yRiR944hM5o5Z/O6Wm86aCp8T0QL33Uk7WPAQpKQPuX1RNDcT7a+Ozwwy
f8SMD81kxR3Z/oKIRrQLQTicOLc8hycQVnM1zDJB1Yo/WJV2Q6studThAmA+/7rVdltLSVVTGxeR
pOVGcr0zGZv2NwqpU9EkwphVAZMV1OX0sly9uDR5Exr38fvdrGFKyfvHth444wySFVK3zo1pFtjq
YGpXRpyGnmSwvUbVLbC10JxZse/gDHTt0c45qq5LKWVTcbsax7CxEJLRp+rgyGUAW4RIVl29co80
rQdinjCluyB22+7SQVJPc3jN3s+NJL+co0tFDCrAMphGXqcfO5RHrStPhFihTjGDArRGPA/gzwKD
sF/ZbxWRtkppE5h07wdFAFj7VZEgiqmeIjBXfLfsK5hN/NIw8n7DnWSmq623wU9mhBcPkRfcLL2C
KDVNKygINX5MleMuzuZePHo9/kxWaPrNo/5O99Q6GEWIkx+USio6PYCX1GyFuZqAmH5lWzKN2sJa
/ymSojrPF1Si0yILl1CFBxmLR/ukOWFvnyzmUGSzJGOzyZ8DmnuqjLmMxKTecvlIsSdnEvUX3PZ8
djK5IFg/NEeZfHLHpJTWbz7efPHWcl/b6ETJ6E1SRoRdt2WhnIxpxrF5Diy0R0+tNg40MlUgkgXL
sdVlS1J8cEH/zrmSvHptB1q3Ld3BKsShEEfBMZEFxcQFsBGd6vR4AzzF5nQVrzf0WxgJZMOp4tRE
fzbZwk3zd6u2GMFyuLy2PEuhsyCtsI/4Alx9UunTXXeRu5Y2o9Gk7Z/ybNuV6hW+OtA9MJGp1H1A
sVjMmw6F4/cQzWuxE2UsIHXnwyHycK/5m5m/32f04rp+dwHN2Xi0T712q6sHvoIGT7In8mcgZYAu
eBo/6vgWKbM2kY8kpNaBWpNTP80FE2ysHKQjcN6CvBRBIuH4Fmj26BK3fSKjhzfWIrhsNXAj3qWa
CKdwfmr/gjmTzdwZFmXJfyrh7UcZjolsEtWM2FPP0J05xrZIrKKD7g9KGYy+0cOOh6V46dCW42WW
PZoyoVrjstGZyRiaLdCnpVHvEvy6zEx6jFVl9NltCRNIlq2rG4O5NWjq+78ukVEvyRCzitkCo3rk
5Esp3CT/e38OQpO6mIQLxvB2Seyd1zhqV4u7B3Ny9k8zx+jktbnOpuH+AlDwZHMsYPFiO4Yis20T
m9BBqQ+nHoyXwCgCW5Xb3Ux1z7RElGwFX7Syrl7x51B3FBec6NykrILfTEzZVdpPMAkOSGwiKvWk
ozAoqw+qRMT/+DPYWOKhmZJSSipON4rr8sAQe10NKiGo9scxKKi5M2xDSPlBtFZM4dCeOeEhk2oI
injzHX8GfUSVa/4QOzTaQP8n9r2zxS7n5+uAuOphJ4RPE8O/mQiJS2JNUH3JLlra9G2F8coZIdoE
gBuwWfzQGcTUlygQ2AVcwz/qTZWlsIgubthf1kEhROWnlKrvuO5pkAWB8k2ho+/l002HTpdYS5Zd
HgJc7tWrjX3cTTPKGigAMTiKNGysarzeNnHGxNCM9AfklVR3OeVgPsQfmrabgS84JDeBXqBLhWPt
xk8jR9p7IljYOhh4mb8JvEOmh4gWdeM0uBWl59ASHQABL9h3/TyGtG5RbJ+hESnH9NoqS7owIYjE
o13PDT883NM1C6UspnTu9T/aVr24xWsmi8+2Uc7aTcY6fdYhZqg3Cb+LOd/mQki2gGPYuDTaAXDv
QvckKHVs1GCbWidMwJ4AcKSGJMFt3Ve7qpeTdnnSZwg0UUNs6OOu6Qe16yS9rC0mvbiADROhb06e
YWqz9kUWTOfUU4nZBbfQm95pvqG7+Rcpl0vbI6ITfQr0erHqmZ2LaA3yCVkr6aT8tXdfof9kwvqC
6YuowXXcBGZBj+1nNL2+QWUlb+920Z4ieampxpBXl4NUWYcJkOencpU52ojDE8u2w+SIjVOWaV82
GpDC3jjnDnUka8v6tOO4T6y6Ro0dlwyzW8wRM/OULQnF87Ue7DTfW2tOZMxZVtaHUna5TEWjmHDF
CZqaQthYFDJHAkHmzp/d5jXJIyOVZ1NmDNQFxMp5qtmPgymI1YnLXrKzu8Y67m3K6O2ITlccsfcU
Y1Q4b62woDovBp6NAnKlRvZZPOA8/5KNvVbOQX8CAv4vfauf6tbkft4WtZhjqUjfuho4clCheO0I
lQgqc1iTnDHugtR4Q3g36sMGTvNqIVhMwnz7JO8w53subwImQ8MC7LRV5ZJEc435YSv5ukde9Tmn
u1hYkZ0LYMwCNXrytWMyZJKsjYf4Cbp823e+YOwl2P5+tZ6FvR3IT5tCCi7lw3gujRH5TgwxqnSq
H/G5jzh2IpOt2X6eDXKtvVqcPThhaalXMCdkbuTsWC46qsg7g1KhKcJ22RkEIy42GBp84emD4nuw
UYhvsuvIVhLDglkbmvjPECy2Wn2IxBSDRWcUj49dp1LklVbtKxEN+P/5UdmNw+ON14m+PiUGGqth
2HewHN3PVkY5Hv9tQ7Y3fNG26gmEm8pkc4moGNi9cLwxtwqlMEXxhCEmBPLiDwB7PzFFum6riV83
wnGXAL//3bbT7b3g69ItZ/OyWUPnRBQe3BbwCJfBYYeapohs38nDFtQlbp90qZfNhXwRtKRzHEYy
p8SyG0DN15rGOlLAc+/w3xtXBw6ldvq/T+6E4Zq8kDU83J8OY7vqyz/Ne8IVu3CqUcXXS7HaRjc5
0NUBc+OI3Lmac4QxVq18ngRYtDRmOQwx35h3NpHmYcCEMibmmjhJDo00eR7jxzt6aQzoltFPWDzj
toe5GUHCdX7yh0Ud9qM4Ephea9kOabynx63+jUKZzCj9HhOo1gWaROYqUKq680kqRG31Dj+aYktG
j483x5CYeMncxuz/yEYOvfmYNaeXgXVzglck4OePtnWV8HatpMHC149FzoMmtnJac1ATcetDVZT0
JUFBJgAqB9zuujakjt6jaRupnWcYmYafR3bbYH9+88xS4AWOe8FN6PrdObtJp1ABdadiXV1MqXR3
Dwd1uFbFkUgS5fT1CVM5NKsLt9P+cn3c04OQXJkhp2lOgnfHPxFl+Pim8EM6JUhGgzH/w4WbZkJE
GLi31LEcJfghOcq+czHt8KCS2ecQ2CfOHQNXzY3k3BULQmaC9dU7FglhHGTHkg/z9Q4ygXwA7KS7
mtNSOhfd7IQLowKxtkRKpl8/eBFAXQeTlAGDtnQgAsNJqavhC41H8tzn3iFmpRmE4DAPjK2NWIex
+n+m+TAm6ijNMSFa9nEuaZ/2bddPfLP8/z26htSyfHyfiNhJ8xexGIfq9TucqVLO3doUZVqbWPpp
vm0bYeB2kiElJuF/zt3BFNflVxcuLj5SGKQ8GmYN0lRFMzXlru43HJclPpwOqFdn/yI9qrrRB3XQ
suhSdo7Lv0cUqYTd3UgQGfwTO/sRiX3dmN2g+v8/G0LmqocpuuPacuaZQzwARRTvDGymaWKXrfG6
X1EV1gTs8pNd4pk6FLs3m+eFy5BS3rtzreIYgN8Tr+gBBj0rKYQF1TG/enGw+h0iHTQnBdmqYyUa
CsbnEvjTVbVkjhQNpRtBJsjxvOgAI2+fXK713VYPmtHjrWGxPHWfZzjH+97mUfkdsnkcI+X5G8ti
L17Ok1qtu/Kp9FTbat/Jn6eIZcMPw0pYHI0fhzJ4+wEvozIdvhEeCFaWDOeARfyCHECedxmJqHHp
ZMCHwNF92eS3DzHsll57hN7H/WNxgTsVilmUvnsFYRFBcp7xRxeLLqhVeFc1V5X+KajRNAE1egVG
LkgQwOY9V9rQcGVSWk22h8DUQ6RzhuXF2AN8x+mf4y+Ush2DFBqbj0C5M6VAyr2UFjEg17Q1mIGa
UvCbEWQWxblk5MeBINJMUdY2MB58HOvUiWQAOyRh9aFNBOJ5ErUDDisoh204pPQd0qqhHjMp0Js/
tdYdvvVvAS5gQNJ8ZiRg09FEip464YN6QUT/xx69KUyv4tTPYCU8SF2eVWxM/owqNHgPNH2FSPoO
jC4SPd/7aa78UqwqYMczgiOPQd4tfnHa/5n9D82fKYmdb6jBjVpioBDyLjEpyjw/XZr2zPwE4FIf
DRicxp5NJgEFEiNxXzPLn6Rod9bg+yvR4uzawepDq8xseMTGD3l87pBoZI6K9lRAf0FGXCyYPsLz
0t3l+MGfwpHsFKq3pwUIp7wq3bHZyk5pa6xjR2ubfsvk8Z37K0GC7y1ElucRpoLx7tTBFB0kicEe
j2v8hhBp8Dy++VouJvkI9L3RPpMrWJWg/o2Zu1/WEY67PTgqqTHHlyH9rbetxeG02V2764LZXUp4
5z3lXgqaa5EQ5G5DhxDRy/KmQnqYXm256jSjZjqgpTNDr4hk2wbG3/b0xmXsl8rerbG1u52I1vBL
AXm4tCkrStwp4eZSYoXuTzPvRjYW2D9URwUd9LKpmhnzYhY8apokONPMXoklO19Pbyi7P9PV+DVO
xER/gYuuQ9IOOMz6JUMuUqGpz2JMyi3ou362H44RbavRJ1TNPT6Fs8UZKfT390dxN7+zM4aQQbk1
IR8k8vy9FyWy+WITjvdCOTDJJndSDaHjUo5VwbGjcZ819sSa/niQlzkPgDRynNNkm7KtN0kF5YIn
CW7fCWDciuiIDwRus8h8J7NxSNBQ/LSqcuD72zwtg+WVG/NNn3GiP9KxCVPc/0rdVMcAqVS98zoT
XOMAz6lFOB4w3+c5vFfCYBZU0T3heIr0zzVndSDi+LnHjcoYBzyMHsRNJbLrCL49+wBd6Xah75ze
hPYEczoyQfLNPcqJ06ZXlZOXcZykJ41yovkga1aOK7v+eWXS6WporPW1F68SZL5bnPc+/kH+vqg/
zq+c1JxOZMlqImwDzC92fXsKBH+L6uvdN/KWPrJyRbH77w2yJnw3Za/Dz9JYt+n8ulsOPihEp6OU
c5fbpHPfhuGbQeljL1G0++QkWs8zJYNdcntM64SxlmVu6adSyA6p1yJtt72gZCEu/7wj8kWYaRD9
/2BktHS8RWTJ7QzSxh3RfjfOCrpjkQF7iirYT5RALBAnJiw14oTMIIPURUGaqvq5eQ8+RHrFFDIm
TJEjnqxq7DL6cmbseCqctlnBTlu4Sc359jz94rd/hkPNAPghR6fGdIN1k/gyeZI9vK0CSF3OtUMC
U2dUNnF2KBzeqLLFqYsqsz+RwQ9jHrf8KZUm2uZjtxHWqbzBm1TtDgGilqXBD4uUtJ8tSMyq7ICN
1ZxC4pc/ZLaSfIDJEuQQigA3g0enivCOWroK69OzGAmRPxlTLORaemlPPlsxRA207MHg+zjASqnu
T9d7v2DZZfWAAeVGEfjM97qJwvg5kYMSWyXMf1POp3wVkHO+IUJp+It0Q4ZRw0iipHaoIe7dMslp
qEsZbe1efEkhtoyBu/xR0qxoODUTGDBzszQllp8oZUs+B1xqVLcMeSdCpyCsu9a0Mv4TPODMUclx
D5wu0hSMkiTl/HrabLzEoDwkkMGYJlLG3XTNMkfoXiztvmVnIEapS7Mbfka5J6X7HisqfNNDFYDB
b+qQqArTuE5X70vaD9NN92FYFRD/PMxGrEjV4aG19bMlE3am6zxynwM7hmS5aB8xGdh/G1y5+Q0t
UP72iqWO7dq2ZCc+qWYTdjv2nVzmhy1SkD3cpf/+pwYk3qD5RmLow0ZQyX+uLqfh1r2b/vTVskSN
Ye+lLa3raurKMM0BvCzUIZVrOnr7zBlWMkRkbgWgS+uVyY24ak2Ugqv/tiZmB/IZO4hBk6e1dkIh
bbZOqzXr6rJa8B/lve3B7o91JkucwbaT64zstMwVt3h8j3RDcOirr54Ey/U3r6UtEiLQr3lR8ine
aWfB9yO707rBkL1naRpGSdd/cV7FzKIQecImCPrGlG4Ipesug/59EnRyfxBS8FUxIXzulEGPMp+S
7j8NuubZHYM/mhG2LLKyLvdkVul6F+OiPl8odDVysqCBjjrkwRreKF8Nzh0TyIQohPB5pW9XIeS1
aD6aYt0CKMjfUsYpE2bl71lJszmJynsd6Sd97o4VULwlwJAu2XDl9aDpq5CmcQp21dA6dFvNxOJV
WX+Q13gQs1pMe/RSXw6ymdHENu9axShsb/E1IN5gdr9nuKv7qWAbLcgKss4dMyQmqjqWEaNqvBu4
PyPEUIX6fwvaeVqDVk7RngeOAcOLnOtnIMlcL2EHJjJHlIh4ceZWe6OevNrc1iOZ5KDdUUP0rKSP
WQdrFaSWgIWeNERFM8igOyDdxnwKRFdk7/hvFu46RgYticUjmrkf3ZFiUiUyPutt3Ked6APTeS6h
P6Cga2dJ1q25r/41aPWq8PnKfKJ+qSRMylS5c7kRhZ/z8Hy5lXO8vI8T68DDz7V2MOIakRN4uCbI
YApWLjcICuWt+3hbU46LXWW/R9AYf+1arRf/x3IMoVgSbm0OkVvCaqzz0z9Ogd40r37r9fAFGZEq
43la+RgMk+ImV8luyaSHOro2yWx+WXZ6abgxiY1e6vQdF9BKvbt+t/nU0078zA1yHx8kYaQE/VRJ
3xK1Ys7JkIhNcHfdXgnfuiQ+nw+Y0yzixiZ1pQZGrfTSPfWljI4A0y3qgQ9F8Y0hT69xMDqqB8Lp
cr+LC00qteIa7QNF9B4q2AXSKWzrLVOZj2H++JASjN38esbegqwVZcR+PL0zqnKYcj5JSpG0vFtn
QsDgrmn6JakHkY7jYzIAHGDw4HRXFFqSLPm4K780IAIu0aQLoH9w8a1mWl9VXB2YFdpl6pZUzjBY
kaGKj13ngM/wpR+hVvy7b5MaEsfh1Ht4FG8MH5setj7b6OEMfBpQ6YtHj7jXDvMijBWcH8yCrwOE
kGOylMmYGHicFHo6dnNigKYWDfD3LBfDz9by63lXKbKO5Np+wH6dmqLOKCA6JcbWQSOIWvEYek9L
cLw0sL6150hwP7SptBxZA3ibtVMyto6c+l/+JoalfhJtKgr8MGy3SVHJ1px8/hGAADOxazRHPdOc
dMPlwVQFczPU/QfsaSph5tDlWwOQ/qMh5pnHXXhaJJzjZ047jQPIQZ5u1owdMRTZfUYcG1bmO1Zn
/8/FZ62iqBH3H2hgcH6XA19ZQmMvAMjtLzG42TeIUgqpD5DkTNw87H/Ew9oI2cPmXRYohtXgc1V9
1zr4rFioaiw6l6zcOKbq09AxnVK3yywn7mneXLhbMOwNTDx+wBWwa+AYUhlldvyB0HzKXSCPOQ7D
uZGe48TX74GTfLOhMWZL6bbKRLlPQk3NiYWFP+JdzeIDIDD6a+i3GmMoLuy4DPXZxBx+gl99hrbs
0F9dIzWo9xNTRegG3xc1dMvPvPhMNSxFEC7i3s9rkE9xdo12BtF4PVjd9wQxTUJRoUJHz24ou9mY
eJWJi+rTl/o3uBnut9G/Up7EwPsNAYAl3ih6ufdPbT01ia8ISUCLAAK5xx9o0A5nkTcInPY6W/DF
KTplQIVDtVOQ7KpThwAq2siTk4yvB/pTW4OnrVbkewhd7kf3cxbRIf0l12t4gTFWOG3BqAYRSK7K
C2YPmAfRMwbpzvwrfuLMfK8wm2ahUaO9y/uTkDdGks83F5783d4KFtLvVOZp9TV04G5x2NKHbyvu
ihDvIRyFi0BsJF3DyR9N3LVZdsCOF4pf9daGEVqLyMwX/j0YIw3pMQ67zwWxS1UL+F6wWvHcwtMi
JeYznlDaZaSPrJUQpyVK/5aMKB8eQckL1gZR7P+hsLoa8caFBOH2KAM6INXpwL3S5UfgBoIV2nAt
2bwTwU7I48gvu31chsz2kXkfLxAYF89CdsjJtPB4K77QZh7WslED99Q+tB3fVYmHfRGyPd0xlRMe
yfCxSd5pjzMvABNQWXdzLvxmNqXalmLTASPqicO8V4MV6HhrgFcNz+1cvrF7xf8pai/WDQTCjxZF
vxsDAgU2VQJa1mRJ8zlvKOj8CD+TC1ZfGK6ppgk4GTfe2+xh0xm+L3/VcKNWE78aGz4dl+ZpSebC
lrCObY1jfb+19gqsuQcx5aH6lYyadKT48VJLVZKsrtI+wbPEhyo//pKFxuEZVSaW9BH2frrWickC
TvFjLCK4sfui/sM/vyJGUnofYIPrwk0WiubV6qAMi1acIonbxRvk2HxI19JQoKkghZQYtxrgiPSg
F/o8oRL2hTl93RSBYAqrDEAf3iSwsu3OSucIFrM3PHB09vBqjL0MToOikhPRdLSnyQyQY3m9nECO
2QMV7RU+2yZ7x9w8fCOfseGDhNZufiuKZY3X7LFgeW4U6DxyUjSthnwsxzOhYSzRAC6s42b+8VUb
OkGDYk/elOfRvR/NQa96HOzySdlgb9COQYkCB0XYjt1L0c+ndlPRrpJOh03SB5uoh1eJiAXFQc8x
PtPFWpuBOiohPmlT5D+XShXFS54/q6xEGxIxG+TXoz7e7HJ82DGj9muzSvXjVtaVUFOOn4F2VF5C
jcL4ycZtPpUrTiaVcoXWqEZSHu2ekSHpdbgEWV8/mqnB+a6O3fKUOYGiCp1AsWmD+5Duk9AdU5RD
a3wyxOZi9JOkfUIF/Lf8WDpHaCzmSPTfwbeXRSKjZLykQNsMBrrv5qKSnQCJhkpHfMJ1J8m7oFUk
RAGnySYIsnoC/4RmzxVgDFhp9nhunyZiqLvrT0Xz9RJzPexM/bmS20O54qtC2UtsCwZs+F7beHNi
A9Mzd2k2lIff1emDScsqymequjBh9M6tFYFbD0LvI2WguCubs3gSfHT62HiA9uZfPvCOagiVLj34
LZElWeVr0wGbcw/Gj6fTusPH3KUWdIbIFxvHsx+qlVbVNcBFCFj0PNmzgsGmOHDgtnT6hn912NWt
EgCcMwcKpSLWsb/FhuSzzza4qVeVJa8G1IYrHuJxIZdwjcO0M6E9lvs5ayBSDEYZVbVW7xyVncyW
UpUZ0zeP71NgOCpPzfmRxNgs7BK0Qirjwsw4pmhRhEhEXSbxlKL+eKsK/NLwyhHmu5CVv88b5Sra
uLEzGxtNPeI4nZPDC9ZWgL9+ZkMfsxOvDcYjrVY1GthvP6Q/ahRF5fJc8QZc9DpA0m7KHr4lPLWe
gRP9fbG6MrFCc2uWlGqWuZXMdN1kEWdh9jAIG+wW0nsCSYzj2XlmuTaQeTOgAFyRQAW0QoDfOnV/
o5pWILel9+54Sgb2hOrJq5SazIeYB/ll1NqTTtUlegnvVQbPirN4AGkTKAirhqfxXOKQTOPUERub
L7keyb77aOXEygIbTvGt5g+ttHdKQC5j9HWoWgI3Apt9uDTT5IrzxVhfVrMfJqSqNad4EmRCq95g
RwqJnhTxd6SkRCNOdfqmS1IlwjdsvnN0Ebx4iJb4o//FzR8ikuwhCWgmBNrGpidLhM6v7HHkxgxS
HhdWT480yaUtR43hvqSlRgFkX33yvZf/gfg5cVclFaUpA3X13JAwAlfCKPfTFDsfbpbMMDqXKyhG
Ts1xYnwwI1cIMcZmGQ5cjO7oA8OlJ7AcQjTZ97Y1qrjQkzU29nEN3fWFvzNLGOaJ78Gb5ZZG2slz
lnZn7Q7fjxzAsUEwK7A61MMy3faTjX/NGhh9si6xfbLKaxnByKepTiHt8jxZW3vyoF0XBtXHX5T7
eAofEjwIJCmMC/dbz7Sqkqlt5vOAFvlDoUZNdUj8sSiTbLYIs9VGp65hp7tuJ+TZoSkZ8QoQ/uXU
wVEhs3yL4e+QKnRiVGIdISziOiLfC7uykRlhelasPJGOhG0V/+ncOUnCWG4cqp2dfEP7yCTs9G0o
3Y4nJUPiC2GwMUnM2OQ8BKns66v5ZVswi6zwC+WXJG18AU7SOXmW6jJIbmqGALqL4n+B0WBKzXy8
B352blR8R3dco+Ce2jj+agMMMEAgsox9T6zJwdjoRG2oH4i+hhTi4wLdiuxm15R5b1DNKs2t7i/X
XlOOiozFthiqBiuErXlaPIzqracBD64njd9Pan/mknK6TTz1myW6ZxVhRqnEvxuc1tUblBAnABg6
wPD7ESZFgiwBanDE9/1myitJBb+EPOrFa7Gx3FBWMf86KTjp2IBHjVfJcD33sMfDeMuvupWsn0yn
eXGlsTXB61PYHe3eb9qXRrGYydGYN1K4RNmVW+Sc8QSplHWMc8anMVa+Q/3TIAXXun/fWlJ1URxm
x2wiW3e5tnibC51VDsXtbV6meD3ALV8PU60vQ282aQcYHN6CMPw4NhRS62wdp0g/3oDuAzFLA0mB
yCdnlKSDSA9907HzobLnos5toaWwmH6Tts1RBf4dUrXUXTBYSpRiKakbRlxFE0fpcJnw0wf2b/Zg
WFUEzBFQxqq6LmD+nAphCbnS/xS+GIXfwLD6PhqH/2p7iB910MSU2ZLBJWRYyTthDReIRiy/H5U+
jAhSig8+cnMSXOvZjQDFkNPGd3N3vBYyJ9lF8zQMpUyH0kK4tfkrOucYvZfs5jqCnAagieJ7IwDx
fjgtDUCxuaLKbQHFURHCY/vjQ2PhtKSPA2AjbV+fWYkQTpX7lypnEQvXvKXWBCGSnbYlNxtMAH9R
YoKf9nq8XSvxuP+yKh7XwtMJHfHwviBt0FcRVkFbxX5FyQGbJlvv30SqztogIrilSsUo51nEVwnN
IE0C/MJ4lJqWNtIx+yMZgwqAUK2V812mIcCA/i1ZChsnJM+9+Tpg2Jg4DOPosjRznf3t4TgoenoF
Qo9HOREXtZD6z6crbph/v8uaD4k8K9d8PwXAEngoSB6LXWcuBvma66yfnqdqYAlJA0pnJu/skIs/
ZTmi4JR929uNJO/D0NpINDQgcnYQ7F9QyXEPVlA8pgoHQvBzCNGVwb9DuhT+46iAdXnCht+MuA9d
//sZbI4LR+vXZNjraGR0l5Pvb7YV2r04qZURc267OHYdU2pdx/WAaWEKVnJbz/NcJUTmRxvGcxRa
Nnd8T11+EqzXQl5NR4fqzkBTfgzK0tXqUoy9SQEZ+K590lVxWOPxLXbfud+szfyjfdpiXaE09s0m
WaSEVPxeCsofEqV0mzmsq3xDGEZW/i7fnH1NgC8puztXepubai9qWOOCXu0yboXDFzq6yTNhm9M9
lUxeLj8C6wdvk3fo2NLAE5ur/FaC72Cs7RQymZBlSzec7W2UWPiOZudVlROepIzBqbwvEoz8/NB4
zbVNbqSIOhhj9qZlpyYEu/lN/tIrzulHlTXmUL/LrBFEMxWIH1EiZwFzUM+sywPzQ+XgOilCpzK6
xHJtXwhe8203j6ULtaI9BFaLBallQ6mrQ8vE/HbvRxZep6UZFb70H/efTN8Yms1B9oXLCU+14W9I
2lS9hQir/ZsWq5lbyxHJ55bgKNDc8Rp4jk2EqWlTBLt1ZAkq9QmNnDZ1xVL7bmWmTf7W9EcNqv5b
I/1Aiss24266Ai6idN5HO1LsPQBdtv4GHKRi1sqO3pJOURekZTHPSxDSL4xSo6CKbq9BffMtDIo/
JYv5Ysjatg0PJKXXU9pTcFd1FIdPRIxbjrtEWrhbT0wQtmQpNSxpkXBGaSLOROfiP5TjLOzNp6Y6
jSMxgzZ3yIXSVo/cbMU0iEchUlyC4GTWBgmZko4uGfLp+8e3JC/8Qo3PEfo+bDLMHyGJ6oVl1hZe
sQZwFUBuZDJPQMhraRSgoCGB5X90BdO6GYTEAfxdNjqv7Txmm3cT+hVTjVPzZwF7qLUCIH9qfiH4
DNUrEbaOhCjgqTw5Z2zmq9rIpkFWFsP0yxw+UPnw4vDVmh7KTzQHXIJK6N4bT9pb05lK1vX4WuCA
DjHFoytAUXntZva79dE+TZwX87N+V1X1QfRBxV7cyHfkcLW18TH+z4BkgrjoRs4r9XOWIalK3GKu
gxxQgizN89jQ2AmGJGk2mEsmCgIH1vPW03VhWCuHoCRWF15Pnm0THgcHBY1AyoIu4+CaUUjIShas
gIvBAaP90uLn3KyCSqre6+8Y2DgTiQYqDTM0SSgORkOf6A/YT9WVKIntValsUpBnprFEFu+PJieg
8qIlPFSBLGQK48fh3mVXMPlRflDeAnV0RzEUa50E15jYa2XP9QatBlGi7Tb2Z9XbRa/6PtOvThof
YP43VbrHBfQQRdnXXgquyHAV8wj/5YS1C13KNrG5Hxw0/aowIWdWAa/UgLGC1BbRYTz7h6u9JZOo
PyGFTFDNjeyyMEHZok80UL9CU0m9WvBOG1NQjd8RgKcWT3s0jXNs2OXmL5GZOWud5KPw9SXCrlXr
FBn9y2y0gxczVL4RJucvlPN9nq/B4PoyLU9r9B9CxA6O1VURfeKKieJQgVgsRtJI+Fp/truennsA
83V9YsAaqCfHnIA+nO/6S+qPkU8/5NzKN2+Vh3ZW95E1BR+2nfnHLEjHtyJbf8oigz1k2ygoyhkS
tGEwk6D3ybhZKA9t4hTx//5JFmdb4O8R4CkokJ8H68QOaptAloHnXVet4fq+0NKawYM4wIa6Z74h
yhCf1pHpV2btReEpR0nkZGy9eNvRBJhIArY+XjucLQj79o56I72FEfofb029CvqtSnPPVJ2kwwL0
4h7Z7sypuMNF5GbQKtsLggQBLqh4U0BlVuqk11mjkk9lqzchk0slYNfwfSmqqL+28TTGrBaIu2H7
q1x8wf+6g3jBLANdVywIKnNC1/oly/mXtqmf0hwXc9B6JIfaEszbHYgrhErYSVzUIkHzTEfp2QRs
VcHMWeTYfWwTf54B3oxdUwPAUkLk8OmMYTCcciEo1fERxEIKB0h7NpB8oHP2DcJyg64YpTgufveU
F34vK1MNNLjMzWx6MmxgmUCQNRTM0AVNQXg/PSNiOxT+nQBdttdH4U2qGB+MjY+J/GZwdjjCve5o
p9V2NKViMxJdCbA56nq3NNkz6DS63cc8AdTTT0Vsp9eP9N76cMpyHCZ4JKszpOfHGKnqM3F9Mp5S
eI3Lh1zvrh3cGcaZmkbzpawCwnGLcYy4+ciLL0flPd59pmKPTzzYSLDYQxU5kl8Y/b8zqZP0Ty/x
SS4yl4Ra34tFGR4aKeFa5EWh1co4CDmei6oCTCXEAlPJoSnEjc2vhk/iwNdOeze+qup9+s9jxfTZ
l54hZTBeNbityaiPFLVJntNoptrTxDocwVK5C//pOMFWo5CzciDT7r4RQ0r2Dif3zcXRWfZiBOl7
EbsDKNRpzO3IpuGn8BPJAkox/puZHzkQi9dxQt1MrIpJ/ReQlYEcMBLemyO2WvG5syj/Yz6o5/np
cU/oFGRzozmhuy0QhTlkm1jB60qC98yFnIHgO+iY2n5WBoWHHbXIwqfybX7by2FIIUiQTBaeoox3
tx0SfE8UnYKGmqhxb3Glnu+iP1QT2aAEq2xAZ2tudKnXDxAtznP28zMv8Z/ktU80dIp2CO2zB0LV
On86q34UwuguQmz0N6iG4hvtXZxopeFC6Ey3imkV7oHi5RY3ilNg01LJrlCJoA2qZRrsopK7JB3R
MbAR57hZuIPy3pThDldhBz8vsyCVrHtEVLYwJTMVpqrXf82x8WPR0tC0UbgMckmKP0F5GOoak5wV
MjYkfMb/PhuYTNnGyJhEDAdS+SOkUOzi851YDMh5PgAj0PB3PxafOU/t3BFCIxCGvHx48vpDRUAP
pWI9ZOlhvVxHq24mngnr0NUzOKscCFA0bXYqB2dF/iBkJAPDoSlzYBt6r+Zy4p3iwrd25b2Q0TSt
04SNL9iCHwfPDN9Ak0oQCq6V51NTk5hdEA4Lg0mGgSKO0Xhs50eh5XLf3yZFzk9ewXWIvdqk1Ymo
QeskS7B2xtohdB3a9ha5GiiYwyyyKxSywsJ8vsy1Ig6gCMUa+C9FDwgjp4Fc77g0lsVulBto1jg0
WGgFaVI+78IOslKPIsmBwLRvDVViAycvyE3HiqHGtkUsaKxHlG85CdS5TaIJ/v4jpkX68i0ZVFbz
FVMHY1AWrrCrxjChKO+Urpol6qkqKu241D0JUhx+6JhtdqVRD8Go/vwyX/RHPF6SbIVae37Pcwre
vVo2WrtZWS98hDWJeMs3776JzWtKcQA6rMYGD9gRqswgarIjClzNE5TKJazkUFj661+TKg2itZEV
tulqbNYxqhXI8COXvMz0INKn3oJCAjYRx75RyJb+E0HWA2VfDH9HFIbZVef5LSBWat2H3HXUlUm9
MYaVN1V4/WJ74G/njVdoFiyeqqq8OswajRUvryfLnkiZHgeQkaKliHzKwVjA8dTQ0t2p9/CSYD4T
CQyrshMEIx6Q7shF+8aaGLyNwcF0u6ot9MvNKdcKEhP36c+r0mEyXE6Ep7G0+8jpiqLaOKmNW0iB
EbAwyQ6aWS99YKehWrcQGsaYGBKv66/n2+lgBXJpwZOaxPQl1QLaJOFuHXtC9JVNHekBN1i5TByN
pZVyaxicUpgYwl1fR6hrm8OcHQ35PfxZD8QTrA3qVwIy8z/bqrk4fqnOSlcWAwWGf/MXekjj3Dvk
Ux+6I1YvRfgtvp81aWFYhoCzCsuZ2D6EkA4vl9UL1Aja0vVq8h2bR0maHp8GhazYi9Zbo85+HNAq
IXPtjo1Y5vW8RlJCF8fHAdIAYmRluBgPXIZygEexl0qNuDVuQfUb3P3TJJEZJ/xJQeliKSz1Vh/x
kleg8/Nsf16+pc8Huxo/15an12TUIZXBFfMtOw3ZiR5YgMfuTE68FznByvvCAhCmFqwKU3zL7GD/
8qSg840pJ46JvyoiG0UooddV8qpMRdrJLPhsG+RHicidKMX04BaPYpEXxK4dHd9bpaDZkYpgJuKJ
Tv4i8wtLBjsU5lJ6uApvcooHGzme3vJ7emNgqhYgpjhy4vIdaGJgAf6JBtirwIfmYbCVfkHWov/4
lLWv4D6KLduIDeW8WHeIJWvqDEOOzRNrqv/iDSjTxsicNh42JJO/r+pR+FfRYtsFcUQkumYt4OnQ
t6Vn22t1mShR0th/yibH1rEsbC0mztxoJmeVYLcQ2TGILNYW6KcCdeB2kEVhOqXzYDwwG1UawRh6
5K+fU3cqZ9uDhVtM+hoGIL9RXIOHkYnG9Pbj9+X+PrwqNXCn1HT3VcZdxG3sB1V/qI8gteLAzYUx
hX50v19mBO7hFTLkQv8pCyeepnbuDOdgHCEqL8CE7xXkq5kOksRmZk1LHlbG9HKuGHF13LAa+BMW
VJSo7RO8kNPh143sgm+tBavFyOd9FB6prri8LpbcZkjl+Yw9CfnB5+mtBcrcQvM8k5nwkfmuflCZ
Fn1BIDgatiNpirDNLB0cqz6r6TU9tykwZ2x1YRTMiUT/cYEjp8SAeE+aC6qDmj3VrVydvxgk6dm9
pKCww61WQh9fpTNmODcwRtBCoEvhUSzfxUV3tVhP+SEIEBpHMonC/DwnW+sHFO9w460i5PqLY6r2
5DTH9JQQfikZEMyZhkBg2rTInRVLNQDmN71R56E9OcT2UYyd8Gik2NKBXmV0/Y1xnf+G98Tiu0DW
D0dnwWWGKe2NNsOq7Hjx5xybXI5AFswuR6niliou546IRG8fLRDb3xvkiQoZr5AKpKS256XiMm1Z
5H/8/2g+crzmUPdpDAwKoQXbr2WXgFVx+zxPeZ4Pclpcb7i//VRyWJmmOS0hXlZt/QWxg+S/Ce81
DgaDAHmMeEJ9Rg3G5WrptXXrzvQJHyeQsRbZvzFjk5MMBfoCBByoW9Hk3EKUov6KAzYiSR7aFyYz
9HgvklnMQVkGhR77Rjap29HSPyLLJwYJDh8T7GPgp1CepYFSXbQ2XEF1xFFk24n2+64c213+AUZt
0Up5UFgVRRaKnqlch5GnxKtIS4Mtnx547CoSaAl1oZo/fUnXRP2XgpVMhCNUhCLV2rz1qf1cfxq5
cdK7BR5kck0CqLQH0xGUUaXVqsoiVzoZW1nfkdqTGfbI1cLlWCUIQ4qRYn6U/MbgSrlvMfj1YMXq
lkyslr9AcIycLo4HrdRivMnJr4YZTQMp6ZDxGYJE9BpLGx8crZh2/XqzWLG4AfqTAIc7r3ptv203
yprqG9xWckH9Bd1JxX8Jk5BMy/zTr5V6oIB2IvXYNMknd1UvTyV7nADnaQLTsPCWEHz9fY/qK7Gi
RMRe5+fzfrKJYmDuMZuuYkFQ9FRuxv7eoXDXkfKT3GpQ0049JCgtRnLPHULR64Iaqt2Vkf2sEzlu
AJKS0LYbDcaXdfcTkQA1z5zXs6NnvFDg7K3qpAvEG+edBG28+6SeAQ1IIAncyMHRkIkEWmyplAxG
W8y75H7QJIYV3sY44OiZX+bX7+NyZ7DL2LjilSsL6QdQjQFuljrkwfpFbhxasbZQ1qIQF2eb9OVb
CWpQ9sxPmJtoHfdMqIwlxfIPC0BlyYhTGLv4J3T17wPdoTGVi5hzshIJnIbPaRcv29wNMmZNcuxo
I5TvduDlYA0sM7rO0OOZDsZrVEXXXa2fdUvTbQaZqCkM5UV/KPJxu165axVA0cHF+2QKXSS+w2s4
3PGf4J3i1u83/SqTj0DDzDh58RtRxvAWE4Ua5i/Py+ZJv200qYbrsKFudJlGRRKjgL3fpOO/i1ix
fVnbxgXSEvzE68SoMG/rpuWzb0Yg0oNQsS8+s4iimV0/NEze+x1wf450fOehwi216McxzhxMI6AS
Vrf+lD9jcWUJXeXuYjzt+qbk9OfMEhRyrQq1AjBwCn00ncsLMDUbmUTVX7zzFJ6IEef8pvEbI7LO
EU7XqrEz6LS3vohtQxaECLj/Ses8tHXvcM5VAg0y/rnP2o2hNFqnt0yicgtmrT+gGoEIZrnLVuw1
LU2p4bfpF4UTp2t59NKqr+/fJo31bQXRavCECerELxSS47oUtsXHwZxsSgT3VpVW1M4F8vL/am7P
LrQSyBPpbqti1/SIlnF6GpM4BfVT34g38OPZ3W7f3lzp0zegOz6jrlH508zsNjO3wrYO0K9uB6Mk
FyGPJ/qHlISodzpGvJYOarb06dCQlsb0I665uLpPG4Y99kUhZHhWp9DyN5GGUfU5TjMeNNtCnVCr
xUGOYVk2sv5hsUMKJ1Pkk3qyMvTyvZXwNwI7nHbdY6S4tbx+pCHS4D1Fs9L1WHCndr2d8bm7OC14
9hpvwfX1Y6jiSL+WiSTBm5ha9GQyIuSbEaMDSPbsm5kL+jiMXruiAsf2t1EVYL6h7vevTTobnttd
DhaEeNrZoM7XT6zyvsH8fbjumiZUWIxqDEL1KdrDO7Khuq7V20uClauDetnVMziEifk8dpyvzkZX
koiWTBIG+ILYPvat1+oe5J39K9kODbdwVuNNaABwZrP9rEaguE3NUjSeLYiohhUcQM41BGKxRrp0
lHXFOqxBt9C45yVTKKelmfniTR342S3E+sLOrKFSatPlkWZnsDH4CmgpRxRw6Vp1RSxavdZswUII
R/c7STPNw7wem5ciy0U53BzwlOGRIrF3cIebYaQxt+p1Kjmiicwk/FNQZEceuEuDmpSstOtW3nO0
7OkRcugSn1eNTPx8zs2T9ulDM6SlFJyJcFtyQu92k0y8oFtX1cJZxtpPt1kxaWDkTGfN0t6TwxYT
FjkGlYHS80rHa7QWiWcijtTLOV2BYVACp5Fa1qgGxjmhHWXfbG0PJ+UnZbQ+Wi86qO44n9euhpC3
OtfpMbJuTWHd4uIqmEjDCG6WkwAL+cBhtE80ucq8COuBjJzcpYMH2WqBSYDeKcmNC+q80y7srBlb
y+Lr42WnBGyMPwzKnbmhXOKMCsx0/86Pwqu+Ha018ph4OBmBxdoQQabNI8wfywqJquDIybd50/FI
utOr8P+sfb+OxXzZptGxbC74xQAEviTFF2zkXgsDYiuIRNQhzcXfEj3WPJMt6HhCiSb1wASA7vVL
97ls6/Xuq8cCSO4gx2zTBgaYxH1Xp6qRb6mzWlyf2YdMb9NiOTGt9JMWMeI/tAQvO+ncjGTIudsN
FkXg7H8qcjTFsgjhjVABeiZQWJnwAgex34oDAwlMimHKCmdy/wChGMXE3S9D5BDH4QLNIjzGK+yW
AaHA6UbjFsEI+VLXcntG7LjYMq4GoSGy3funV9zQwcluw9lQ2nmn3cGWgHNqBvrBkT+vscTMaAEX
5un6pA1pHzggT3licYiSpeZdWDh9bry1p8veQrKEgiz+MKmeJztakDTibu7SzbedPd+1KdcqiAC+
bXzaoivJgKWPO0On59RAuxkG00bQBFQvo6U3FQwkTAgRZXMFbI73Xrknfebr91mKPpF9xmMHL0c3
osLzbRwX0mAzL3wHlfw3eoxBitk0FYc63j1207EUvawfFd6/aEQlY7pjcZdlnipVW4a6ej1YVJIS
yQVTsoa6qc8yKkqktRGsLuPAZmmpE53xrHvLY6oX62pzuC5eCHNC7dGW4sRPIOLckGO+1m52hTYo
OTkCBM0esCXzYi6DVCRq3lmT80Xtgf3Wcu1CTVX1RtzwRnaTWj+WxhLDJpAxSOTftfV62E6N886m
W4HJ2pZsDjpW0vZ9Zty8LogLqSYez4blKpGlgNGC69pQWPlrLQG4FR8/3DN7yfGR5Mb40P1Hh5gE
jkXXoGB1igBwLragKzyK+LCQniD2JgwACKP9gdwF7Rqt98Oguvwr9l97I3cn18RwjE71/18hBG1z
TsOLAolMxBTq1HXLdc62j3EvWSVV5Cw7RDf5u4uDfJnWUqGOrhdAqrGjjld7A/uV9UdHMs9W302u
Qja0rmtKSxrGh5Hb2fFV/QBjZQsSXJUy09k88FwqxU+zEUzsx4g9y5SuYlML68mmHYDqzAsSZWNo
LSuFM1faPeQvWq2H9WbgcQvcu05SmrLpdLwwxcHegidtNt1uTLx/1yIm4aXESJ+N+wJX8dorFVoo
kZD2Oqm3WVuHcS7gnQh6bdaOPAuIrqMTvXg/OhwHayopDf93Ff42k5l9LHcaoNefZA4frZJsBTxq
m71Yu7fK8aisqa7g0TJjZOjByWgqx3z0eUH/L7vBioA47jxVfwmprW0GZSH94xf+vMoT0B3W8iqw
pDOylT3OM/K7lx21m+beaAVcJZ8/K/UciXwhIf8lpXJfsYMcWgWzjo4T7NrOFRXQ/+QzlNLK9SAR
/aesWV9sbJlYmRb/SAv52nN7cRehnsi25sy3aeCZ0JDPCEoBXjnslnfBXXO4jBudLO8UgIdpIy0t
YYh9UehW4kXe8rLy9jcTKMnW5sFSBktYfS6waq+QnDVFSOqJKlqtmw4tDp3kywUlGyT2gZrX9NKq
+itzu79NHUoAr+Ej9PA8k2dxyF74E2zlV9p3AeIB1dENwFFmxAFVlRAxxSnwaqNKKCxukYDKp276
GykNV/7zWxCBi0A3QcVltLc06qA6aCDcGzuLZ7AlqdjPMgfP/FdxzFcJhOGjfd2TKMJk6WvTfH0i
HwsijjoKynz8MGgWOriDwhqu3jbzEuYY5IfHJQB0N5bjk/VweoayXxp8CD9uqXVBAglfyaQG7XLK
ae0JYmeNNuUx0b9B3MlIrEYn31WorqeNaj67WwQ2IaZq1K0XoUOkDQFJf6f7ckRidIKMXbPfjCSM
yRkJGvHo38VSzdVowAyizKvKtLNsdqfED//n7UqJJ1wYFgSh5MWzQ1YsK5SZnU+1EXFa58VL1Ceb
uV9WlSUVDcoVUL/IVaWJBVSlhfTmezVAs9c/QGMsvPOoIO0YlVpwuzr8ubO1EnDKp6frN/7QHS6T
WVSLqZoSKzSPwBz/CuTHwZ8oT2XVtUnsSqLQS81lT/HAS4UBrmkEIWbvUYIIvGczTY894tMWISXd
kfLh48cwpQI2kcUJpsRVfd2uka5xsbI5QJu8ncYs98Sz+dXO/LBSKNbu+YiaVfdArH2nj4T6BmAj
6/Q7A6qBNCjgYAhnQb8LdBOnAHV+dihH3qF7Jkh76ycA0t3eUMPZnt/OL2mfV0NbQviBakRm63x0
qz7szgoOW70MnHG/WAx5zZ2O5cDmN1zyxuJcn0wSCbNA0RsUZd+xWz1WihXtmQnTC12+t8m5Eane
+j1279rBtoy0cp50l1pC7TOhyZhEdfet3+bs+DunTUFJbVdXvFmfAQEc8VGtZaDvKVqcr47VNjkN
9eJpCSJV6NwuLMShNbPnPobb3GvDP5z/pH/uOC6LXfNmAXIhKlNvBriRu9zNdSMMSUYXsLkVr925
wEXBjflL8qIg3GsVv/3uUnhRcVGsk1MzKEFK9Dz0BykKCH/txAtAoUqmQ+LdIwl0ktsHXLTkqlom
QY1aVrflX0k4tKNpWjooXUGMGNwSm6m06i/Gec1s4QaYgHtywfHAwjmCpcQE20uoheVJB2sxuy0A
v7ODJ8cOsZFrcGEfCloX5Qyyoqb15ff9L74D/hN2OEfQGoTfhuq+bFcV3mT8OAwtCnpK0+4sf9Qn
TSQGZ7Jh+rqufTUBc+AP7gHUvguSUD/ulauwDgeMvu5RFikFJUpGmOJg28X/foQZ+WQEAvUApukC
lC0JHmAPOteURuExqqdDtZqSyHqXVfHwe3mkjOiGHAiGg+lsruNanbqQb1Y5JmP1Bjs5DTr0VQ1h
Ab356bUCyo13SEMLqzMp25DvL4aKP2daBtXqL+Za48+vq9CJLEBIMk2beQc/h2jD3JYn2so/uA1e
3ihmHPrlIfR7WGs/gycALtCqUpuo1/gjs4zcT6mdWMJuX/M/cL/XcrGKD6bosaE77Z8TNLMFXVG6
FHJSf2oVU/4NIdsrr3mZGv0v3HB+qXdqGlnh78q9bpHWCTLG2VG31Xa2FG1/hIg1uE4mRuaJ5Q0+
b9/gZUnu4otmwqFdhGXMwP+4uU64NyZW8fugn7J+0w/ZmhKTXOxxsLr8JbNKFFB9UOJVXN6whiJ3
sdLji0O5NprGBM1gooMh5yA/JGZRUqkkeg9oSKoyy1MAQZAqZ65ugMuS8c68wUqTktulsoOZ2ZWt
MVCQfF111OvxLOnF+/tBrawnnoHSWBVC+UIBSzeQmeaaV7g2zxY0rWwrhoXwqWfvSHzUWZZIMxn1
RAqMj7n74JnpGJSDYHI78UAcdMqxtsLn1UsTYzRvZMW62hqrFvfLiSmAaU5H46aMhKVSvRnPE3V1
HExr6X98Cz/HHM304YJSCAOOqLSVJKAfPsytQgNzGfkDOwTGTpht0R9EIcOIhUY8/O5+ViK4gjYI
Zli0ugGGnKZ12dLzKVL0fUoDsi4QuC2Sgt73w3trZ43CGB4PQV5TrZfYwvrIAoo9dFZPZO7d4pon
YMe91YIGdTfmGRRW9d2cVHT9Bc6aCkseon05foCElWRiivQktxrk3c+JmEFy9T8uUCEV3Vo5VpRx
w1yhPA7+zm0QtAFqSVRhlgjhomLVilhlkaclbfxNyVIVPnd+VwIFURL8mO1Klt7mY44UtfpSzLyR
waKhKRxiihqRYERew+UY+qeX6tb7mWQIb3bFSjTe4KJFhL7qlwZIm5jAt+UCDpyGGrFXqFY+bXeP
SYqN+SVvw0/HbZi8nzCOlSK1X39rZGOulwU8/4pph8dQhYLDXXRbaqwwYB/yarc/XNf0J3kI6riU
EgdN6YGDusaXFr/2q69hPrnf9xOTY4tuNxwefH/Ldt4mUdvWOD1stYvN7S5wTmMEBZVhgsFLrwOz
7MrEIg6JrUgJC//Anq4uCtkTicqJhZGVi7TkspL2ucB4e5YqA00w8pJ6Osvmg4ISZcqRZN68DApN
5QCKVcHaMevDmQK42aAL8fNncOijNHJu7HQcOwUCrkWpixnsWpU9W3WligqXbadog+XdO17CS824
J8xR3+mHQ3DD9PD8vALgAYtA9WTWbS4XMFBYv/7bmCMW/E9K7tdEixD2vWj+Yg+LISwUm45XgjfE
y03aa7rBeIn/zUazsB+0qOsZheffJSt+EuZY4mcfM80ikQZWq2edrdI21IEYbUo/6XN+FCjWymTK
liELIT9Yd9pMjR42cqLA+XwsgUdX2Jz4iNp2E27TdlybrN8d2B4SSJs1bPMokQOXPzBSnRDrqCx1
YIZvqh7z+8SIXUer/Pfm+1MzaqvBcnrWwG7SelPbt/wROrSPi3ni4rjvaZNF+xIpFGAO5qhiY5Uq
WmJcA/rpS1xQitSKGp1SpJdQA2ZR21ZGeG+2o25Xi7RtDAs/JuHAjPROqVhaU4vuaXhOAOJTH7tG
ym+iMRZe7s4wRt4GPNasQgzHSLrGbpmHSFiK1Um5hVrKs9VVYDk5ubFIRWqFvgYYEvuln1EA77CX
fYwLw3vpxb+g+H4wVUkVa0Pxu6wEbo1yYY3MYWQOSxQPR0ocSTy3EulUTjwBrm8dQL/lNnhVASN+
QpNlpU3w6uVNyX3cIDHI5Yv2i4N5OBXSPvsGI2BaqduVAulv3yrVO4HKdYRMnZtR2nq4yWhP1oIr
fzPY9qGTEuSeKP1XdD4kkT8vq9S/B0tTcXdur5pnMulIKTk9I+tqMfOXL0T4RNoiV6SGL3CU1gj1
nAz0D49HkbME2J0XantLaqJuNFw56NB9r1QkooG9ZZY1WjMj4i3fSqjuLryQRWZNF5GunGZVZf6d
smXO8GimlI1yHmntL48b08kWNSdLphDkUESg/HnCqWZiQQ9hbyzbgtAU7nBbKfoZSod7DS4Gj4y3
yqa8VihdIuw7FFP43+1s1J3WNwjCWZPWced9laYNnngdtjVEGrPNCI9XudEh1mV9xw1fjr+2MtrY
ET/SkUpk/beu//hA5xo0+z7S1vdwT1mA1TWk3c/lFMqunsKtEF7FQeGH/Sj9BxtP4NN8QX37CW3H
Go0q+PFZK2gfpnaqMlD5ctUphKuibiVmrApj+/aD02Ouvp8s0OY1lWSte0xTIGwmgW+B+XJlnXEe
a9afJYxzuX7a1hS35e28nCt4LaJZRMPkcTr9ywpmkcLgjI9AL/XmZ9g12edvA9Y66GGvrI/UXd0I
VnjbBY8lDK06oQYSQsxN2E22hj1c4UbQx12gu6rjPluBaVjK4d/5F47c1zZnGrpL75ocRfF6z6KA
Y4P1RkVXjt3D2SfzuC4yxvKoI9Yc5N1NzC6UV+aczjinsskZaMDN0jNN9y8winvTeExIprp50rRu
YDQIoZaTIN0NjOI76Hz1FWjcK+1Ou/vNTj+3GyhETIehRVv32Mw3e2a7JNw/xvZCA1O8Bw1lWI35
kFlwKDH9jUcQAQX27niOVDswKV2h2v81r8yd/GkaBpZgpZC0K3jkZt3vH9k4e4RgwMpk6krmNG0g
3arafgqJ+F+EOZ1wcXyYW1hrjLnQysyZEdoOohy4OQVeeuEExEkZJT1eWr1wvkSuZTvg0OPkWO5r
XpSUYIx/iNaQWMCt/TySaFr9Ni96tqI93NZ0zirsYHOEqvpSzb3N43GNwiFQYS3K2BcGzsYoW4iB
l4UwTd94it0d2vHE10cPpEdJgZs6okVew2qLaQYRTi0q2NUJQ4UZc4MolHr1aJqHb79WTqqxI/Fz
Q3jF+WmUTo6zXH/LYo/dNgPpFIO4M3ylccOXzyWvKG4xWQjhpG1cTvaHkZjWQe5skYG+S2AeQh5/
r3pj8CJIJCVzroZln15pq9iMk5QpAw9liDuiDHO/nzqV3mCiu5bWrEXjYZceuArocniuXzrm5smk
XcVbuF3LXt/CihICwQoFfPzWoezWpuWwbx8lWqVJAZ7wfVcVQTopjQ78z5FKcZ+bmr0Eck+7qX/n
0sr7MLbQoo807VyVmkgBr0a7SErBOnSQVs6jQ70+WS9Nv5XiFyAPGkRJU1t3pcwDkYSmLi+weQLV
MLQI6tNAmRJ+qHGVDRQOc48K3bHzjqBP0zbV/na8js2DQ+V/NVOSvB2BmfB7WiJkH7Wx51+ngnNV
UctUAtv2CxSsXTNdza1soXDNRXab4GLUg+2CDRAFv1Mg2obv1NGx0N6tCv/KmvXKznmHZkGRxW47
yo4On93HRIMnyo8nlau/7JBZGcSR7SrNTmTl14HA9Je8Hk9OpGCqudEiTB5+Wc7YXs2hx75ERHMP
emoEmOCHMtVTcSl8Mi5AKgk1yQBbk8KP85Lf4m0S4MbILdwZTdHLMamlZnGmxXXkI22TAvjZm7Va
WcO9vnB2lB2pLM6hVuiy9rN8hoLu+CmIWFXBMhYOCoFf5dg+dp76ViuFcPfWH2PAQrBeKnZ0xO/N
z3EIGAFThiHN8ltiEr8dssjRumZfC7HpRtSXxxqSAicCxneyCtlPcQCxPdx4cexDsxxZPHePPtyf
+A4YeNLHVMHRvf9BAe6fR1qiFoNcglbkk4LeZqoenOfGo7cM+mcAtKEVcPwX+RqeWo9zT/wlDOAf
hSngzjN9a8AKRzacQt9qriWyW7Phy3/SrPLsVR7i1txqMrvi0HCX9zfw1LUghhrIQsucUd5jjq5e
N2JV+HTjGsYtXxNto9sikJr3NR4mtEDUV2UowNgLQusFveYxCT0ulK5lMTmzeR9DkZ0SMBYPQ1Bx
HSPeZ4PJpB/T0wRdQHNB3riBPAV5jFcbnqbXAMJXNRQyQzZpd2WJn+qI6UQ5DKo2dYNvgDDqi/tW
bJcLwkOJpHmz+ZFRHcTXfJE8pn+PJpt4MkoKnhlXhKMNS5haUNOkzqlCDIHOI8oVnvflJtAvKHq6
7qJDvM2RF+XDWkGTE5BHEJbuob/1KP8WFpuVvcNg9cyA7FrIsnvBs3hJ+g2xckAPiSVMMVg/UVFg
n5wDJrveFwxsMnEH+WOLaPyP3JWkbpQ7NN28u/XvrJPZxkaK/SzBEgrfT3La4qr0MMV9h42eTUK3
YB5lc5aYAUEphkZqk3PfXpoIhhY1TAwnxGmw7LRMgadjjWI26SZZDjsRVznDZUmsvlzTzSyIzG40
5/3fx1dTdK7Yp11A/Qp605LM1YJF2FE0KipI7OdIl2aTjXNbBGuHz0IcGA4ymjXczCLwtIti0f6Y
W2a7bipP4tMWYYQDaEve8C8piD9Ipf93CBlDePWmwAiB5m/fUynmPUm1+eRaVOES4Latkp/GKOVj
PgmbM4TuZclgO6M48oMSzBCU/Z54oMk2s3QRzfxk/niZQoG8TYQZSylOz/YFHrGiAhJmSZxhwabg
4L3ut0dEnwmNKGLACBlKWnfQJf8WLiKKyKsyU35xyndbKISNJag9z6cdZzarqVUE4d1Hk3vmGLvE
5GLI69432k8Hrww1rAQ51b8qaw6EhB8r1zmamVplsE1soT0bdOaORJp68H9U131VI3nfwc/nx+wE
YUrRx63hTDUcps9B4hoNHfBmnYR4EarTuiWH58tqau8Z9/dZ07sWMQSI+EJiyRrul5SlMz/w58c4
dBWPvPmyyTqJNo0ZSYLDnxjy53tWoDT8nJExx8whmez8YDTzm3eakaFmWH2hDVtCMV4K1SZCP5CX
0JYDyXLOZ6A6UMi9Rgu6258HE6qHXDrjdYDLfxSSKBm8f6+DdrJvY8Ia55mrBxfYJaXzWSgwiMjA
KTUZL5ga76roSsdOOtr+nZKsE6uOxvvqmTp1PDA8oOR6HWMjc2B27fotI72R8KhR+FqFMgfESH3x
H+pRhX3cVBI7HAo8v+qhnH34rgiDiG/3iYw7mXMJ1Qbi5mqMj+4H4NEvZbbyFPQE/8xeDvyEEf4C
VCWbg8No05PVkIrOmtg4ADjTBibekgAFzs2JkV7+qFdJkhknFX11rwKV5P3AmiHqjrmCCL9IM5+k
XxuOljf5Iv3JhxdHvGkXxG3iJFy33yZOY2sVneofSTSCd/H601JhIWtfa5zC113nMI+98dQq7VAL
UwpmCauWfft/+VIiWdmau3xLK2iQCpGI8Eqc0C/pOOUztgxF1H13biOdhZNjOkEGQoszMK5nhVJ9
9eBT95/eXfXB4tc31eQz5cXyp5OI32VpU8QfRLo0DS0DHPOPEImv6Bj/J4haUc+cUHDdssV13wjx
sK09hOj6EUPu8+WMj1MI4tSXhc0laEsceDWoiS2KxGgkKZRgM/SM0JeKeXFVabSPc+vGWSjwVc80
+i4h1uyI9Tr4A2KEyDxjJAPhm5PndLeaVaC7uehvDd4kXOcGYPkyZNMVH35KMu0ibr60UiA4MfQj
5K5WeVstSMnabZUtzgv8O+Jrn8u1uBkvxFAqBGe8iafDQCYh3RiCI08+RAvKrBOyTO2NiXdBkL73
TWLScu5a/EDSV8l0dys3kzqo8Ybk81M4xutXup9hEVzSg2eb0YuGIosdu8KNDQIa0Php7J/GN4VP
Mj74bL9qf71a6+L8etkOMrjmHTD0l3+unGgQi09QiTfyJ4AqOpVAKrc/46Grdz80mAl+PUKrt6O2
r1SFipLCu83XYUmY5j3zWq+F0wR3SCv5vZJKLOR+4q+77goIXhNH2SvAnkbaxi4zItasezWOuOwY
zYJc+HmHeiRhBZvJZ4tROWRXAfgaGuRtuwey+14caueY9pNE879C78xi0sebB83kG9+p1dS5SRTD
jP3Cofop/YuMQYetiNhL5tMIuMr2AUD1PpAnoC9/iKdLRJTZibc1+G3oOqsBP78wJbRpnkewuVlC
2s3kFjHYPvkqMAIykDojLvTEWY+ogpFZd3fEr9eCOFEcix7oT/QLJ+6yHSJ6erazyPne/HxZ7FYK
wpCc32SO8wvbx+WJWzHl0wAcKi8br6PdQ6larZfaNTo1gfZ7JMgjZ/o0LhoaeHrz226gJXqX7zta
XbS67Hz+nlaWoeh9BfLxcLpp2Vqd8x6FYlVrcLZ9tJ5CL7+82vEzHKIAKB5K88QM8SAr+C6mFKW9
bSilMmwwEQOCjMIZyaVNq4OSs82Sqg1EYn7sOOwZM8q8SkGEM0zzlBUxrEt7N5cErel7pigbMtpG
o8cCJgGCVeC7OeQS57Qiucot6AYVMUDlMoFNBPGDD3iXEfactPuqLzDsKtD1GOc0Z8N/NlFrEr2r
ensKu4uMAFkUn1s9M8TNa3P/dYYhHoqXUNVLRKhRzV3+5zjtc8a5yhE2PZP4a2gPMQXi/QFHfc75
Z5BmhPwX+mzZ3G90qpzKMts2CWuphwPabCfixFEc4s+/URcxRZ9Jo2lU+Lj0BZpl5KtP0PrwL3pE
szi1EL3ayscJE/po2BjUn5/gFEtNVrgBz5bz2DjuSimhkKqNU/0X4UuigAs7wZb67+vlIsEeIwFX
U/FxJNCZA5PEDo8AHOngkVkgtjXIDTTcY1sQh+wu2QctSgTFKLKtFhY4fhHloBRlajgG2LOEmIeZ
RtraXd7hZ1xt/jjAGlSBl3hQlhLqTI2C1sy4tXZen2gOLlMb19JZ5O6ug9GHWhQVAvvg7SqoBotd
XQr31hAe7BPO/midb/c/y61EsYz9Eh1X8JJQjG/8xOfbG7CLvuJ0vH32Gbgy99zp2yU91xiS+y9O
LXR8lh5SVQYm0iQ1Tsyq/wtthOYuqnwWMGUTRhaMo5j9e5u8QiuYRgeJ4VeksyETPSqH5MxfkrAW
4j7SZi5ImH41eTBJwKgvAkBvYHLP09oVk+xf1hzGeYN1fP/vdPPJ+WPAp9tQ+0ENkWieMc6yNSSi
Y38MS9C1nZR38g9M0Nc5YKY96FsBczN9x4P+0qM0+fGQpED9mQD8DxlMpnuArPRCvdU7y7Jw+K65
FQAXygM2rsmZCXGRmxSYq6WBVNZV/2aYMyiO/iRQ4AoikItmHsMDh8QWoMQ+CtCeYqdydWYj85Xg
MtrCogqKwPz332wyjWUtaIOVHhHSPFBCw78YL+3LIPAGzbFtWXNXEKOap5Pls9+keF9k3KSoDPLU
EkV2clSh9JOcYaasN//+3fjs5+8JuokEeraaP2l53clkqNJC44voC/aKGLjHGN0ATqBmgGi5IznV
ISXqYtLRj5cBjR3nHYagTBFVBIYZr8xSlRAwtHifV33WOfxaWGdFlJaU8byKNahVzQembtS35k+A
PrWpjDjhFxqXBpRhWf5Ixkc/UlIybMk6aArP+IBX3gS8xjJQh54xXxyN/KHv6N+AbRMB6mkfsy6m
UrAXdR28N4ZEz7lwkWguKnaH3okTt0B9YwFxkc5n14h4gxwDpqnKY8Vvo3skd6NjF11Ex7wq1kYM
LcoYrpKePpl93y9BFjdbUCV6eQVY323QsC0m70DY78/n0CnV84k5DEqb6kS2/pP7ZDz3vmtasEWh
l/zYSasf6nbCFXu0dfbWlSTob7F+5vKia0a/hS8FNCr9h1mEkk0T8utmDDvD6oju7xA2wYo6zCrh
BsBYyeLsmst4TY37VIB2zoQM49W+FFBUw5uxPxwbnbBJdifn/JGgnSaD2J4J2D30iMwyR3dzAAUj
bHcIngCzZiQMZ/fjzFYR7NTVkjo5cgn8q27p/wBoxPUuXfwHOuxbLt3MSzNJgLLhmHDbQBfGuMwB
uwv83a74Nt9L+mgYxW3B8zKsfcKqHM7d8pip6oetW+vvYwcx4hPTj6FX46rN4UcOiW9YP0eeCA6a
EBDNnRi5+XO0Ioh9fP3QGCjIDYywTObIcLm8kRe4TUy0TWQgXHRZtr9yQlqFaaouf527ceVzh9NN
Lsrc+irDrlJ5a3c1QB6yutfkiedZsi7i4DNjZaliY0dX9zCbSJjbEoo+0FB/xvZfBevukDrtLIJ7
gxibtadLLeBr+0alDLhz5Y/2U0Nfj1XDHbu2n1qhwS7Obh//szcKHc9FWKfXtWwoeXmN07t6uUls
Ese10jIqTy97GjfJ+NjNO54Xjlp2ECgQWvUQYl4FjjDFj2TS/5W3IcFF6WHh4xT+Mj5uDTYf9Qeh
+u4KqKf0YvTTNfvnr8/loDdBJYl4D/VYi82tBu6haCDxI93M4udMlgxA2iwoTNNVUTRsXOjHsW0k
7gJ4WhTsxDHORBz6j7Rbj2PrMUyTsIb7Z7hxPMwJferxyEcE+CvDlTvdFsAtDuIfpfAHxOS/dyWl
W3u3mWS+NFm1SygTl4DayBKLaZtdxOFWZCcWYfggQlwnO4LLVbo1z5BQQf9XHXgdWtP9wEVsySgq
SHXhAizMXaVTsVd0k22Wp590HGClQWBFIVzzCRR5LLnIm9pTEp2MKkJOLhNTTPL0OLHbwvPEP2+q
goZ0oF0GY8pjX51pDPvoxFq97W5aL9NN4S8cwTTIKN8/d60VrgzYxQ107OjJvX777qyTb37RiG2V
OcRJqd+HQzeUGXzy6IlP28tvnuSuVx5cvMs0Cif9RhoPxNezT+zoiMsspk6nOPjtUx13SGXOac5R
toTxA/YX+YSiqm4AzHe3ofcrDiuhkbKfdJEgzFa8cJu64lUgxmDyGtW6SDP8QAlGHw5cS9cRMYL7
S66jFEbXYikxKJBCl+O9adz1bQG81icV/rU5IjMjldlSonIZYjxrOK62x78WvTqIfILqgHc0N4lu
8V9//jARqUK+CsgOePHMWN0A8y6ytvuciUIcPYxhBU0ezq8qT0YoTmdJlREx9n02UD3lMtts4/MP
qjeB9dOy4Dy/JU9oonhOWlCdcWQAcxdozng5sjiDBWnnWVZklgnoO3E74gkDSoj6ld0Fbb2olcHy
dZtzuMfCpvmFxw9oE8qsOUM0yPCMoO52yy6GwqdPIo1le76xxWVtiK5xkdAahL5oSDg/qwrv7CwC
zzLqfcDeIv0bK15bJQVx3ELQPphnzSwaK+s6fEqi9+EOsI/GHLhe/9GUU99gKXqrZ5yLp0o5LpPe
5AqpFJdnr+UVEIwA7VSS1i+kvSa2l9hlcyhM5QjotablX77lXFd6PYVdRlzqnAAlC8dkkS5GEOXD
Alr1Kj///GIhD5fTHJbRNxiDflIKqDwJ4GCdiNV9uJxRCPh3w+WvWDd9H5sIAeAmvrWdvZxHt6Gk
rKPLUTMLAaBQOMyTsQUNbA5kSqbIbYwGP2Dz4S8yqQLTcn9thhm6aFdtbTBIibqcQ8Z5rBmn7DDu
sw/DVfPId630ye/Guv3CbjIM3rffhMY0H9F18PA6Ji0N8slEI7MHjm2mOtv7F42kxIHloIvNfFuI
N/2cZP4hnWOflMMpW7kaAfpXCK7Ge5Yc37QQ9wJr1g9/JCNTBNeIwyf8rifqKjGGWGDCT+Z1HUlC
gS6EPU/jXYy2bnJlXxxLyi1iprWNzQAUYxspq3b0CVfFi3fbJ/3gg7vCfK8RJIT6lU3stSYTd4sb
YmMWtJN/d0Tn6abYyriSwsTnr6dGP60GmwJObDJnjxKv2+uNuz5oATpKe7oVGr71BrV6mglksuZF
7ydP/yzKrgHfClkOz7ZJeiEd+CphD34XuPgnfdymTvspJHR0cNWcHNLKndqA0OTimOw55eZNXxq+
kvddfRAosCUb7tM2Hnwku5va92VOCOxoR8oFs+5rCdaSTtTj/NSmJtAL/479H6Lw52q17najFEG2
BkIQCV0qpIFI6DQtnhTOC+fQBddumw0v7wpJ3TgTEkzwI5wlYZLEyTaB6v+dZbvFxgh6fndcyvyZ
r8PnNhslvcC4OyNJx564VNJ9unB8ov9Nk2HTEUwOhla3VtrF4wJ4HxLSfyo54cFVvR25FMX/mXOP
mG2pXUmvvuPpPxeqDnaka5fNGRZaHV7045aKko9V3Rpav0nQypPNVQf+bn3Ti0CFQdn3eZ2UOeFY
R8DFaDN1vvrqc/B5EPDI39FpanraHNai8GnoDRkAhQI1WYaLA9pnZuiYS5YnfddVo2K+kmS9rYdM
K8401HzPdDp6sxD8X8VJv6yZdi1GJmrncVJHDmKvp3rkcSf195DvWBRPdn/czUXk8gEVyffwKowD
zKhAufUgerh8id3t/eOj3BwB+4bKFa823Lk7Apb9TOrY0c3WzJt5RByMmXVvpNnfW68+gQba077m
dcYpfqxdPam6EPPIlJS4zPwi9pAPZzoz0FPTj3v7wHdVPMYt5bTRfvHAbn9Ui57A+sKv6fRK+7IM
g6qccBegBSCD4WXFud0AfaZVTeNMzCQnjfaRrqaI+37eKOQmpBmMTuhNCPuBdTPU0WW/Kk0Iu/U6
LtptlJLT9+GWUIM5f1QWHF4N8PQOxJZ1Bvsn0qDnTE44EXF8YWKcC2gALjL5/aN9E2DcBNNew3FO
47t7Yvy7LmwQKFYJawkmuDAGgrsowqEX1cP+cHMzFIWZ7e1l8ADyqCjVKP0d+5R0IkRU/v1UrOmQ
JERurGqSf1/KoM9dns1WOLC8ZRlFnq/4xy01/RU+jxhRwJltUCtpyA9Nr7L1BIlLnvtV2INSESoh
GSdlMWH2hl80yIFMrXvIs20YES+qS3drnrpyDZZAW/T+okIvoOLmSsD8ZhFcwu5zGVTOFXYkrhO3
zyljYBBeyceQK9ZnE6qvlvsgdVZmkX76cQ+r/S4C/zuBnj11Xeeu0VMJBBWa6gIwMkPhHxCh+lsW
q109sarTwvErZXRf7xt7zKuGo+0glV8yVe7cn6LfcQHQhLtU/mV/9/zQKQY1Cs3V5n46rf0u9o3C
4HN4bLi1CQ8Y/UgWZknUu0x+m8N60uxkzM1HWhyxY5MQ9t1c8h7B4DpVqOpyxWe86z0hsXN+lbzx
8HzuPSM+t29PuDJt/8pah+LVCaR25TxowGAS18gb1YmjPaCkN0hvNZq7MIf0xVyF4Ep/mam5qRw4
w+gMKV2I6R3dYQFtFFg3oDm5exze2JkqjFHzezoeUixed+gbe2nqH4h9aJXR4ZnpoRu5ePIue+P7
As9073LDXhvFRC2DjivV7/Pe/6Eu7KAlBho2TAob5ag+efkpd9Iq4NWz7qhEzf3pTGAcfuI8K9kn
T0kq0tuaryE6Mnp+qd09EuR/eoYCtgLg0xAzs4zNeRMiQcXxOKKAULAShJsl3UDIKtTmSxT73dFu
5uIXF31lFngs7Cuds/ua8rvr7Amy/3kNg2WtWqCM87A/Sum/pg/awmO58uVzVoauuyujrUKM1Eei
ZlS8NTIuMPu0vizDtfFaxjBGiM4R1E75+zUZMZ0x5J6ziMNhe9dU78c5E5CjTaAINnGNVBZOHhz+
h2jNwGQdj1cjoBd1bnVWadeoyLFPfzm3catvsLWFfQY1CLKfaXHSiI4qUyF6mvmVUnwF/ijigCNq
PX/vFOKGJmIVMswMmLsFfS2mfthuMlrucIRMA70RPewxOqrTybYnmGhjhVBLmPOsmsOrmfmGp80X
j7DzMnkFMDHtx5EtpXL6zr2pFGbR2Fettsh+50KYPJ/gGrlNCNuwNJX8nOEmau7jrLQY+VW93fLd
4mJhu019ZB9eUWUWbcNgIUsk7iZmElgBk/pYLQAGL598ebOQj8b8QsUEl3+5pTnrYyYLIY1krGdR
qRqxP3UbXK8QxORRH9NCtGofES7KaSR96JOVYkuM7uGLN5N9KWjscjkrt+sxZyDVF3OJzmXOphTf
jMW0JBLUm317Cj3/JIB8zx3cYpm+Zrxx5xtQc9wbEVbSzhzpQzOgmAnbjsTWthqpGjRXrqT9T18V
9kL6cML23h3e2EPtdNaNxTX14Y3xM7KEcQQHAKNoxqaLuX/lHZKuzy5C0RGOKRU0QO9V6yL/c1SD
AQzoMgAW0FJ4nLPaKoeOzPQIvnqGj5SQD9G6o9REljWUVz3SpET7bVROJMeVmeieObqgRIo8vylQ
AK1O6XqbyI+A6JpLf3mm3Fq173r+L04Nch6y5dn2TCd18QCATS8OTLMNaju6o/5DpSYHMf8R6ffk
SPyl4vm0LzgfEIUHdLK7xxOfgclBO8qiNJA1KBf+8NeaFecQ00rjvCUNq26M9YJT2PEV7LnIwO2w
00LRBlFqS6DRZtz68KLUk1kE4rmCf/wbj3IQq/jVLrmlV9NzP5+jNvwE1fhfmkGODIaI/+ZVhU4G
bB0NEa3ohPmdB0xS1PWpUftdGGZT4CAwqPuU7O5op6SxHoIisiq6DJO8bGPxzuJIxMSWPc8ylpN1
CDs7wdub1bS2oBR18n0dEj2rmKSHWkP81x9/9hrigLiX7pQK8IIPjfkQCZzcvwaN/zQyBdTHUqEn
vCe96oXxf58wGa7oQuIVNUk7AxunjfZh3GVRAxq8wBXfJc1L1L1YLFKZ7jSGCD1DT4vfs19UlAob
xzfLzmQggMN036j1iOzSIwarOSiHKMBQhcYJ88dhGcJIc8CZ1BU5WQhoQ3ckxGNTeuw5OBCV1ymF
33biKuTZhg2Lcjc9VT7E1QQqELBBhnLwDAvqx1xynU071exMD0yBpy9PvSqb7H1vpRPd286ptoh4
Rj4+0zAJkzlYz+8+YD2XVn8gpiIFxAPCxXWqyA/pJaFikfJ/athUOryIidluR7Lk3HjNk3Gk83ir
zhkMeqmlZnexUmk6BBgGPsaw2NYXsYwjoyqEl8D7yLjbpe5ervGW70zpB7YgiyD69fw41xpBYWMR
XoWVxw1pCDDI1+oillB22ODlqZbEmiXqKceRoHBVoEVXE4pJzg3AvCfLcRwHPnpAte9wiSHV5bgs
QwFQddTPobxUdTdak2aLtNgqvWDC5gS3LuS13G0f9VqDZ5QrJTtU0bcNtTS7V5QlG7KABZn41bLY
egKv5t2U/1MAQEIjGW6jb69edx3Bw6PKRp8RBSWXDViabz3gCBTr9Yr9MB0EMC7ARc9Mxe1qOYTE
mJWSasiANFgoGJsrNv/IAJxsC7uz3S+NFtWnZl6gmCHApXUoktOzWRuD2F8tBLLbdqFra3gfQGO3
TwUBnhgqpjisUEOtSMHyPaqKk7FYuM8B756Hcx7OWKlhPkmPa9lV67XVsvS3RHY9TkPWYXUoRioR
c92BN6vFkBHNqyqwZ3r21u2r67tGSFkZttXH9qCKrXRI9sbk7bDMSjle+/P/iVAp7ylO570CZXQK
ruZs5VI/rZ3i92BxVmNJLlCTI2q98LrUDJwPfEv9JFuK2ymQtap05ASmOHC2A0xxlSQlPx1FNVwm
BeCEucv19VtdoiyUIjXt0ynKw0QpDzNykSyBmeqftbwtoACfxDn+8S5V8H/obwVzxcgaHNylo/qJ
LTIspsfbRnS8rlYwrB5aSgxEL2wdPr59mo/1czRS5WXHzu0tjA4Xku4gmcOgJFyiUGygWGNd5gBh
Jo0j6nJw6dZrbeDB6Z2dm7CVIUbQitME4ATWH8+WKpfXFcaJ0+k4GbS6kU2S9dJM7odNMElgkWSI
jP6efWcT/yP/UMlR/Qr5QcmaHy99UgnTXA0aXnogsjz1kUXSaMMhaS1GBjG4TvsUhzin2UgvSMXA
5Qhm30hx8nZWoWgsadJ7A+Z47fUo6rdMsWpD3KvTEH1VEuDYADcVTpPuvH9Jdt7HKA/OloI1uQxt
324F3S1fzrpPLvxmNpjkxU0KxhFRGGEn8Y3yYGoVJ/gk8cM6TFx1mb8N4FgeJGkT+wuBDBnh2FES
x0y7vOKu8HIvMUR0wDh2HKafqniNcdsCDpz03BQ92jYrXxtKtecClffeB4oBnMD6swwRVdL8PNga
g1y3FugIrZHL6D14tyPvI3OwXhHySuQ9L3ZcPkHPnIftHaEOEv0zpsnz319KxFVvgI5eRt2agq4k
oMbzW/K83JsFfhmalcaxmJrwN+ex1w0XMj79IDPZxAU7/P0Uvuj4KSAEsQFXguzbsyCkHvoXCOtu
0Wvj6jH4NQk5Rh8CcGgCxlCmvas1+coUzDzYRJ4Md5lzukx7+cX40tq3vj6b9kHYMdZGLn33sCQD
IHAWHhoeH7SytnHFYDBYE1cUTXk3b35uAz6mzn43DsDAE8YmrYd+Jp4Rm4NDnjQ5LrjnM8AeMwPP
eUa7U2lSaN20fpyMI1GbcFAJeS6lnLloTTzKJRfNH1HsOcC6GdFBd536A8Jx7pql0nD1KPQYA78j
xjSHJliXVNTBiZJB74ZLuj7m3WamZNVF5n/N1op97nh9MwR79Mk1uBqA2F/r9XHIxsbvQh3iwR0H
paoQHvWewgJsZn+H5qvV5IhDSJZ0wBAwZRBJaTalA+dC8XAwAWfME2GIH0er0H5J/KNJ5nbIQPLW
5wpLEC2aL7Mt8oII/9Rpxn0M39WrQw80VmlfF8Kcjn6V2NxKyOKBHelI99Kaujs0tAMlPr7J0YLp
Dc4WFaak3IPg+/6udNuJjnAZHX9OkPF2girkvS8OV3Dh+JJxhE4gIfbhi3MsksRjCBynNTZxCnv1
3cYDh5NVwc456MD5mIXvSshsAF0TrAQZxZAhZxQajWmMx4NXUn3Nliw+GGYUW9ZNhWg7SOJ8757u
sBGvFT8dGEz6Ff/0ZTy72MUF58iqRlP2vQCQHfG0z29mE5+Ho+TNgrQhbjbE3p6vP17nEcxw5KmC
XWtcRYDOyaNrOgxLn7BPNEP+6vtHJod2EVES0j+bgiCXpmHZlhXtu+ZE+kVrLQ24LaIu+e+bYr2Z
c21jrb3xFSiY9nVsfOJnyLbkCyhfroWo82XK5xzQL0aG9GS9HZerrsCspznbxBcW7aV1c89ZB9N0
1Fwn7hTfSTJByIhGSN5CG4maGZBropsW3pT9Jt2EKQuxHu7FIXustDao6J5CwzAGKEoHPR00IEho
ZZUgPqLiCEEIhcuJLwLKgFKAGXeT20gLvy4rnJYbLK4jfYQ81iw09M4S85pI/FwSeTV1xgDLrLRX
U6UvTuKG/YTb6RMEMxOKb+Y88tj5CWVXO2mSyfUIAXvcWSJ+sdDxh6xjiSYM05klescZYfPOh7Ih
qP8U+OQfDSRgQengFRUHQ5ztim+4pHeDequd0TnnI0gRnMyghMY/fUZJU6obkCkasBCq/b+7u+s7
/ZrCwxM7O1nOcGVl1aTrILTnSLNjgNwDGuUHCLppvZIFvvWOs78n4277ZrTe/bn/4YaFundIVCRD
PM4N5wjAqmggK7y9cdfFLHUaSK5VXr8Aq4vGwMuhKxaXQTU9dyaOtAb6Ebim28AAQaiWTXhe48FK
nqVYXhrzSr9zy9XFn7bsBjy2YoYxfqcymt//1wf2n8GLRMnWHnJNFO31Ghwk0SXZ1+HEL9ziL5C/
/tDj1Sq+wtCuoEhpaUIWOd1uDJ72j0LaebfPRA/PIwij1cMMnNcF3op7t4nXp6Bwxll6yYrEoj1C
dbi3s/VL+hyjBWTi20vVliPVef9+uInFM6Slh//pTgGKJQ/espxH/yNBzeacG/ibPXW378jHxLJm
0YvmcnfEY8+jjC3qW95nNJFKU4LAEJTzgCKIkLKA+xrtaipW7bKENDiuCphrlOWZmEKfJ04KBgsC
sSL/bKmLnw+c+cPA1psmZtcRQE1TKCxl7CJvRvoXzvyWt2UwP3B7bCT9gjt9K5R2E4lw6te1DVI9
9QcuR783XitQLg9r/IcCCFbCSjqT1ofzA9pgo4O+UDEgHnN0znBYy+98Qeas+VdSqo4PPApxYWou
waaNe8tCVOxEgL8Vq8UKwvKr2VgvFJhM7n+lyHs62kCPSHHEIE+sclds6wVc9gF/3yJw8gfyu25P
FayfotbRr5AbVMo7razkaK7cReThElCDG4rLtaqX7QNv847MLJ90bfbyGbG0doZ9rMuHq/f3u1wA
V3df0P9lT3s9rq3Mnt1u7CM9p6wTdLwQ4EsHvVV0gXaLeGBztnBgxYnPmmMeqig70n2T4AO/gL1J
My+YZ7osYtp/PMU9KcKZ6IfGM1PqXapEHt05NOVUjXBEhfEWU7DVbrVP1Xeir+jKXbcg+bakP5kd
aHgS7ai71rhq7ZAiboKvFyvQwllrnGxBR7HZ08mdk4Y5Jy0jAnrkEEknAIDdG6VF23yU3Pzs0Sk8
z6WXJr0LrtZqj2ClXSozmHXSswCRwbvZxD8z20CpAdL38W/NBfkplcYh99EixOJ7kP3A8i7uRQLK
wWCzz6BXVMItobBBSbJq9FMFbVvaOIdBW8weOcgAGoSO14VtpX8TDqWzer3GS2x7KGKGAcbAaKjG
sZ9tLSvbXy0NLJxtws8wT8TieuV0WZJcUBbV9VUKiU17CJAjWMbt4JOv2bv/qzenf95QPRm6Rfvz
oqOeD2U9MTXoeVrbiaUjc7S/47mGGxTz/GmZipqg/gD4z7e+Zhsj+FF4a1iuEJfKDFqPzp4hx59J
vMS/w2xogi1dkcokkX/MiDSd3u4qP7QhjSHlXO+wFbZf3OpeOG6a8RlTFuJHDIn/9gMFIBlxktKM
nlnbN4SJgIdO4SmRD04JRxVsZQeWB+EkcSedxJb0jHxmju1+jWjJ28D0pafxJflBOI5ig/GLY3AW
Z5Bq1SZlWYuLsoN8jY+9EmH2nEhwf18T2olcPIV0XHYRll3COnbwuNBW8A/3oLb5DlA/Zryzvu0H
PRzoNKN9f2Lt9iLzvgbNc1aW5E2NOKELglcuZq0KhYe0GUI5BnXNfbbN2NSYf+XRJy8bii7qJmtB
ZjfaB9/G4UMC69hmPW0mOU+EQgpONtYmO8Ugc5r1DXgCm+96LnagDf0erR3IEjYlJJ49Gx8zO896
rtsQLpeDg2YLoPWOaD2Cg/z6HWmAyITeeFjAryWb8LOIEiNAAN1+tQ0ib5ufPLihJVJyNX7I9xcV
DOHi5uekFOtYuvnKjCHW6roJ5nX4O+jdDtvy9+MvWQh+BBIH2oJSv9WgByyowxnyq6Her+syRdWs
0KoVjgQ0+xO1iR09QUoZt1CkHC3SyqsXRXf0uhZDakDX7Caj3DOHMcg3veGYgm4tY8nICp8TPkvo
gzsqlDcBdkfMsRkWH3RRWegppCYbjtAvXRMFVB5pmMb9b0wQIJ/Iu8zbnyko88Rv+igCmJCi2ZKv
1Z2g1x0rGYi2sQTPsbH4JTX7zD1NssVxZCGIHrLFOL1llTwbcu7SXMmACD5FYnYwjhf48OUN1nRv
Io8oaqN9yeCZeY0dMmJyeqjreNvhGINwu8P9dnHsXnO8h9wolYP4Ixrb8xFSztHdG1yMTM80RDLO
/mG454Hl4hv4v6d0PvjMarK5HUFr8dXQ6SKGq8F44RkS2XLzKhBK/1Nx0NLlglqoXr4sk9nbveiT
tP6hzmFK9sMqt5znffn2CgmI/Dlu8w9O3xGmPlKRYXggLAN9NTpnQZP2FTERpiq32djnXPCaPtvw
sdCyrLLk9rmL5O+OnbAebC6TA+veQwzfwE8TSLDIS7Q4LBX3UNZll63vYAohb8zq4SLs/weEg+yD
FvW6Rjzlt4OGw3S97J/+0qVXPQ+1LnZfBxsGGAzG1HXLct4ETrSgv6wUBeh+CXELxN5cIdTbKmyN
7pQvo9IAzSi5UD2Djc8aPNVPVGZk/K8TaGGpzYEPf1ArlH4aPsFtMxBUvJrsmTD8um51ysi5Dw+t
nDLZGduJsOtBVVBwR+6F57YX9URPqW9j/ZgEI++s6+0GkT7iYW9AupzgsIfkVpYtl8tHjBaUFnCQ
RpYCMpVqowhQDDlCnvOdJPF7h9TCs66xrNpHdqaT9DRooB38zwRh7FuYQUkcNBZcooqyQxhnVOxP
MrhJqE28XbnyrvaGdAWtfjx0qePrKrXJeJhPkSr6OGEohK41wgLXm3WXVOKWil3rfXTXhDeNVzHK
bhDY8oN/ZMlEtv9RbqgH3ynBKe+x+pTSDQnY0dYi93yxF+HpbkN/FCMJglfOvU8VOTrhQv/xswRF
/kD+RovoB+0I9zp8iw6iuNknvgjp4ofHb00QY6Mh7H74j8Stnd3JcUZ6n+aK+WHRwP1erdPsIcL4
oQnn2uiVrNfFSh9aUzyBvyZ/UMlksinx8ZEf1aVM9c9+eJErb9n32EpVD7aIZ9CxT4Dfk2LShFLp
c3lQbfzqnYCKfQL0/pRM2Qf/jvgai7OGyNdBJb+hJeGMnPiP7mbnb4ozTsaQr/H2SSZAKb/UaiIW
k87YlVtA+8rXx5HZpiO2q39vjIm07J5ai5fBsNHLuGM9CyYpvxDCZzSmBu4HgHUI8b0HHdyRyG2W
MRPIddNccvVMO8AnTOqYzv/ReCJScj9PkZeoBh3h7lF/AwdcWk/+aw4+/GPNsekkWcNJYmKM48hL
LGdna76MbHcJM+qSyAIGG1Qi3VZ9MxEstTmMzo3/UJU5ei8DC+4Ei1L4/zXd48eX2dl0lBZXOcpN
XldC50UnifAewoVZ13nCLRyHtmvvz88BHhGXllUaNbsih1/BBQknAyTQh2F5QWXPOlNR5mC7TJfz
nyku6A9WxVVwFjnxGcyFTni7IHY5VEgEKSeA3fO3wTIkXgrP7vmsOcpei6I6KmHkSpFW8XP0mcLa
gSZv5FGD0Vnj6YnX1iCO8qRuPHRlzy/+SPWjI+7yMHp4cVXWl81WqvYygI+qy8whfqmpcFuipXRI
RLdpxjOGLkhO74tA/WFHGlIOc4kP8HCloctfRLuHD9iMx9sIlQJEZ9epg3b5oz99qjNMpLRSxhgw
Fbbe8Boe+qfuipomS/+qMinpKqh8yxY3f+uNRAtTR4WoLnba8AgW36NggEsmJSZfDyWcEZGrcHci
5hSvFpSlvrBW+WnyQ/460hCwcMl8HpE7cv23Rx47pKXQ77ZBiCjjYphevBUk9ymtuiQo24JTHhrf
nVCRfRJ/DsBOtExuYVGIOtYFxVlRTeGLu4pNcB1v3Ycd0ihXJWKTRS5WNruVZJhjjKLrfKNatv1U
vyH3xAZtnR8xDliF3iAWceqyC5yh5qopuqQcOZoNZgu9WmS0iXV1VA4TOuCZpt1XSffyDeRCn72h
KrxREacyDnVtlJfj+jCa7RJfA+/ZUE41az9LQxauWmRjS8eHDqCpFHgp9nWC+IbdLvCv5vVxn29s
4BLeHmFyMOUZuWjYPdeOO8OtEuC1Q5skSphEBlfwgOyeyYkGgWTQCy6N3Z76GA6Opo9PVst8Mdwi
+KN9xgFGP/+Oq7FUUSyLruWmlQEZ7cFQ7jetZKogaEoHbxA59erVv6BhmLJwbNSs5ZEBgOUChHQS
WaDAZwz/J43uxCrQoaRTIfxWprC0wJpkc7c2fmnej0ubvLrIILW228sMuOC2Ur9VplzG1f2ERpAl
Y2xutOkZzSf2zWX8Q01nR+081tVwjsY1NqN+kOSxDpuG2N/J2sCgEhnGfISpQvN+rPP06+GFFyum
m/qwqNYiyrEqEtv8SnwGiZRhut/xqBCr11sTIKwcGvcLJ7a0+3xtQeyJ5EB6Amjc4OYEnckEF4an
wVv9gj3L8rfA1RrZABORiX525wNcBRfYBw7TDDqMU2fm/yvtA9rNZQGJSYj7/t7ZN3K3FSjTTOp7
3eGNA7xoTD7NPK+9h9WoME6Iw3Yt5+v1M//Y4k7L8lVUnKvlvy1QFAFcf9D4SlWuSRoum3SO1YCC
1M0HwYij4IEo9grp6BEDLPFMQOWaym33Or0UUAslSyAcZK4jzxy0oKBv5mLtTa9XVQbPZQEf0vxc
Cc/pNYIHT4COi4wTvyTgU8qhcOkBMgP+Dpl68DSl/JOq20R8UcV9BMfvYknXiuCS5JM9SpOkHzu0
YOe7QbXSGSHM4o3+IF5OOe2EL0effhZsIqtLlFpbxeGg4feYVTFZaILDRIbGgUywj7XfAgGNTd5z
DczGBQZTix/rTI0P/oC6WiY8NOXk/ngEk3uAEy5t2vKVFJWGSBZmBM0gmzhj7x1zLrrvMyTvPaew
3gLiWoJKcN0Mir8ymE3phRt4NfE+9g5KF9I2gBrka438SZ2rzxKpImAzDApYexsEc56FyKAShd2Z
FnrKYR6f+Tvh7qiGSERBKB0VyHaCkVO+OEC6yvMXHps5YirSKZuWLD4lVz7bFXQGlIZbbKFXyqIx
e4BxKccZEsULbSwkLFFwp0jSHmq6AfOi1tQHMJCPjCVRAF0k0lfR3vnhW5wW9mA2unEgACrahPy1
x+PcnusynKxZXzZaT3too8t1dxxrX27iDRypfE8J67r7bZguxJGxlweKbGt6PtxHav5heL2UIz6Z
XY+rOfy0QTuAgjmI+TqSzvcqTOt7Ko/XGE+LoGnKBD6kIMcE3IdcZZPbKQlqQQn3juX3eu7YPjAe
fMGwi5RQqxKyMH+cvLOrUAU+5CsIPtIMPkdcTWdiRu+ayo3NsDStcsVNtyJ4H1HiaqX1rgwsBfgQ
Vr5epA8d1J15su5RORvgSfCZK6s2fhy3h3EKM6LJbKvKFLgsTnALa7Fsr03xz1EBteZTAnj97ESQ
qt4LlwACSLM7g2II9aosxDNMn0rp6xVCBdMaFSVpGnPizCkcNyZMFDo8zJdXLoDel+YJfP07WiUh
z6qtdJ2kLWtXm8+CgExAf9lXAegm5sTpd9JTYENcboV6t14SIH71HELpULTKYujIzr/2ulfrp3ao
DNogwIRCKcBJURjOIOZoou9XsxeDDZs8fGhKLxs29ngeRwhTAgM1E4wSxRON5OQ4mZ69LRIiNA2j
dJsKnubMns8BGOBxEVelJGFOumu2gjmoOO+yK73wTmRhg6+tmtQq3WI3ckkfynvbX9LcZkxQOxfl
/f03ACxtuQUT9ub6J73ciO3fYZFl1S7W8VEY5XeHNsbCtzzdLifxp8x3bSnMPGSEMFerUVL9I2VD
UFqFvnH6D8cLCpwnmv4NTfZDx9RqMeZQu3FkQtG6ekJ/OVj3ovKKu2P5uP7cIfJKXx4Jon/tjdGz
9yUEY8NXPZsz4Qa+SpuC6ddwiU/YUJcHL0JU/KnAOFAVo1CFzcegytFVbaHqe0h2ng4alLKh1sop
nygdBdpE0YwN32A+kXECFqCoBfpGymVnKYA1XjVAHn0YeRu2FXUjDeNfwIWq3AUx5lzaOmtapVpQ
vLAWQ21a1t6sxGyiB1HWiHuLFrOSElLHPvarbb1r3EkUIQrXOEnRRJKi9giX4uIBZbRjBtwgrn4R
C0zRyeMFEIXwpdDDG5OYp5KQrSMaISHfCJ+FdYGYuACaMloE05nDzYAY+YcDkBCtwSuMlqS6EyLg
STd7qR7ritx/8W1uJULX9ILVuIm1YeigRCbzGNB194COxCLg5NMTXDgXxFjdVCQ5E0JCjwOOJlup
gq9/v5u0/eJuS9SExL9b2peIREZw5ocGti9W/xMbfJG/yb2e+jYJUNV9fu19O6HMVibm5QxCPzxk
GMUMWysb4F+SNNQwkv6823K5gmyJCGr5d0/fgk2BLMBjoF/J1nEVt6B5hd6Kq+O2qd41632NsSpZ
6/9zXt9xaxfvwocEYARvsmgqwIpDQ1RXKZpXJmep7Q8q8LyIJsAXrA3ktlqofHLsi1Kwu9MFKKqn
hZF5U8HO1CP2XPliANJdeDGPn1mCoursSwju1zfmoHO2kEOsVN3plFUyduFcCFeMk/ubnUg2+ofT
zh8YFOgXT7ZfB1mimUB8iPjJGGy1t8ZJAR7C5wpqjkuwraoL8FDaVUs6FGvCoVSvbPD+V/kDvodd
3mb9QkAlFfTHy26B1SKW0HGU0JAwZw/1yytGAqWSfkHTRV4xvCh0eke/kSzsoC0iLwKCh9o663sN
5Y5l8FzO4NPBZztS2iF1czF+sIfV4Vxjv8DrUgL+UK76fg28OwMP9y8b6N70vOF9TZRAj1LUPG5s
YPQvJWsFxA5R3zqMUv5XzD6CN3VLO1MD2SqcIkYVIYoOpnkroPiXwXcE8IiZKQqYrc04aLk5oKKV
wYPVDiXKYGIP+2HHF9WbDljmUct3MOzV81OOppCJw4zbh9qUPezlJla509Rfqy2UWGRwuWQp4kak
Tzmi8F4Ji17giRGi6P3QGQ2cTmuMupjtfX2tdvk/LfCzv3CyxjpnC4pB9UbcpJHjmVSo39hkeFFB
ywJ5s3Lcs08GvfjiOji9GoriioOE/SJHQiCudZSt6mG6eTKjlOlwxRkiL2ImTyVqRfYToaNOQ0vP
EZQN8EFsPwAI1b3wxsu4nh9tVhZg2Q1hLbJXGfdRiT+kKy61G1ilbAOlMfP8o9LyeeH0tJ57kfVb
tUafrFDu4uhVaxhSRimHfVV4XjC1DEPjVcG8htZpjiVy/iWq4GVozTCGrr84OVpQ26WV+uvxYpCZ
DzuaGg547Tpr5CIIXTq2p5T6c4285rf5+08m2hxMPxH4GaZ0PkDHXoR8hS4z6b3Thmh+EXyFWylV
wK+w9T9Tug309ShPJDccK2Ee8jwDty5QIl5xRP41ovlsr0cx6lJ8pnCI3bAtU+RcyKD6DWgal2Tz
7vta7Y89DyAxlRIexh4uTQzntApWpMBy12KuBdQGe6P6kgrI/7yTEEZLV75UJREy5O0CntIKpdj1
9wHwAwl4dcdR/JWVmjJ2HuAj0klwyMM9F389jssmE2C3OkGkw+66/2tl2NCcw733WxNfZcN6Ezt5
JB0ShC6EdbZRllvoodNhKv2sDjGYs5Bw476m9hu9hY/52l4ReXNguGPtlDKq3xhsNgP+w1JQ+2v6
KVJk35KvBj1DR+vL8HE6YQ5prxrP1aadf3HsS/3NIF+WhTor3Esen7omONIaRj2Wn2KwzBSFseyA
PNqn/WQfs4AFu0kALcGBCOObp822Z6yqtrzvQ2RQ1JRxNhuSOJgdI1yA470oT+fDFLK9+aqzr5LR
IjOnbURBMcBmH/bTpDEZjjNdP57PTyp1Qsg+kTe76qND0V6hlNP9fUC82HAPNuW+szJJTiLiFtCU
m/+PVfUEIwkpvzUruoNS1v5LzXpLuk4TUMwfqWqqGh81WMz2MwVVA1SC5HKAHY8PAOPU4NDmfnIn
4OBSgin1wGrahzJe32pody0p3p4+rnWw/hdHUV4Q+BZ8DOBk2LNSqeiYVD/tveaMpNBKfWZ1rlAL
s2Rf+j/l79XWb1w9ipzWP7Q8spr5cqqtGW1Q65btoGJgZ/Vp57sFGyMXl9gs5z5UgGcT4pWB9/Oh
QDwo4OFav9W47QCxTgnq4zoc4iv0I76VVUhhUb8gxDQwN9WZZ1fTwCn0kJb6/FYlN26X6Yousglv
DGUKcIFvbhYdKYtE/istDiBMMTxiyDYcg71m+v0WvyX2vrLOHl8mhNaKchEFw9/mexxE6NPCBlO/
Btj1SxAXZquFrvJ8A7EPxuFvc78QjWnth+Cjt7oPtZ3dExe9IkyrhUD3Yc9gqBHXsjl44ncf12+v
bU9zLrJw+GgzxukgG3NC0xJXWoJ0LVmJ55ZXxMhD9YFhXyCoDZG++7cdY4RS+0i4YTPXuCChPNC+
5sPFE7MpVf9z0oEW6IUUDhCNuTfTwBhwnJo1mK/XglHb7E4sIbQ0lBIN8JvewFvutnouqrfq00QU
SFm9bnGcJ5zInLJjTQgdEdne4YmCM+oNLeeCBwF+kKIWqJkXXQ5OzUxBlcBEIvAJpJdlkFSsE1Lv
EV8tu62YPBmy/elEFr+C9h42pzXpzfXFnKsbm8AmMI/nNYaf3cbsNXvQEqxw0t+9Pgr8pt9sqa7z
JmPdMCXmAL+ULmPaBJy4Ohkim5WQhELdDDxMSvMFspldmbIlY4u7M7au9zMRxNfYrC8Oy7V13Yqi
8FIgswzQlKtuZWlHPkd7VKNLqAH/ZBU2qMqYjcJpTLNosIW5FZQCsbm/C9lG7aI4BPVxIv2Vqpxs
P14Xmd3fE/Oz2QWl0wEvq369uDSGK82Pq+8TvMRmuIoYG6edJzv6Js6C/Ur5EVow05+tJv8l3uoY
apO5g23Ze4ES8c0Gn7B6mieIwqOhQcf/9I0DLd5oTVmtFiWCxaAO61JL2dE3l1vxP2lUjPYVW2JM
0UF28BYWK3YQMrYrY12SMx3nzoLdmkR/Iejswt7QKvew+OQ8bV7HmjZJyvIrzE1pxinUgnFcizHj
OAyFZvHF1TujNpc13FeR0p+j+uueSFiYJTgy50sd7gtEy9c7mmZhKIJXuNkWS9728Jl4xqOtetE0
OfWfEgvvVBRb3ukCFgUpEIpA67ppyNPyueoQ9kv8KYYIHu2SODS4NfCGWqoekHUTjZcf6oL/d/KK
js0s9oOOMsppAAWWDq7iQxCoJEN9q3ZftK5NwZT4SEsbqwfXcSjZP4MRtCcdIupfH+doJrfLxiE1
1adZmjJAVWMP1lh3CStCbLLjDBB9tYR2fWq+Xi4z1fnrTtAiWLUHIdibAL383dogQc2OJ64QDWVh
MbcfZUhvxw8Wzd2qq48z70SxXtkeebhIBldw9f10gOQS/BD15X0qkFqYO+F5N6XkVLUIGukJce4n
15fwM5sEPucvUDQCd/UF0zuD6H0eTYkvcsblRA0q/3MVbvZ+oBKHXDINYzS5fcmChMoz/LjNCfny
a9ZLV28BTSbkDCJQRZ2Pne374jvUAdzzZxP1mQSUhb49ird3QJ6cMUPyL1i2e2JEgmq4oXjFd8H4
jrR641mljCqhbfdJhuvskzGPVTvNaeWyG7SFDGYXGLCX6RZ2X0LrKeP7EdWskZ4stjMhYyCNr+p7
VZodmdz1orA3XoEiMrMes7bd8/kWJbFjBIDxV8hlpRcKKV3JPpgxD6u5nXDOLDh7gQpgZqhV/YKF
OONnn53OtG0kAHTbjaB0K+JEBo4sy+0L/1+/mtZgXeleJbVea8sQwQeDsR3X8wIbnG1BFHjKgtTF
0R2MmVVfTgWGNHyPp0l0yMyU9MGQ4vPby+IRJwkHoPjoEqg93O1GmljoAGIm+1g08GiJO3lBBN/u
cqppPzbA4xQ4SpeZoDC4mznJutFbVfmA3/atOTc0t24JzwFAmubcT1744HxsX3oCwQUBdl1v2KuG
ZRJ/CHDou82+Go7lI4egQPOYyuVrobptNQXKa93pq54NhnYttZlpOyGNFf+Gss/ZXF816pW30kt1
VsoVE9+rvHWhRMh5aj3Edy0U8W+aBCFDOifICSPmDilrFHC7tYZEQQ2Z2mKC6juIXjeMDPMahWls
sxPJsrsGueBz8le+8t/yagxL0f0kTfRszLuDeXWVlXkvYpKJT/vldPg8RYAurMEapiOKdk5mc8dY
5aFfDNeDv2XVwPv1Gyc1e/GLfH7ixzzrhKWP4QgEEHjItJDSjSvWQcnCqPAdo9V0JL7Boobwx3+/
VN4x4OEfqAob5ex2HTrD+W5opXJRI02bi17BwzTxNAYNPAiO/mk6zhE+hSU9LM9vteW5AS/WXIVN
aOEDsDNcg517pwCXRmbZXHYwSmZhYWUEus3df4hOKoIWg8C1mjtRTPAyHMttD18UqxtQdBggmLiH
4cGZnbB52e/tXlwz0dhGE7t+r2jzVG/28fhu0NBDfEB2XSuAkPdbDiqlijKCbk1q++4XyPCrCtFq
b8EBUa4YFYMURW9RrcSyNBqzIWy6zCK+/14Nd6bqaeaCogW3Wg+sUizkK4RLW2JO4EA+MBzt5ijI
166bpEF43Ra/z4XqFwRIrgx/rp0BB8tXQBvZPLxgFM1IW6ewx/Pc14NvrIJ5BRVzlywTK+bI9x+j
GkRqKpvobmdKrnde3leQe7rdlxQfn+nLhslY1XOtTC5v2LPHVMn24zbtd02K3OEC9ck/vCBplTuU
p98GKRKeShhaQ/5cA9EVfU45nBVXyt3iB/j1tW+wCWnpQAIWrFtQB2lXZ8PRL3T87N4NE8m+T4OC
Es5DG7cCLYKyIxzHssoPCbNf9/Lz2B8HxvoDAgOZYaokdWmRQA7uZWCr8CmG6AIKI8TuMmABDqcr
xy3qiVUDJ6zxWs0LxvF+a/N6RkxnDx/mfo1rmju4Mb8zkwlRmb5zhmnUE/Jzp5yAVv94M1y64ky/
ySlGSUsd5HzwNrv+A5jx3Qskwp+xLgxKPxgBu5jeqUoumfpyfHDw98KsTjvvgYc2FUG4iTfRE64Y
wUHhx/J7h2rRJzRcscnzu+W21Adnr89BpsGI6fMrgA7c6d/7BC8GeWHct6PO7Lj3gWf3PhdP+MeX
BXrChxmsgVifVet+mnI3iHE1YF97B3oBgrXN8R5W+7dOUFp/Zule8Q3aSsgzcEavMj9FNbh3FksD
xeVJJ4y8eR2AXyKXTLHQ16oD5XGHVef9X4DsgO7dSsFBkFFv4FY1gMXTBudSSiWaZS23Rj/YPkQi
Q+n4/CYWzoTci2Ag97g/HonxSxmUcMgYDwcu3AHpkXB68pz8xHAczSx8TX0QvD0FfuYrhW8+X53v
o8JWMjbVAVnS01xQoosweMnrUbAPiNYHzWu90EYMNR0Q5GVU/fhhOZhUwh1Y226nPwtw9hDY+PIY
usJPcopVxayt1Mu7nzUe8aajrwThfGoDXv3Oxu1RGSVM+/4bBHQzIeJAnbrMN2T6stO0IHtCwCbh
tvX4sYex1AFHxslhvttUO8bl3fbP6KMW/KZ2mJBzlvwvL+xYP4MTi1/zvL5UC2wAsnvTBN1xdfW1
oxkdYS8bdWL9i/P0PlJ4ePTpU8sqJ6TbCkLy/8+vD6mN0I7bqdlMNO+Bt5EJn/TxDlRT3PXfqPok
sbCHZ5lksJKD8t5nmxLnv49w2X+ELrIRkqcOpwY90/t8C/vdByeNVyRzinuBdRgeXu6PjUVKvym9
Oq5bIPaQ3FHBF1XTrv8x5wEk7mcZmQwf25EEJXBMEUXbjzLhBbbnD1Xo9wD52Nn7B72HdVn8xHpn
9hwfwtywdEXoTmPZrYg+bFkuzT5oknFAVLZYaN6MMyeLnfKODgMqBYZ8Juj6s2e7kCH1uEzxO2f2
rI2zInpsqlB59riAqTm+HOJqqfA+VfUn0LDEUX1FVHHqMdTL0NoQdRA0UdFDXKHmgZZA1GnntnQk
gkDz+6nnh/xyw8dMWnyYwLLGHpRc7Dy/EDi3mUTga6N+3wgarpivHdlqB0zRn2BCoTBld6N9G8Ct
pc+04val08Y1mGVoFnx4haWd+bOnxD+kMafBoRObmqwPBGdpmhEU5rr71YGtvKyzDNCFdUxSPra0
4AxGsmmP8GjaL58PQPrUZCEI3LEwlfAUp4yhXh2HS7snFu89ILI5e3eMMak9t6Y/RW9TrGM+TFdw
ZyNL+g1LGW/udg0ejQIWvcVS/9oue+S0WyyPPYsuIHBoOfjO6BrDSx3Oj+7sa3qHSepiPeIKGU8z
lE/gi/NoQ3xM+Bgtk3+lyiDREc8HPOw8b2YuaH1yGDpgM9mjyXN2RBId9wZh+jurcf8mmJeIN8H8
Gu70bvfT8yd3bBHZXDRe/Uy8WYR8Vi39BY5eXGpNFsq4UUvX7sWBc5AVbuYyHi1B3n7aQ6swXmeC
nu5yLb2vJ8T8Xzx4QEW2m4jPF5vTmGenjHNFc79vgJ838DsdGmnCq+KQvfkJdYmCX56n1jfoxvIg
ftOXuB98xVocV0L2fcsX0psUYJ6cq/vlSN9DkMhZbFj8V0kpE3VOJw7O9o9a3NuQPWjp41rfV7A7
ijBWr8UsmwmPAYp5dv8FPPGRzgvz31FcRPgEnbzJKz3r4UNVFeK+dpm/tW6ajpdQLoVMff2qinWF
qGOBHBgBPY38/t5XxJz/7I7AMXOd0jnlYV85FcjzQU+yiOq+qgcnm+/gEoCw74WmgTYFHVa0EGpD
/RUBtJNI5oGDldxR01TstuQ0u2v80mmkCi/7kt3IUHWPKgBXuqFO3Sg6srRb6Okvwm5p/SfGfidX
wAvdHFv9BTK/OfB36rwFuMw7JgU4Kv9G7LLGgCXSBBWZLGbdQmfZ1RqCYNB8nLP53QbEF8Opjhad
EcCxzs8fGxGhTqwD+w23sX3fvMUa1IwrSr4mIjSMKqLLX+kXV49PpNmExYC4CHyou5y/+J9ZBnDh
UUgOy0l+DJapPkG+38ZAVAo60c14+NVpdpd3ckHxalyzLuy3/Jxl6Gh3vESVED+vTtlxaxspPwgt
CoJ7M4rj87OgmGZZjjVGoEptg6KFUya3keKvJBgudAt2VLbByDFxlO1dKKT/dfgDl+6HPCj6ggxu
xWCPaFIA/dj8zlySgJEVa4T7LyiqJNpetk2wIFhBmBDfDF1WyF4Vl4PrsKBmDRjv/74cCFtSOsOw
I/TSqHtBO9kmYWCecsmI0QY2iqhZ3MGreIudjZxmlSobq4g6QYD3xChwogDmFJRkUeklNoJD5xBo
ELf9noihSgkE412gzdgMizZLg5Xi6rGS9e2ZbEX+Buyj/TLQ6ZZv2FGBSjbS3zdd2UBuSf0XKOWd
U23vUsGQ+eZjA4ReOeDAhoNNVSNjowhzUajnD+rMUjxQD7XM5Kr5Gd3n8MuPF+c+6vJ5LtTouKNi
PUvey9ya8WT9tlrME3CJbpJJdFSmYvUddJVYhcX+5c11sU7fREfReoUMl5etcYAkBf6cgRT9sI6Y
D3SPPpyfk8izheRdHdZ7EhCXKDkJd8nswE7PlW9dqt32FVJfH154N++YzxX/YWUG7BOxz8OzbIqg
zuEkAIfT2CQ0mhbln7RkQ22lzUhIixhLkq+0bxPhyfe/8D3k1Sp0+018aiEXmBAymyEJUSRKrpSb
HZMabLofg9qtN4hSbPXviVpL83JD6mk5DMjlKlugcsQaieieu5Sw8f1noEAjKIifZLYZAw6xHHAX
roGk/MCUr0jOHIC2jKELgVZnrHRoVNdmqKZZ8EY9AgT+EynpqFrDiRC4Q22zprv6Uzc6f32osT0i
SQEZv2CGaaCPJvikxrP/ovQ2wj66AKlEyBkL2p71Zm6Kc2ybx4D6ucMC5xhKsRPXNEoG6a/v0QLL
JWpmW++iywWm/BNjmPHom5nV5N/u2tqB7AocWT9SJxI7s/cv0SYF/vOJLVWMnBkg1j/OZPUcVfBN
AMplJpmTWKvG1tdyM/zva99AncbK5zcNWkvq6ItYGe16JgEBgQHSw77J/e6s8+M8TJW6lD6R+WUp
pXwiM032qMUP/A+JeMDL9kE9+cHV5evFQCckOekOHQrpX0KbvpZ4WubzRKRM3hqNyBmB+aM5wpCy
ia3YECJDt9AemSqamg8+XswBkwWBPQQesk9b3u0VkQdbr0MYl/ajPP7k52PzgOSEVEu2TBtZeP6C
xYY8rsSsAy7Dfa9TqKsJshej+LjPDxm/P9rC0J7gkrh2BkD5gTUVDyB3b6dvwrHjeV3RqncleUju
Iu1NVFBQ47cgVjfgf6I1XF5CZHXx5tQDkO0FuiLKecqKuqOTViI6tH+Wc+3NtcqrpA8lVGNKeVda
RkjxTd25NgyBT+jMwr2ntBpM9MTO9V2khpm0aVx/Bs36u5zv5aLloUrb9gFjvs7BVQHBIITf+IEu
twVKiyit2r+HihBECjyfEAdR0p9wkgNFyrWo2jEeQYMTyLZLJQVo09utcylAuvS5G8JZDeAKwic3
sbwPxMbEady7QuVe8zFCKe+0kktNajsmdsWVweMauVGKz7OmTWkuVSj0N5KTE/2MM3iU4l/XS8vw
rC4/ze4a6EQwQMBaDpc2CaKsAEGL+fWCZ4gfUnLQ+oTstififfXsD0+mAfAsbQXWuvvOL5kam7Pz
+88JGDDWYTMmrIlslFhD0OhR0EdTRVQr1YX/S/4xq4v6rTVxr+doJ3Vx4BrG+nvacMkOtA23nrDY
d618z0BhMWW/GMxyAGkIdZhHwYJxAnmQ+rMfABUCO1AVfMujnIN7JciVVARzbbLy4I0lQR4ZIQoa
qsQWzYUfRvGYC46bfDkha+XU9K9VGBxalOXYpZvljwEDsnTUFY4Hw6o29FwyBNYjF/otIiVJWUe8
9tlo+r4IenSu1jYEI+KVDX1cpo8D0HO4oV5BWIpEZE+AyqMBKrzCSs+BByd9fMliNFwgriFJGIgt
BmywDbFk/Bkv6JYQ8bH8yQQ026iNkRpdFwdTOlWCHUfd/oYPFZapNT60/n8GysbWB6SP6yWcLE1Z
30wZPD+NLCGIaNh9dPKC5iqV+NurM9GIMI79lZ8D+kl9HMimQCROc2paj31c/0S/GT6YfTAeFrRE
jNX4EC9WjFav1HNmhFhPhrGHFpEoLChoUTYJVzdTqGt2W7Tq5r3etrjlzg2WVbhkscccp1Rra8z0
lnsMS4DD002XyJuvCvFYxt3MzdCCdgtpNO55Pplr0KEjRZTsABRKqMeUkdHtXptuhEfCFRbvnsZt
YN+/JQNjh7nLZn2NvZSyjR9v8ailVrCWOFuvjATbjmf0rfclJ2XPyHUDeOIQVSqQbaBV71pYy4BD
sgwN7mDROy4ibWckubcnPuxw2qlZYyRehjq2LSOqDXiDyShhZhf1RIcBZ1WB181trtR30e8VBL6e
NgiBtMw5l1wTNSLDyEqMniK0OUOAuIMrMq/Qc69I+MapUxOqyD0FB1s6BAzpy/sbA9WHI6GkgSoB
mzunLXBKco+7rGPb5R0M9sIiF+g5RKW/vVSPuOqWNoKF9Jn6dzTGJxVfApXAQ+XRaJxJYWbUw+yW
QTlVMsFh3jmPNgYqXqHuN9IWRJ2eMobeWZYDNXlfi/XtxYgF0g4SV7UpefKPHAviOS4xUyeeiGSC
T/5iuehXCLhTTmXGCENWcSwWuBgqfTcc0/WEJLJqdRiJUTzQMLBi8Lv1iB/4uV6nEg1aIW3OzPMi
mK9rF16yrpikTsgHnPb+7upUYiSKq2+59gE/kFmBRiaK0gis51KUxyvCSYCINUyshlW8/qTNpbka
oLWPkOIQujAffY2wXCKNNYwwdRiQsixszcDSPnspdGLQqohV7sQ+CwX+OOejM/hqJ+3ViBzSUf+d
wrPP+g00w+9axBWfF0+kUd+qcHTzldUNnqE2kBG+AmlvDSmRXq9zMSIOkoc8D2/ItNqTVjp3MrbC
ruCGzCW1cYh1XcnWfBnthQ6yWDMsEojVWA7D7bJop73XlPD6Wmmg1IBgFf2kL21JIbT3qoVbJoDE
Jse0z91Dm1cEJ4cKYSlqpGQJQLbBA3YZi380qg8Ve2Bq7a+PW24nAzPCL9bYdrfpUSKaodTzisDo
um4dVVOch5TIgKOmQ2ZX+ZNPwg3QHFmJeYIEGFLvO4CJscs8IVNJG4Z0VTD8u9LV1W6kcN+cNdBl
RNbbBjiMkrwlGxhAjazIdEeC64QYBDjlTPMaNsK0bjjATVrvxDkZnGnuojzMWKVgxK33Cvsf4MXs
obLGc8ir5ii3Le9Pnbqy6wCLtD69RC3+04iNbL1maqVde8hmpZEVCsyK1YVtud//fAfF71f4szkM
BsYZkuCxodSKclpwyygtaEkUzL1PJKC8FbaZiHG0g8rHbs40WNfY8bgdWZ/817Q1XwPLyMCduz2T
7MrlZfQWlvaVEUNhsBXBiWWdu3n4AkUYVygG5J3kIRhNoOiwyHstUYY5b6usi+UDgfIwEf+ZZwCC
7tOm0jmya6i9+ITXPO+ZN4nF7vwSzSsUJpc1JlsVchqWbD1Nm3FIZsl1QA3TVQMbLVVR6ISg3Dua
GD+kBjrQ8nlZ7j3g1nbBrOZuw3H0syXDExrqqOhRd/cmkadGpSSW1EhCNXBqsS/zRfYuPft7fqOT
P2dHfuMV/cM5EuqxUTDJ0romkyDlNKdxsSt8oUC6ameY671cScY7CGTVNeZTzLyKOq3T2k2gBf5e
RJNINxb5DJjgd+St77apRc8lHFPc9m5Q2xwplBpSepEBIzcAO0j+xgazGSAorWm1hgwVtSGcrFtr
eJYcsVkuqzTtxKeEBjTiIS2fcZ8+A0eWAMSpOsrKzAdLOHIKR4KNTQrk6RFuv1KUwaSfw477AWB/
WrTbm10jLpVGG46CxpoKTTP/uP8txdhdUpYNrKLVetgJD+2Wve2if6U+XRJqtU0tAQ60ylMnWgYU
7U5Meok5GKZndhVFt/Ff+HlfASPrji2prEGkVpCUdqHKMA7W/syItups8c5T6UeNxvWT2a/IHGzt
6XQBDCa7tUR6KHYfIsqbjy5OXrTpJNlt4gk/GaT6mIRhHrmZeesxKIzzbBEI8++MYGC6RJb+nlnS
QeD0c9K1FOCKGeqVqHB4VZ5NNev6E8y3vfvI+S8YMh7q1h3QKRhJJlj0QbcX/0qiTZv294qoXUSy
bLTBUPITCWRwgRzlxrQ77Cwmrtw5vFX4z/Gl+GljvJK6+xCreQIdzwJHxGiyNOfZzwrC9z3k8qDf
w4d7A5WDBL/u7qGL3ztas04DGKWXXA8dVFTom8UJhRz7rV/so3ucfu/i+EcAKOYMpkO1GSLtRrX6
3OTAj9LF/9dcM0rz8hdDnL3YAZONuPsH/2HiuvSnTi7GhmI2AJMmDbySG53ukajoP3PlkiShGrdW
NVRYCqjvx2vJGsvbg5ARaJZ5xI8i4QP6dtXtr/ie2aYj5IOQo9mcnt6+9kT4btY3Xz787fYGzSCr
14F49G8ivRzhaql0YNwgzI3Pgo7syIY3L1gCtOeM5Kc7oKzA2Ioah4EXqBlllxM+HR+Op22MqMnK
NFt4eNm/6qIAA3Gkmz0e9Il/yanCj2zzMqWbJiMFzw2wJv1t2ct0RAG6eKGFyvAgvhPDAu68jR56
9WAPAj5s6iMO6EtIYFF8263SF62Hb6G0RHnhcP3SlsBjtb55fMO1CZwjPmTUuYAiwWX9Bg8O49EF
OCX2a/kCd4wT3tuRwpTycoVC/YRz2RaVqKhJpbmFPkz4aqAfPZmXI7xd1BFRB1SEK6c5uonm2TuA
+5TyDN/DogMdYX1TaqpZcM6pOaNgCO8pJKTQUDZJIGd5/+mNy/kTf0/aVOq7ueTl9ifqnIAm4pl6
asqpvcKWku6Mx5zIAlqWgwQae+UCK+VuYPJ1H5EnRB0f9Nk+ZB+0TAHE5wxmeJWKYPBzVu4U9URu
ZzQ56FmBbvgk+Ne0zz25eGf3fpYdLEV8iwmIGL7PkWniv5seANyTO/nXkeQ0Xpa9nmsm8Mu07FHm
a5JQFMSgTOmPb5dgz1/01rvXt6yP+OqjciIS4B/NZt/kEvccJq9pceqD4HidOAJZHcNC9s1M9BMu
x68jJGiq1NKKFSvLhm2Gw9n9kyftB5+xx36cFhcigzjw9ia6R+xHKiDHLP6trHIknl4vah3WEtHs
D1OGvm9Ht813uX4ka8zJyrT9OGnlxL/cadCz+iITbdulEliK8Liqq+EwJC0Z4d5YB78FrMvjNEeg
B2Xlt2CSn4tBq/di51jmlntfDL4TaO2SVMbBQyjSEDX+yd56NsidSPx++l12IgBhK3K0jB1rNn4I
QMJ67anGokv/2bEOj+UbGs1A5ZirqYwC1W3qLPVBY7Q2QORLmz4GH85Yhah6mlrJXS0Ew7NFWjuP
rCtOxN4wb6qtxxNMFq8i07XKAsxhE3s0SC2wa/PxqT/oh4oAsn8HSyNRidMNNr1uzc0bMNBB4/8Z
OCj/dahu16yjJvKzrWQBefWzJ4Rli0dfdTr51dn0ALywTWCau2pmuIVkN2D4/VWf/100XJq/5m5p
878AhQiNR8IJXsgf2wbfPArABzVDmEVWQKd6w6BBBY+354HDI5TwvnlQ5LyCankDfpO3hBI37TZz
Chmk9e5IVtW2/kf/3kKjwxlB3fYGi2hWIFqjETvg7Ru9ixSwwDZGa+MNuFiP9FT4cCU0pRi5C31S
1VUNmKc8K0OnciUwUWZPc2ZrogmiEuK0VZMZy9nd2rPg71UF3zv6z9IqU/1XPGkhlBimjU/1Na0W
/sUzya7GP1CO+IhCpgLTlaYVgX4aaOl4xznAFi0fkBlhjVV8YiNQif0yclvA0IczM2X8n6MO/Qbh
+hl+d21tJBPgDwqIJihgC4OyMSa6EhZGRZzvPMS+atNFrB+f2xuqj7KLeY91hNHXHPCXYA9ICSNT
HNp1/NSjL+QZRPTP/zhfTEFKXwQfHRcCMxv3VeZghg4+2YUHF53uFHmLYDQItadGtu2ZalLhoU00
ufnXJUHYQwv8s0RRVcgVflC6KP6dzywd8U0MlyhcuTm9Cfc66u8hVxGkoHZFlM3XB1tSI21BKchP
psABk2yux4MhLxbLs3ELDtkfoLobluoqL1HNLrvdYfauid21dBq9DY7cnMHkHMjiEc0lxQgoWW3K
sqxUXhON1vmd2AhOPPE7eEeEeDUT20eMhP2IF2hAqDUmfTRvXw0BIf7uoPbL3h7ScwNYTd28uQNO
LbgzuwSB1uJPb6QsZNmhWr1voigLY6pEroTXUq1T6FxKW8dVwJltaOwRwrBpizRgzLcdwofKcPt9
sVHX8JPMrzd7RrCNoKxMAA66XhB6yO1rg7rVZHnf6FWHRB77hib9dq4orwhf7yzRvtaJSJZOMCQ1
pjBUfDJT4tKUNETtpeMSroaVpf5CpJ5GhEqUxjvVtSJtQ7mPoltOKz3QF6FLoI9i7MNGiO5NbPfN
AANtwZ8Jwj407/IxyH8+vW/8VU9/UNyflQA6VrlHg4c0ZFbUCUduGleNffTTOO6Suusgc6hiES4G
UXE2oE7OPkULPP8jXWrUHraaW34UKuYU4IV2+A6c60uRh5RboF0jr08bLoOtAt3LpYHMqpiUnHil
bpkeqH3/mLGSivPmqg3lktOfSNu1UlMGmN7nyTsqfUdjF8k/CDhOQ5RCRdppxZtKBvZmLKNTlLpm
k2imTCLcmnJZthcOurI/dmChvzbMy2VJU6+KdInOCceG2/v1fiU01g6WoxgBLPmJYi943w8Ibcpp
wgFfApwiZkUCEqhbNX1FCa7SnA4rWkk6tK3y7aQoo7tIFcg16hp5zet54ftYfn/rl7ulupf1tVQu
ficNpXd4fpoQ61w8RGUBYUwNoJWuTpgCSTg+q86DYmagQmEP5ypRungXnfWfFjRmCPEcS9Mw/NvJ
QF1GfDkMw4FVhJmvZSrbBgJFBeiAJr6jk8lmhwXCxiYgNMXZq6ugD1ecILr0LWae2xOorp0WfM27
/ntXRoFw0KpVcVHA3jXXD7ihOVJBnEM1zY40hVqknxN4zM+k8qKP2NpUomIzHSAQfPXsRuPj/5Nc
yZZoxZUiVtwQRJuVn9WV8KkC9O8I9e6t/qxWAffKuTQc1KGQRq3z1JenAmSplyfEctUMYXEFKGp9
ir6IgTq3wMG3npol6mm5+RpxoB9+xHilK7NcDnyvj41y8mipL53Q6jinstbUgzUjUbyoYmrA5hZH
F4LwUMG2WZuH+nxm5N0xtM5/TdffIOfxq0x4ty1lTiyDWe9yYPGvXi3ENbz/sMygG1W24HRbaSaS
R/QJ2Ma4Z1vbGyEauynKOMAkHj6iJA+qXWf2QvVxHJ+nu5qWe70k1sZhZbfr/j0OiWXtRVvAJseL
Ef4dMdCXB9xQQB7cthI1cseMY4lQcwJNWMPHl6F0wcnsgCVHW5bPKgKq5Jbs1Fm5gICHwZsrmw4i
hGe+m0Val9FgnR7WSZcGrh6ufIBHA6yOw4ROMLIxL+2RZc6ZyL2P240kaY3fOaEKWAPslv0lSDtZ
yk+STr2JTwq+8ucL7+h3A1WF7isg3QDAbi2jeoolBObwsRiOv6t0vxiQs7rXQ5QnJ3tJm8kVvI3o
jKfjviQ5q38mJitF9bC0z+KGdvIfzy0A3vc9TdGg747Lfv7wXlGV2J3emU6STs3LrE8TfyiEDVHd
KNu2VtFTgons3Z60QbB9puybpXOaOstzS1LfRr0ri6JyoJQoM6EFcxS2LW16lr6IBGduYxs0Kx6j
GNSgfgKRxE+29zR0oLhpOdVA/VaXh/Ee7FXWz1YDmUaeoN3FTfQEhs3LpmkCUvCXBfvjPwFYcIia
fFSjXbQlg7C77XzUKbGP4MD3NKrpG9tQXEZNUPGoO+rB8QQuwQXheutFrdJJ1vJO501aIfsA8JqI
WQi8itX3BmsiZDIz56sZjpnQCtqxw6GMJFi2e+XQh4AmvgCFflaCejw+7/sy5tp/k+gJWjeEgloS
SH2fbapOgzaC0Iiku0O27c7FyVonsKL66SUBql4bmRj7SGhStpc5NKWZ6KKOnRVVkD3IA8jewHEy
wT78A/4n0vwzGhgJuAQy9V/pXJbS/rVT2avraQDUW/EJReFV/rIkINemBFWW3gGKH0cPawmEGxfS
UYDl2EoQhDNofXJA+2bFLiAY8ps1hLO/6enOMBKqq4vUFT1IYNxMErWwNOen1V5kOxnLA/P1WBla
vp/1uCxo3D37S0BILI3lv/gGjslv7arIEN/knMJMkYHuMlZi7HJHSynw3brfV69Dw3Phn9oyCkCW
TE9OaKoO5kbDxzUcs55AfitTXU6HLzsHwam1cjOLYNJ2NXl1KQdBEU6xEyjSbLnTVA49idcNJsUc
WXsu7hKs8bMUC8IyuvM0gcYsFwnFnBDl5q9R7CKjRaSV/YCMR2yaeoIPCjWftsxFwaHBAADqqI5E
hy/7bhaPzR9iA7X/6IYjudl0Z081YsUf3LlbF3xVRwkQmIrokpelbWEcFPhP0lCSdiFl9ZA/O7lj
ChfiZZovXuU3/4keoCkvfDs5oMclHWoqhWeLGUI6cRYLNMTRP+kfYuk5jGvkTeb31BJfjF93rBGF
5Tk6aPlec1tCGJc9F6Q7PjjAkR8/K87//XlTaAZsLZ5PnHgSo+sUh30yhcT4tQ4ctVCS+S2c1oa1
xO+Auxl9aetT0T2JsDfs5WwNSzoefgLvCi5BQ6DRi3NzVWWpZbuF/bcBVHEBsN6uPA1+htEJl3uz
0kJ/m590xT0WwdEVlGw62BiN9qGiIcZC+xP3bSWrZ1eOCNN4F3uXcWcoFSY9rnjaHUuR03I5m0A3
IbAR4/r81CBp7TYE85MBQ1fMMB1vv9ZHyjiNolB0mqU5b2AzzFTjExiCdNi7iib71q9MnpUwWYy2
YY8G+kWzXOSUKjM1mkG/nPEW5zkI/tEzEI5xBwjoVxEgiAd1PUaywyBsXY+UsIjodxPtMQbfUHQ5
4Q/NqnqyCzB7mir1OMOocVv3uogPSTbvsY4RKGzOYEHXWJHoeUnQvira1BAtVjx58LbBYXdkkhnp
ccb+ixMwtW/6fg0uD7WEVF6dNXN7sWOiShJv5KdRHYLA3DQwS5Ve4giJJQxzBy0zcxoNsMok8kNg
vuVlSNB1JRiVudf3aaItA2sMpSOolShjQMSvm9RBzJFY9GkBebT/O10F/V3/P93sH0ssJ/IQENRL
EHL6JDydbSZ0+n2FPi11DoRHts/EmG3TTOpMqRwI3y3mKFdY+NoKhKn7grse1UC0bPOGQYSBlcq4
DvDDc88AqV4M9eXhIr7xsVn/NM75Kib1k/0dXyPcCfSHlRtMaK7DCWb/R9usxW7+1tMHSiMKceGf
DG3jmjiGtYICrRuShvYKkgrg4uormvf0nVXqUu21huQu60Q9MwaC+zvECoB31alljRDBw/2SOUTv
8QwJzkUIqS5VZ5ie5gyMBAo9Y6Rn6Jm1MFfrKJE3nQGUO3EGzwF53Z4bGH0v2sfeV1qLIsqXai3P
L+BAUuovOwNYA4kkyz1PWnLeaLAo0BvP1WNLJ6wrhUkRFN4EaRuFE4ZpjCaPHhelqSYQa0rZxAkI
b+kB7QTzCq3Ib/rxEi1tkRoSUJF5qOPgURepdsWDXyguJWyOBLHXyODlIW7Hh6ClHNiI4EjIR1cR
j4pq41NdAQF7qfVIry4Cm7hc9kIN/kTVJ+StAqn9oZfoT/+m3wHle27kf8GifjQEoF1vfX3ynOoY
9xeC7WqlZUeFwIUOnIHccILJPvtSrNFWuNcmvxq0EQpiJVmgnV6IxCfpEQ/o98DThjBLy6oavr+4
ato50+YDHxiofc+A9Yd1ucvF8kVM9aLMwkJWaThQ+D3Bb32oCNzqtiVGvmpUpxhEtlClpGztL5/U
HgaQFR7lr4abWdDAiBcQLcUlNPoboX1rzD35ghduXAhtPu79krYQ/BWkuDjaL8X7ICe9adz8dIJC
8rUuJoIO77vLCuCdtWFiD+D8VPTOaOcOmofoUKd5y8vpreMzKTJm+CUtC6jZ+WdRR6io9iZGrIbv
N+g2nkrZL+EhJ+5NBz3YNOXAn641ks55Oe+lqQq1877179CTxXzHrE26i1zp4s4/WudGnHemvYNw
OcMmP1+ZpFJN1eydgNC/DgdDsGZodJe1Vy+WPhYrqFUu5/GaxjuY6hQItNBrYrQzIMT3la51in8u
Vj27EVvU8J7rl+s7m1SO2OvrrZON8PuJp8bCBYKD11DOdwwJxFc2d7SHRMU+mfnqi+o1MY33b8m/
n2NkXha15MdQYxJSNUeax8feYIQEOBSzmTCdHWFhDC2tW0HNbnXfIz+n6l9RvZCWFGJDL+yyFRnL
ufEngWheZuOSS5Cmi60rumDj0swVveekfeygKNvgcVBLfcdyqZeVhj3N0L611SmK5TA2lZVHPHub
zuvvVyq2zjpEbqOG8qsgt6eKcze8cRRqxZJ8/uVW1ntq6bxevXm8b6hc0Ubnh07qc2v6eUrPA9pC
5bqDgewDdcBjeL6+nPufsxfuy7CaOh2k44txMF0bGOCarg66jScCbk+yRPx6xDan/09LnfIJMyub
Krh6sQ9rU0MWkruwll82eTe0lITMel69Gf/5clPuN0GyEw8qBnI7FvK3PmV7Fz2b0qHzgLBuuKzT
7dUuUm5dt0mknIVo9EGcX3M0TqBX/PHicnknnGoHps5ZxpPHSH2Kpn+9piUT5Q3WmxD3KZKrRLuJ
74ad5erVI7lb5JmF5rc+TOmgs8oJeLECK3QgRbUK9e7yExxqOnyTtssPj9tmVaR+4ckitJUjY0KQ
1vMV/8Y2UUsBga/tMlIM4MQhToLjUYKsLhyb8GBeI0QHF/Dl/xNdceXNfmj3WBoy75W1thig0oqr
lY2uOGMB3U3lB2dF/yHi4HErj8Gd8ZZ8z/SmBbtc6M8dW312yZp6qHTa37nWNCTxsK4canWfa06e
GQhNRWVCzF4wFtizDE2U4o+h/s4XVkrIYpoe5BIAcFf8MW9/kqe4gpplqqMR778+xKqAYNPqMnLU
HP5XXLTZI9Et3S2fZZ2iDbSuijGCA1/X8JmzVlxcfCluVqQFqr93TOzvtMeH2uw31vfE0PBmJgRu
BGH+qoEFDM2KG1RDIG6OAHbzgSCHsMShLi9UziB77lCjn4fkJbfWuL8aGNNh5HwaDVbc0iNKz7Mg
y+2jQ/tnviMC683Pt8qLz5Rg2P937bXUWe6tNgSUTS61+fkBj3HtC4V88xk/KjKOPKazY6mlPKYb
ornB4ucwOKkLN65yry5+qoZfraP1bL0JXl0jzJAzC5mXisABSZXNUHu67jj8CMcRyAJWxPG+0o0R
3+kTzu5tmwO/oPgEtz6E9JPcle0RmFrYU9/MqUpi1R5LQ0NeU+/GBnm0fpircn2nqk9omLCq/vjN
HpiCrVrz09RwLHpz2/IbG5HpbptVVAB+Om0KWvu5fF7xtHA0UGzHg8ltwiRJHe8QfU6OgreTcvHK
BQl6hwlyxSwo9v+egrpOzGOz/28edaufiVO0Dg48gi27raz3crML6PSa8W7HcTZW24g/8zOrd8B2
e6ozeEbigRgdm9iVcHh+Y38sY21GT486V1ZSHF/HrN3YJcz/aPAjDNmf5tIPWbnfNPKFNnImWdi+
kJXxtqsCj7ha8mVXJRSdhfoejiZ7OEZymiPWfgZiGlAbC7mzvY0t4xXetH/rdd0rc2165lwkruNJ
YkUITlpy5As7WNIkaCw2GeFosIrA0pu5PHw0Vep80aD8Aiscu6IdjMafCzmQ2sdl0JUti60ubEl+
hd+zEwz4BUc0NZ/Am0txejj/tFWcRvNdUMhD0RkKjr5Wit1qtcftojuuxz6nQAlKAEi8ty5k1VVB
dI94d2BrVF/9pO9Dji88m2x1aezISEf3TiENQ66vhD6JTjGf9Snc5eZNglw/oIS5Q0YD0Qyt/e5p
omxTmbnW1wz/scwxfAgDejn5IxR6sZU40gzj/bN0pNeUcY+qFc0ZA+Lew1+1pr5S2kj8fUL7E+wB
yr04WqOhabBBjefjC5y38V8zqC5REXK9O06dFuAawHbOIEZ1JhVWDj7hHuPTRq7aDB/vyZAMFYro
K+TrfiVoC4VAM2nZNQ24CDVKJCSAvOnOZu68GAKFWV9B1aKqwr21+/fcvDuBQ1ThkEZAOr4oc8k6
aJlzjzebu1U+dOP+VjLhw/ILcjeNZ+gfVrG9wsyoHWr2W6n5/WyBOtFlUdvcAepPhSewdCFpC6CK
ZR4kuP8Ujce/0jcz48fBSy8S3lSXEdD7MP13ysUlCQu67HkUfO5rLdZyNQhm72L32OhJu3jmVnzT
4zGeNwoNccdpt+NGT7x7tBQ5s/Z9POfBArwNb0YaXyZkODzVrVo4S7syqy+7JT5esbEWSQKCd90u
pJibtzPSFVsk9V8wqY06l2mUrstqaiVIq6YJQtyFdlTBCrrkitUzUfInEkBhAiMhkE1oCpoW7IbT
ucQt3auzKEaG/RkL6dbkkjfilmEdDq8El/oiwhTnSNtFdemhIbJBVuS53ue+aZD1i4HdtUdz27g5
QX+cF3J1NnClJagzLOu/CYjHBPtJ2gqF3FSHh4rIJ0ea98okGhCXFg4JPKUxwtfeC4mUfvtoJJk4
ZP8saUVoZOH6CQVBNRzGuBptoX39Ck35U9ZFlyvif1BGf38//i7FfxM9YaJNESPgH31SXRLiglfV
/g4cj0mhD/Yzizb6p6F0jRjTuFYA64bj2sZCsl17q0zIHyTIPg8I51EMaOjj7Vtile2kQUSyhmHe
xAeBnCZhUXgFLT9HALiO2/WOAmYxfgl+5L63dMOY0V2lHlF6JD+xkX598ZPgNx0wfhLrp1QrxDVd
DLEt9aTPjxusddgm8BjBPsTnwkqcQ0ustu5u5uVxBCShGJeR/Vn40zlla4qv51jfoiDJysSquD9b
Lir6hy68xxZgeygw9FIKdyEYB9xffcUxY+o58LZk9EudELMpIDykptcmWmrjlhyvHVDPSACcxdHA
Lxs7rHOvA0DDy95AU+5S6u1/nhOLaxg1aNW1KmdBz7RKSpBDqwCBv7/6+7S6Fyxx6QOOrs0PDcsj
22BoPjDJibBekL8tcz2hqfCsFUJxcMJMvGwlvuWRrkApLh7IizF7PsknYMQkK9AVAN5QEm37tTuM
N55u9pgLcB3agSMHwo0EdPDrIR3zNLIHYPqv6O0Vvfgg3pYTnwbZOZPJ2eMO7lEQF92aLA0d4iKm
X8be3LPvGo9Nm7xQjpWCh6zaEVHseLaAZhzV+pe5yt3Lul5k7cYVT1l9/2HvMuHTCJzd9z1qa13Z
3aG4Fjl9PlQyBgir1O+RCT10dbv7s82xrtdqqF2jZf0AHBJsM8+4N4YakMngXIRHof25xFCp9Z/8
soMRb4hELvCwmsA0m0Wc8w/kUFejDZbS+ezeuPUIMcXf+xn4yLMvqcJBj02nqlO2NZQYXxIC43PF
h4wGbYHRxYs+Rf3rpzt+kYQ+gGCPfk5YrvXJXB46GEtzWIhl+D6hc+lJuD40dtF9WFipO8ud+sZg
4QcrP1Mg2fjJ6Bgj0u/eLS8VjwxaaHV5LIZH7Wa1v4gatg4thFbsDOMNJfp9xdDO8m1eMWXpJ5at
34psyYadxqaaibC5TUHTi5DRn2KoaBEyqNPRslizt45fM+ez9et6VeenGm/vPSGYtwKOG0747Exy
GplMwVCQvfeCPBkjWIcXxp3u1iw19/FPoECeEUZiEGDTwxJz8ILfiQ36Tm4wnOxqKlwqvwoM3iQq
l8EpufvBq+MgemnIOo8jZQhMQ49ZYaULmh3+vYCMiAtJUbm5lv9n5gAgERLOWGJTMn4QbaOYAXCT
mohrmpqkhANVzHbvZ6L1nKxeJGRJT5U51/Vjv56q5VZ27prdez8sxbklEd+nDaYDZLfcz4FqIqGx
4xc4K+9Wb+AWk2W6y2sMZmaI3Bubxh9CaZi/l9GLTbmreEWnbTdvAAN0qvISjGgaBTUZJsWioh1E
o3vDjOD/ni+daDExI/3hQR2uGdKJPDd1IadDI7H0fjSC/BHK7cuvw8sUVb8V8seMTcoqXguGt3Dk
YxACVNuEPGHjpnTYQgfVOwZqB3xF54iJNaYNAz7mTbuOxkdN75ZElxwiapDW1hYO1zGVcRCQ2t6l
rhrY/iD23hZgEYMibt1YxPNgxosTUhcfTR5U62u39WWLzFPgVNhMX6oM/FnoGTPl/dIW+WupAjgB
bp9BTVFYK4HzljrPlC8XEoNi6W5zWNwbilx/xKeSA4W+y12VXkAGvOE5wcwiMQZEM/Lg0ivfTr2x
mzyG46AB5UbAACYkhjO+1Pn/2Ny0SpTV43mz18Er4NO4iR4HGKfoSWieuqOqhkm1gCSyqy0u58Jc
e/cSsnXTvYy9OISs8fTls3ziGfcXA90g6XkzjDQS+RwH04/fGVCw/HBRcuWUlXfA1Mn9E64/UhCr
WCmClDyF20LbG8V1hx+6ob/NtQXdn0KgvmvgHX9Xa/0ITC+j/73WnniSWyl6TABf/gVFGUchiIwe
BHzksjZ4v3r49PLFOiO2P8fwGQs8mXa5WYWOVS8JFsI4lK1m871HGf3I3LZ1fINwVCo/95rrNp3v
3mBz5/xsyISeF0uj+e7No3AhyFG5WTc8kFpIpJuaMgfemDWDHTk2YhjKGZg9b2C/VIL4I/YmRkoP
E2t9F6D2CgDAu2TpY2eybvD/vb0TbcG0xmNjMgTgqnIC3U0s6t6BEP5lhRI0ouNajELAnkiR0BZk
czSGIPqFdxHkS7ITR3oxKPGQTmSbY3GLIuW1LsmeB5/3No8Qlo2Zy2E0Jjt13TbH7dF4/g9IAnbd
Uwot9RFyNZncQ/ehxyY8c2mhNDIiYVIwYUydEbx4Lr7anVr96ZR1KcYNS8i9m7mLO368dW1LMAgA
nIOzSpq9VI/coLUVzHuY7mK42aeakphq1QtLeF9uFBTrHaw/4po5todGSqolxHuhU955i4ffTfSF
UEBeUiNZNLFxzYph5TaxaFnH9YP8N2JlIBIlDJKF/WhGdalj4UAzdRWym7RPodcN/Et7k+w+uzm3
Q62UhxKBoZ6sFgHbRdUwr/7cxRDoHXF8eXm0w8Xfk5xs3gdsY2Q+6Q7prNQy80fEjQOG87++m6xV
maCguY1ZtWI8Nmvklu5cpzgNKuF4kC6dmEfUkMCPxNJmZ7THRKBZIZmitoPesaSPqdB2yiU1S3MX
5u15PeuIf+RYZjp4UJxHc9IY54SBW5pqlJ0bF9KKeI87rCoSt1lf9QHLzl2xRLzPeTD7PlODLHTF
0Fpk8Po1yRuiBFUVvw4GPOpBjBvNZp8HuCA9J3x/0k3GOtcWRLzq75WHW3WlpSOP+W80qeqHRXbc
0v9xPrLI3BjLlhLiYsdisjwePyUhKz7Pte+faTNdHQI3SCbVG0r+amJxN/6U05KYX8/PH6s9FfqI
XJDAXPI24gXv8r/l1WvAtM60whkCc+DZ38deI/JO3ATppM1bG0OiV91mrYjK6HVwtiKNjvpm4bcL
xX/96QYWtXr6Jn0SVeZWnDYMJhXzSDYsqZ6gHdToJkF2Lfn33Vf8/6o21hOr/EbrX0hcpwOVNiSy
WUSeiCnkFDiHriomlURLR7jqt5xFxM1WgTJrG0VEAIu/Oc3rIXumta3tx3KlIYDBQp9L9MKzhWC6
JyEzO5ulBCRbqnpzP8ihhS0/RNSxArC0rTeWv5YCvdB36iqal0VYtRATfxFmAUdiHNhoDRImqLZS
EqgQvrunEhH5uWPSh8Mz+FcUdI46r+fj7ERjqwuHS6bxEf2k0/RfeUvksVz+9IsykfSdVaz769Bp
wdrXmP/ZeBa0byGoS1SraSKIeOvufNDcOt0DXOpCFzNf7k2ue+lgNN1aiAbstKNqEWkShGbfNi11
IZfwCiIfzxd7d4EQGGU5ZY+XQNDRyzRPf+xF6sIdRBa6ENQU7m1sPZBWhv1oCy6YAUuoxzxQs5iv
bEC1yMU2Nzg+d+GSVNZkY+UelN8AqdTwu3sRvgcuvTgsP/PlF4hA1grWkJ/edB8dKwzIpB5v0HhH
cGO8U+aeZH5JSOjZsNHByFjRS1YlfWf6BxOaDtFRI9XsqbyjOCHEieaSqgxfS6koWz8gKP4WuSId
LUdUcOAoIItdA/Brivz8RxZu3s8o3xDoHCVdT9mrf5MqxDrEJ85StXGkldkBQ5Ql3M877xVvvPEi
HD99ZjMvt1xLLeJ7PI4zcNDrHH/47Xci+z5Qx7gg2tZmcXycp+wrA0/3CGTDGPWjpXVldTEd/2RM
1Ec1TFyhmrBBilbnqBwaGf7dU1wo2hsyvY9NrXz+FdC5TyR7mOkJq3EnBo9Ehd5ZWSXJwGLzBH81
iNA/fft70OlbkkXjz61pQ4RYbUHRc5kHtwPrgB2Hd3KPsTM+YMvgjqAfZoL+fp8qLtKsRwEGro0t
oDlOuq4Bpz0kuiKnajsVHS953tddwDRxFgU2gTcyelMClkW8XqKbCS7+Kh3+RjiIu1o223pTx8r0
VbWeiM8TRoBlsIeu1Y57xblxNLdCpZEKnUv3Oz6wLy0V+o0dF7qiwoWqr9ZgmK74rQu88FtJsNqF
8Ge0OTo9XTUtYJcHVClbsm+jXu4s+9dLkkqRG3iSuqtsyQd+wvT/T0xl3mhSoI9qJJtPfGZ5XSCK
FdeirDcfzN2g4YB+/XB/HjQO/pgKgsDcudHkWTQcn7Dj2DEAnBF+EVJbsnjwgb6NcgtZbJzYMiUw
LiD1Cd4YIqL9C5TyMfOo7LgV3K3x99GghXECZP3usANhqM+HIk8/ZFqaEx5aVUziiJJmmSFUkaJq
ilAX77rV5P6QXb3E/WCTdMl9MhvKIKO5FytYELLqxNTYvJ8Kt1IRLUF+yAxz2hO6f8lOkhYxCfDm
pEY1l48bwfhjkNLnivOs4smuTBxwM9gVk+tJqKD5GCn7UH9VA8sVzk/8PvZZK4IsFgaSgXKGNyhh
i3VCocyGT5IhXZ3yk5P1t6sjbDQBkK7NbUIUBhuxND/a3s7evi6yQ469wQnDJWrQA5+CO+5w5wx2
phrbnxIyufSztH/mmIPF+9KgqCt+rMH64S1jTJ86LxU4PzK6lambDkAa3dhfTRRxpU4VSSvyIomg
vzKXP2mauClhKGZ9Hrz4Gc7P1eaAuBZNNzTFquSwJczrsa2UXhHbKi4e8p9ssCyXycLG8Su6rhio
0cGyf+15mjQvsu2IxDcnplIwdTAwbj8wTwZJjj//SkQE83DtYwPU3yScqwCATgqZAPWPsHkJEtnb
2ks8DjoXjpdoyOn4q7QNP/9JIpXsPOodnpT5Fztfca0mgsyFVyvaZgaaXhKj5AqfARtD7bZMbmk8
c8kRLxKYGvYG0IAzhj4l7ogYyZ50KBlS3PBrLf0IqaDukGHabeGAgJjiibC66FaFqi1m3JpYxHAx
TBC6rH6+REj6H/hvqPoNZe+L7mnJ0mzZPDnU/Be5Xil9egs2l/FUK8Y2aliZ/gH6gwcVU4O6M2D4
Cs/s4t836blpFvBbJBsWlz74aDdE1vEuXaziqX+vOnqbwLwtGSAvWY47i6CNqw7j8PK37/UGOSzY
8croYL+cY9zhZm1Fe8WHmG3AfmOxoP55W611B037XHoIXdrVM1Oewn3zLGgJk6yDt5vlv7C4pE8Z
zeb0EM/LIx4gFaHns72ay9AivjKRE9zaIfW2LeIHRabVjl3ipAGASxqfwElfov1P+gQYYlcD/IFS
h3i/EK5zEbkhxsEtw8sJIbv7QPYEwfJAUe5F0GBUyHybaOMsV5gEARBbyzp6CLSX9NNr6/M9APCO
TRT/VdDDrsL7o9i/yxwXfJnZNC8TyVGTW7MNQxAIgNodniijn8186gSY3W3DE6vzhq443cPy93y2
IIE3vIlrJs9UeotAcNoMzjrXFecRvPybIr+m7WIe6P9KZvOtdQqwm9SQZARa+/RGGdajd0K9f0cI
A4MPl9wil7g/EM+bhGiZihkp1thuzl0TJYaX9AVPaLuDoW1KTv4DL2F9NSP8Lt5aD9cuh2Ke6V31
BBj/lL3fxPZ6+iLGxDKHHNz8Mv3dqzFDlxhMRq+lHw9E7JyeghGsNsk+lPU9/PP7AjEADcc4atti
LwU5MMu6JTGlpvx1xsn1Ercy1w/roksg5Xy/IvOSiiUzcW4809Z2PMtsgSsNNQNT1V5XiFyMOiC+
XB38TqHw+VvwUDOvq1TfCxdUHWHftKIFXTXl5v7+EALQ3b4AQU7Jy6Bvry+lEceq07Lb19+mIqo3
gSFehnGtyZgAwAts8Se9caB8bP/ifKgMElO+bkE4gSBzuIMMwqciEA/QeVq+I0W3SkTkwEg+LtT0
ZKSqzxQazn8Qgcsmyw4fCw86PPrvca6g5W3qbwTxkW9eCEweYkX6LckoMcGw3GX24eVsc76OWlga
/ELRKwZc8ENdEeZHTqZOm6o5w8ISW2lLIeBK1yof1E06TL8Q96wihWaivY251SxZz/McQfPsOBKB
peCL1rfsKw2hFjogxP1nQOSJz3H0jLJ6sqpNph9FeTwHUwl9x2WwVVf0GB6EffeJ0AyHjLyXpg24
xAP8xam5x0OtYj3tleosf1DX9ufxNUQvCLdltejpnu93AncWcHqgKx7s6HdLtWepIdHcFAKcUzc9
Kn4EJme+PQ7i1Vg/WrM12IGFB+f5Bb9zgmhUyvJtseiXmGMKzoKT1SL2pqyUeXtw669ruJL4h3x6
bLggJIAU0Y/HYSMrjZPO7jHggeOOOabtB1Gzv4ZcyBSHOE244BmZJ3hznzdpcYgCKPqOH22cXPUz
K7klNybTZ4UGh59Cg1ET34Q4NQUmfj2AWQ4hsjLD44yuiPmaAsamvjTbdpuaTj4SUyZmzSp9KDBD
acdDOwcDJkQ5WpelFP8bl6IlmrtRQKHDWHKoZHoES8A17UA/drTH1PMU9OmIjxj5t8cB6fFdLyLe
ui5lcndBOD+D6o9EHnzjLaOI+4R5Tx5DWwwWuW92Ny37BPJlXI2jDLBamhSUmcNV1Zkk9k6CoQ3O
suCv+Ytoa1ku4DUREqsz0ISllJyIL1FlgMhPPefm/ek6J+5bUV7BwhgWAgKdvrLLWvKBR4g9gJtf
oVcglb5Gupe14Uk+6SV60TeXYoTGrgxcxeI/52FYD8262rJ4CW8HPzGqBeCk8SoUAkMir76d9hNB
DFXPaqBfkyoU7izkVyMkgNDqYwRMGP2nT2AraLAmIUfTpzFd8zKwZtsk81+TaXKITY0my3gfgGNQ
nQ9StvGFKrOFNJi+MX7d95upJW1FYJgF2EakdeplwXVlwBdT+fy3Bl0QmzGwgJKMERRCwLwu2Ea2
p0H7sO8UcO8APKuofoBenOTGGoca6h+HYCopFDtBEM2Vmf4/pC/JBk7cTgtBy3+6ptXANCyt1syV
60WoROrdsZNeEV9oIWRPWVEtUNn8fDvt/oq94REu52EF8HdL0oK2uhRJhT0TObfMLSycfUNQxoKd
4nai4jA3aJZ77K+u7lm0HpzrEtzlNKOebB2O9ZxS1xm5OTJdBKg9L+swweDA6wMFsgdV/KS/rGAr
D1dVErggIdDAlztlxJ7nr4rUGzotN2Yt+/kQg7m1OUxH+Zp+tiPn1uvXlYt75x7QW48oqdEbBFXZ
VfX2zSOA93SqzlrQ5lLAwn1+qmFbLmpjRXkZuLxpxV9ZV7N9o2dfoqeIsQ49KxZQEBcbMZRQTdZK
99TCdtZNwvuu0/5EyUznWNx68+c/+UHgrg5Od5pmz3TSVCR6DW9IywNymhZOsSif61LyQs1sRnUB
Rp98Z1oiHhl5nMfJMqvvDpLXl64txQnC7WfYX0EnaaJ8AWSD3kRPzBSE2BIRpY5f38ukKmE9dMFm
Tu51DeF6hQ21To3H8HnPAvi3eG1l1vRhDGry3yRzOR8S7gWa7DlI0/1qxy3G+cYDCA+BSIzOTDIn
M9abqe8vJck5+XgR/MzLBhh5ZFIhAr22TbYxRWnwr8Tc5ssfINFhElvBTn0qGXfYDTSnq83MlaAj
Mq94YqYFp4NyUfBcUIUDNGfvxVdLFJ9Wyri6HTvESzyihZprdJaDJ4jr+xZHR+8SaVGcpoae1HrA
CbolW5ejdG5GVlpzpxIrDW2Bi73HCXlQ8Z6MdnLgvVc4EzU4P+fR+a4xF/YDvARPzeeAw1vE/m8p
AIB9Z/yP9Mso7RwaHJeSSdjhuZhI/HrIBh4nO/uk3lI+t/c6WpHlc9gP6VcHwSyE9zwLB1HGGlc+
X8W12kWp28Pe2W+z4nJQaontc0i2P6hMrr5eHkdY78iWjYbZj4Rrm1aa0vkjWSSyHJlSWAZZSUbC
yTqjvIW73LLJYECRx6X3gIdz2X28V5ExqLHMv1gE9EflySw34EIFxlXKD/Jy75emTvFHgdS6AoW8
lVKRRtf8/popro2TY3WtTwht0o7AqCIkxdPDK0g5kVquMoTQMEgn0KyzEJV4bjkJa8a4ORoNJkaN
uzsT56qackF5U0iNPxMAm301es+DdwPyUCK+iBiUXrveHVdjsQHu+SedZBeMkdnDLN/adY9a2zDK
DMokBaJvIrdyCi9F8U33cVZkGOBcurDIXppG+5Ew/t4uIpBkYppuVsDvNbSg/F46pywLfHZAJmwb
teNaPjoq0dcSOaiBqnlrSFWRsPm8hqY1K1FUbwIab1NBaZ2DYuPpYkyYyH49zbs12+BqCiZsJhLY
omWbfpLur1Z+CWK5894OzsqO0w11y/y5asjNYbLlgo8QyHsGjBesEwbtVU5+ZOQbWxX/KxqxcmJh
ZjOlscnGPob2VJ5kVRA/tgvUijaPfX7+5e4CJUeqYassnLCUKB4j841I10r14LMdpofFBTSbWkYw
WJLNHqd7uTBDZzHc7SAx9ASiN3BvNdtUq0b8cmUoCnAIugqZwfNFmyNYwpo/wfwCqEt4CtLPLtWW
hN9c1SEyoWX0+hnZDNNVhwLRb67tUKE0YBt+7qfUo1CWh/wn1sCGGeybrUCROhF6G0el26njWSVt
yA0ZkZK2zaFfoNmUtE0bkKdKsE1ChyJGGWDtcAChnExEcUC6QgvR8sqMU2O4Yp2d5QgW7+Guopdk
bCsp7f8EJIcznL/d0CkRTfuFIaZaWBRSH9nLei6Y1h6bj3i9NrWQkA681MDx7E15bTHrs5MFYXY7
uPkuZPnjBFYf5rzDNRbB54VakORCfwalJzAai3CxMXI5HxLlRHxM4aTHEa3iRvYMD75r+gKbiJrn
BQvxW82QN0nxO4nJwL2BWWL4P0MIUkFN4KBLm93qzswmIrEToTVTBcpri3TiAT6nHnEl4ZVOPOk+
PsAI3jwDLPkGgmVqy0L4sA2/47WBtEH87Q/+013d6CF7GhxV6d2hJh/QQnTvHh5Dim3uwQhxSoLw
UrcF9yx4sJYFvG5RM5SqBPDcIpuexgPH0DKShaZomUEAgl5usyvUJQwhLY/mQCWx9Vn83MaZVKu7
IkBWE80QAJe2C0ZncwIadScZCEAwg+xJ33o04oY/OgMuplQh+iFbSyoRNoUxrZkCz9xB0A+Bg66U
SBQJJGtnmzDMu5O4S/Ig7m73oOotk6j1Zu/xZK2tvF9WM6EadKUgwlMWeoAEcXCO8LyaxV54kx7C
YU19CDUbhwogBl+BQXztMGvfeQw7RqG4FyUtTQCoImmZIQsIvZ1gdgjE+MFxHhr+9lGiAFwjUo92
B5K0DUdsyuoOwbaAAOGhdXOruo6dwanZ9z9c+33cF+AygiRdaEkaRMIICeRazFN1pZkUy6uuWBfD
NOMcjLog6Q0Xd+yQAStPG2FcF/AdBG9Uq5IAk27GTH8SDw57otWF/bhc/JKgb0Q0Khb9xS3JtMkQ
00MfM57S62B3cElG+MHVkMgf+dGkmwvzVqaZD5SpfXSyipi5jpcFDvvzypwj5+190HL+GPZFiZH6
L+y1GISJkDWcoa2hFjo5TaUxEV+nueYhIi4qY6hp81jXLcOjgf7yBXDIOLCUvGGrzKzBWIqU281Z
1BOfMupCP9fuMcSmkUldsJRRfV9OwDubgXarmYzJ5UIiED7zRr2JOPmeOSVGaToa9Oh3m6Vo+zWP
x5BCh8BeP7m9ZBAqHgfwyGVvPWg4YiwMFuVrc6q839nwMds13ovHdz5GJGVLi3vBlUubTU9E8RqM
/3jVFg9VupAvvC9ShOufseadBGU3LT3IFLBEq2ZBXDnEJHjykQKMUNef0l0uY7aCI7Jf9Jk7lges
0iCpV5nYOgGjstGpGwYwkPdXwHCJKZ10D5uema2mTBzSXMY8nQ5T4b/DKtvxbAQrbOwLXDJKWOUr
aTOlz64QIgnP92G95NSJf1wXneghzGQPiTBHCZBSsZoZIOXGDAjH2gsCOCxpNbaZFJke1fXWMIYL
zFC7XjWLsby4Y4sH1Qdw0eSuxgAuRmeMXWYDHxOpt/r+io8LM7VY0Rut/pMnrdmzo/Y3i3K9UaH2
UTOAvf+IRa4h6mbxOjiGvtg6Ev/gUws4xHLl7bvC1OSU1/da+uemcfmMVVFPHowH4yC8TS9O9uz8
xkYhmn/bKyUuQoOFGKOHfZbQZF6sO+Rq9wfgmR4LV7cINtjyVmYVw6C5kxeSmyTBThm3ZKLdm2aJ
foeTJqGl/4i7IBQe0Q3mrBuwFpZPmuz4ADrXrUu0FMCNn8vbY14ZPjsJEICGrIO+0VdAbjTXRRgu
A2XSxQUf+AuYhisSsVLeSpufJNLdZUwXtkuqBesf93qx5UVDJJDcbDgcJSv79IQ8pB0LpLn+0yrm
K25Ft2dwNGOCNuXi2TUpzfCBKg4/SEM4ekiK+LYBXKYagMgMWuHQPEY2vHF/asQfGYGnRrDL/jlZ
n3cRwmFxsvzdv1WxOhZYVn3i5kRoualcCfeEHxHKyIABpW6Dx4N3/kxjT+Cqg3Vn4YLX1S4PROmz
NZINmL2fP77gzFitiBQRRf2LmRn1CojIgZQ4q7+kkPKwpGASSn1LpCk77+dzoM2gZUWaTQP0Nsax
oQXxBh4UiMWwSLp0XPNtKopfAhexhOQysrJWcSSTmGumPlQfjsrkMHe8xEK0gu5tvmvl0ZrcN84W
7BWiWlPYAPm5tX9COFws3Dnq81xMWZGRyRhH3fhe2XXKfygyWE39b4dhKgnfZ2Oz3Fux0bTW+864
En6j2NmAQ3nxeS1wjCSKIm3gWQ/3yl2bp3RwIoLs24jAFMVu5AKmiLrTq16F6B107Rl2ypPtgUN2
AUtDH8U/UDDD/A2EhnTQlyqSadoJl9D18ZIi6XmBK2uu6Hryt3FmcqjYeY6CpIE9wf5r+MpbF1Q7
nlBP2ir/CaokF+SiZgL70j4kvA0LnV3Uwy+r3gW+JDHt+AKhmHCCvSJMqtkM/ZqO4L2zgLtufdlS
xf/DUCQ6bUOrsCHRYPVzVbaDz3lNPfvWtcB0mhvaAPhmDbLh0I2BGvnaFvGRBE7OKak3NaBXuM9h
XvPFJyhiHQjy0Jj06ekEjG/BmJn5MFGiNx1gLpnMm9+IcDMBwa7sWrmJXvBjxAWJtrwnQy605i7l
hskmjagKAdnlILGMtM67dtMVThuVylNy+8FVvG9ipCMeL31fsl0Z2jqHv2buGzbN8p39xsTUQK0u
5EOtllcVfC/nuxJa2QLehcJP+ROCkpEX33JUHL8DHr0jWxnlfmDXVvNZqDksGG7QXW06rG3nRpG5
J63ivhreR3QYWH0ujTvRhXgYwzriTZoSnlxrLANrkhvsy39O1a2hXdWbS+PItuf757t4+qKZuvfv
j/8V4mOvTPopp96BtREzesevsuh0buJDWOv6dPGkH6muZhJqfbBveXFoTFpMBKjRa7DVrzn6c1jS
jPSCyoKBTej6m+WblR4Im2X8UF99oru4/oH4dGItIsFQo80YB3t6nW2UsJXcBfjpYSz3xK50qtxc
l6mloQPLPyTEBsSTwANsvasc/gWgEmEvpMOQ533VIbUgRV2fSJK3LTw5il/sWTOqkmqE1yVWuvt1
fInev1S1Xeq1/KdjD3FoAPpQNbOhcmUeg8j3YfsRLqbNggsD41vjW+B7jZ2FNRG5DCy/3oN3X4ar
KIUsnsu1DOblM9j4GkfiKqAdFMofpK9pOi2uhTrjgmRzq8k050TYl/ddP9OG2kyRV3hsHyWVN+cR
VsZbs4YC8IoVhKBLSgrakR/9oBKzu1HvQSZB/wRUQRMlsqZJhsRr/1ShFqq5jT3Xyxm8ALl4Nx3b
BbgagMPRFpIuthnMA9OBmSx4SnzfGtufkD+FuEERAf2vMJbup3VQ4r9SmWDsNVFzYvOJk3HyME6W
UOiJ+Bg68qedLEjF22RvORgEfQZaJrMYYAxRvUoagnL4Xs+hHadHhcNMXs6b8WSqqqY9cmZsZZWU
D2RrIPUcV4hXclg86YNCL+rOy8dUO8vIuWrx2SpI8OKoKrhTbYOasQIszmu/e1KVAvwlQ5sOVYEs
kiCDxPNO2zwwKWKJXEDwlUxN2wPoGBztdQR3jhu8sJUiHgdlyPuKo01Vtt5xPEZ18ssOn9Et3aTE
X8lOW7eJmx+Bb3iGASWw7eieImzKcowgZCE+AvU+L5ER7wQ7eU89KgxEV4UHP9tSqayChRGeaqyq
JHEtPorptfbGZoW9Qqsf76dazbnLkM0cke8rHk0j6Jyxoj4wfPOZ5IP2ja96UAAebo53Kj/fXlTV
3YOaALxaio/1amLZL0wx+nDEm8axyenj4i20iFVUgZ9T9T/BuPyz05pfRSwvoA09JyU2vt9LH3TG
Ep13uU9CwHGzq24G8CEWLikiU0IGrNk1QmkWB15JgAxirNvNc7USgY4q+W1rV3TcEbAVPEK9rcS0
95CQLctxAOieqDW9qURngn4eLrnptxrrpA812xOccjI96Y2uZKKQpPLh5fxbiWORDR3hXfqkIoo/
HrZRzkwOf8DiDJXIH6xa+rWLr2miKBGuucwgOs5eSeyX5hrRNkZAF9Wd8XgSKQnBKsw/dEzS/9rE
CGIAzlL3a6U/onf/Gs2lELf45u3vUiANIjOLveNwY32v3DS3K8puFFV1yA0EVXeodb024i9tCeD1
c+S6ya3E7HMmEuUm2Jiuo5pixNRucD2MFrzXogPPcwqvhxwBZyHRrS5VHe+zC9wRnjgsilug6w0X
7Kl2+vgx0yPWg7GFO1AQzClSpC+dIb3jGpaWMPEOHajQiXm5N87lORV43wyHA0mf3XLut5rWFQLX
IUbAm7i1XPxw5vSy3HJjPPrRf0WKd1lpw95NIEJIRAhtrnPWFvzb63F48oyQUIfLavYIXTjveLMP
NO60D9s8OeOI4EXnSkuH7B0zpsQ0sArAvNANDM9UJiT1m7XWDENrItb41UFAMVz3qjqj9II+pLMt
j/kT8uGM+uqDuglS0tQYT8ltW8RfU1LEv3r5xvt+vxRZCy5D6uPfe6y2nZ/+Ys6eP3A+M/sVEEhr
jakYPsncg82gcTZpJ8ugyVH123wxqrQH9g9T1gQtaZCAwWN/Sn+CxnSS2XxzMkfWfQmqLrzAbmNS
Ut14HvkbLjAovPthJZsjmfVDmWhmFjc9SqX/EGsAU7zPVltAEWOdfMHr75u4WcJfNrNHGO+8MTZF
UDo4FFPf3fKbTUjUoNngtZAA1xaqCyuN4TW8aSN57BV9V4wu4IBM0mqpF//a4Bn1yGfTKjGzcmRO
04cplcYZKJmTRfuMsxx3cC93T2yuHk1gUxpJBFwXPJTiwpvi0QL3/qIwhjoL/V3En2Dl3V8UB8J9
2IKDPLrEA/DXYpALxbQAmw8lCfT1pkNwJR87CkSKBmgOQB04SPIMtAosyR2HdSxELNOQxdJN2cfB
Q8FUeQMJxufH9FT29t7gCmBW3ivrvTtp1DI791xQRw7Aly1j1bfbtGw7Ni2crRmg0oRqtnL+QUE+
u1fs1j5Mv6KZ79lOpVkVA9ea5Kt7W/AdO7GyVdH2agne3nxHZ1WZL7I4XYog7rzHjc+xh28sYGv4
cz/o0YdMgZKkiLuPHyHUR+74vLYWNhpM7BOkVh9rwvLLYhtx2W7GiQYMOV33GdnItIAeofpovgKa
bBauEF0kohmUslGIE1Vo5R57bDjIzCG7UvBOpZBe76wqEUW/Y4xz0jzrXax6dNg7haqJJep4kXQY
rttAmEKukgQFx+/mw7EOdmxuVDKsZxK+TjkW9mUqcS90xcb6KSQBLoQmXhOhe9RXT8uWl0ZVgD7d
ASwyMAG4uQsh1kVM1yxzlqJmzvnyGAWT/zl5vKWbS3qua5I0yH9uJX4+XENaxYhdkH8M84jDRtjw
U2mvg9/gt01Z4Fb096WPySIAMZVtN+yTUu+n3TcV98cYoDQaWbC6+jWl88pQHIXVhDjIOvPd38Q5
uQsYCAX03TC3azKz41xnI070M5gTCezK67nMaJqrk4FMuUem2vyww2XQDbvXM5hbUmUzDE2PUdZD
epXgmAWjX0hajJKX4Hocb8cuB3mdo/KOHqBJ7V7N5KEXQ9S848ckRbrhkBhlB25O98YqEOgaObZM
ijLEDEeUEm/NhtoJSBdmEaXbyrOMjPeOg9HGIh10G7kiac63yymv1lIcos/xxlQtyqWRfA2PP3jX
jpwl6Tz9wBjP6zwfVRO25SjA5O1PW+zuTjMAxW+ZB9EkUg+JJujXVVQ83uF0OAZxQFMR8MAWni6g
K+2z6wsZLQ9kgfPw/LeYzQ8Yd0CO6okQHl9odGd0JQgfwI1V4T7bQLgKy3FQZwqfjSV1XNE9P9Eq
jSZz+CKG53levawny2Zj51YE/7Ufx3nuqC0dXHp3fhiAB8izJJTOuAobU5v88VP73euqvgq2r3+R
ITQylC5WZBJokwaSuTN/oAR2mMJw6wvrpzdHFHxhBKRwc+FkU4Sgl4c7s89WO1qatNYq5aTXpXFS
zAFki8q6+dr31xxD3ssPsrgnvNvh99Ort5JTsJ+QF3bdFj2vn9DuMs/GEr5c3HYtRY9d/9YLBSQk
A/lghgpuXmGy62BMPaK/Vw6UWQUPtxwOhjeJzTL6HlINu8QGQWgGbGyGrv0JbRYBwq1+CZUAhMeh
KGtbFnRXDSHCUZUfLzYc4Hus0DLNjwBqsFc5lqIsncBk3+xhc+LHLarnvz039u30s4DJIXYt0T6r
ANplRdg0D9cKAGa7AwmnfPe5LM9JWzkD5/0gyltFsCy2BZfnhzhjP2YtBNQrbU+nCg1YauOU55NX
51RQP/guT0JSQKdxYx1BrAobsSRv99aIEVFgQ77XzZsZl4upoGAVYkd79y+M5baSlX0PG9grw/sX
fKTCL0J8uI8rxTfwYShFjdAd6N921PiVaUuzKo20SNzE/uH274mIz1w+7j34yt6o2mj8gIEVD8dm
eDOe9WSJEaYxozExKc2xFvk/+0BaYuFqLf5vVnADZh4hec7JV9nRveb7ORzCO79KoQOFkSvsD6QG
/lSu8xG5PB3aN+K3mSfWKtuVUPMPKQf4cu3Fxx8CK5R+DAMdvMjM2nzraaQTVueocv95obvbId5K
xq0dhtu/6pkBmYbbN6RrS2hAsp3iuvQkwqLwKHExWCGhQJCm0PDhxtnEu2/a2Fs5rmjgCcMGf/fu
k5a7ugRHDkIdpJyNl5yK1HSrP/nxcQELdq4FnBBvnKZiS6XjPark29Wfq5GrkO4cQnZ0vQTSx6oF
Wpi3IMqENNjO7o/c3L8MKw3mT+9KcQntubHRLfP3C0Ww5XGBVYYrSTlsz1Kcb79TD30nr33PIN4x
pCrT9IWGCFtHU8UXLs5okbjVTmmpcDJmo0NiVZPA6sIC/PpHA/ctbd3p64+1SxfsMVi7stZ+2ylh
BJjqUh8bircGe9ocscdfsUcD9URcPjnFyikMVLVEuDBgK6FDgQZif/zpxYfwSFfce9jFUoE7enSi
xlOmpO82EjLgv7b9C5LByeiUATA+bO7y6D/LoeSeyfX7m9DofvlEVeANQp7M/Hueo/t5f+5Yen4G
773asC5jmX7aE9qgUrdm8z2UhnM2TaIqTQ012AEyeg3whc1ywfTooy2cL21QxcpvUxpe7dWCe3qT
2jd9xRa0uzQt+IVIlWngkgAkd9VeKbiSttGhBMBs5cy1ur6aHfVW2JU2ZEJiZIgXLQe0UeAIYRNI
lkgT3y/QxAP1CyiJWfckiXCF7gXFCkvb8ibffqgkoU5awe9MOKVFui8UuvYC/nMRsrcQ8X19C4PV
Cgl5S8gfIvid1OdzigeEW/bf1WDMMw9Tzefo9a73iwWPXgwEFfPRgBQzXRnjOc3zaai5ejIrGz33
HVPBJTBPXNuon2hLj8sImKVtSIa5J1VU/OeWmZWwYkdb/tgToA9RZpuczA2wcqgOizTsWqbcM0Mm
5UKqSRxr4Brlyz8IbnwLHxRQhk4mKdd3kimxPe91OXmTpAEteW0GKGXtN3gkfXVKzpnkpScisFPv
4KaVdPLdQvxOsFTSMKcMrewZvs423xamUc50RF0+JUMPKqwAj+BJQkcy7V4IaVX7wtCjYmJdDm58
ijlPQrRSqqGM93Gg0dYe6kTqSHWdsHPzmip1pW2DVs4PEvK+jbgC+QOB/rLLJSeIIFHwpg8ebhcI
j3voegnxOsNcpwbkYFF1FrSJhPFyORu/DenOlQyifbWQFwk509PpQm/SMZn2T5pwU1xw8yu6H6gG
7QUsMcquhO86dxf4p6zvXPcy4es4aiLIW/ToY4W7/ckKjy0384hCJFRAEwwtZjppns6haswmJTCP
/MQp3QZcZm3+8uN17bTdzjvk702Abkr53pui+r0XEeBZzb3nuC3n979MF95kEPpnqSAWCcaVz2zn
Yzxq3ycStZ1FJMdd8tiYXON3jREwEgzBUIaH4T67khsN9AqZC0JmiK214+f2aFy0UZiH/tm5D/eF
vxaBZOEMPDszMyUiNCXpMtgV6/WGdg6ph+mY+FV96WTdEmqUuOUtWldN9xXF5d9URODH1GQL5Dp2
TIi74V62agdAEd5Kd5EQeZ7ns/fCrTVZXm6uRBKlh8AqluirH+ZTg6rb4KLz24Y9t5Z7QJN3af6t
5rxuu0J8nr0j5DMXWCKlknx4k2oAZXbYzOd9w0iSJkcmILw79mIfBfgNWWK83bWh/JuYMHNiLQ1J
C60VvYs3ePkRzH2JZ83SxohAW6n6C1tJLXXjDXKBppXP6gYvgOghFhq+GVKzfkzoay8+aTWO/WIN
/K3SLsXpht0kV2NiJGFLtbfc7IxsuujW1JwhTOGFESencwwBoK9dySS7GCsgxTq0TU05eidMJJ2z
xEaJxoa1g5pJ7ebTW0taKDhPW23Zmx0vip5OCk0PxdbcIbpWVf+/c9W+RYPYu4guSVNzP5AK/2bv
inPv4oyR5qp7pyzqrMxYmBpS7o6CTAmaigs25yik6eqQBbAPBSxFmPd3LNMItARq1M8PkaYHPaWJ
IpLoTSSZ6Kh/Ucln995PdP2t6RWNgiCfUm0Z1xhIfVBpEz98AEbbjarpITBhLPqucCAR32yqE/Bb
HvhSl1CYyYVScpsiXpywNt5RA3tKYEj6pOX3AYV0cHy2jULWYfqBrZS7XY37fpdtvodRY4BoQqR0
Zq/9WsRrpTvX5eid60qqNjLlDOWPOj5faV/Mc3Dz74k+dYl7YL7MT4blSAHGdsT4g8fKxjpxYZ1w
rnVxqItZoWU/QD0sV3sS92WIGpa5epMaUmfWSuisVDtk8SPaDt1HcyJ2K2gOtvY911QOzxnVtXEV
ZukGbKLnJFfbQ97sb4Ajw6KAPqC44fU3HxKX34n3aHt6Tzj1fgSWvLyE70wWcNlcvOr3eJZRn0ep
eHdzVq5B7xrKD8gXfBfJDay2VNyImWh6vKYHm7/3vF9TvFIvrUKWO5DTua6UwOryp89JH59lxMS3
D0CAIQgCM9E5DcEbzP3wMHtcLEM2TEqNKyjUx5pLHBaOOJWmU+MiO9xDmoIPvVAWTOa62OqcAvJq
dhXjCbfhgcYsqDbEdw7RlfZaqbBfSH3JRdX5HsdKgCTKpbBX5JzJWsfALXIFS1zH9IW6yoPAxw8v
dkq80NhEZr2W2dWAC0lmzM1UzqcZZSokxMnrCwdKGmtpO+w2IiM5ISVeBNNXqst9UnO9N0gxSL8+
oxdkvylMnuUfC8qUEW/ClNz6fXos7pq7EkruC60PL9fdc4isKSg837H/KvcX2i7ae9Z1uRIgnhLp
rHQYW0Ore/c6nnXbnpuEEywXFon9CmJ6JFVFBjL0ThRgzMMYCpmWYqpH78e7nxRnkXMzwYJ7au4z
PvBjDZNYEfTHa9SnBc8QmyEqoHZUHQ1cNPAeeUVuftMT/qUWsPk6O2Ot1qsWDuucYUvHPjCdlwv9
BJJu+fra7CpGqmpetw/bk9EgKXDuiOBA8+egmbMOOM3XLIEmfTNmr8cVL7gUEbTUYxZjTmYpi/Km
bwz60GzvaGj1lb+04DFhbwkS2EI2b3YKcNWSzKt0hI3oLs1TpAmkosXBEh9Gsr/2kRCN/sHHUNdJ
YCGBQNlDoelSxsWGONDBBHJWikdyvuw+Oz6D9YMeIbOBEWn90CPqVEyCMk9/ceMzRpvgR5wEfC0u
nmdI7p/1fjYBTxfGlGleuaw38waMeZRkB3Nq7gOrhLwBU7exkUg/LlO8z1SuElPgk+AeLNOFdz/6
Ry9TjHg8fwP22qiBRBASlC9Bfb44vWXHflhxsBTFWcqJ9F0XMTB8N0tpCwlNIrnGXhKEsTTzMsmz
2f8ObCZ2zS0egnR5ABzmoiVX2pbsjOAhla8pVp58xm8A1COqSLWn4tLsjgT45a+BfXk9rfGOr0jl
zzTcBqOTlSP+BvVG6f92lU1+osGLZtYq5mGo8bdYNRPm1egs9cFX1JlV97b5yX4OX9BUfS4260JC
K8nfqr7kKQFF9uzYLBh7jYxerYrjZW2T3999VVpd4h0gMnI1SqHR9W/C07Ae6MQluvOrX+wvtxTP
Z1Ss7al0741GWx/RLg+jHnPY6YwdJCvrSCox0vER4S6hdCX8MEQLGETpT+tKwvz3bUxIl4VJak1Y
XpVJi7/rIianuWzvzT10Hpo5i12tvwz37e5pMdohNu71m9EHDOQGPkq0WWDH8l+UaTgxWGgNjcBY
vS1PDILPzsSrKvJ9wvcMGVFlK40VvgqaIBwXY8v8BrOWYqKKcc/H/Nybb26WvzQbb++AQlg7/7c8
pwba5auI5XolPj9u/iMi6bHXx61ydexH7jgFzN1fbvtiea46XPuUak9cfJ3TwqCHhgSeH3K4aNwV
2jiIbTM3jCjMAm23Vnhpyk3T3rsc5lS0CfXn32rQd7VSIwdlWIs4ZdaDundahP3dPJRHqCRuA2Ae
aiN/2YfoFpiPaDy/WGo1P2uozTr95/RW7qmKb/AZZYOIUi2GGASQ3ts5zK5RDa3RCo2StA8AfJJh
RSQ8erTQt8hVkqJ5Qf9jJYXf9k2rmv54qmXK+Htj7kgVubNcmWXicZ74ySUWOiR6iFMoXHpqwXKm
zc3IjvIeubd1dIWnZZyslM/tGsw1Ouvpm94oZtLkLK2IpVk2UUhihFFI39gnV8tiIJ7A6pL/gvq0
DpQ17h0mkKkCt87AWNg0BvWzIVkqIjhSQYHMhJuvipXNDZPn1VcO3HNuQDri7T/8vYTfJKwaziF2
hpzRv3AtBDnZ2pZ82XlyBYbOqGpz9QsfFD9mTe0gIAyotsbIWXedcIFei37FZ+fs9y4Dt1jf4wZt
Pdu3lt3fvuvEdSHkuE1e5EqdtLWouU6LLxZZXSElmI6UIaoERJu8VhI8d91Pz+VSiUmE0Wj4LQfi
imA8HAh3bYv1FSF3yfKOCWcV1rcSKkmvELl6Di6ElSxoxfQcidNCmcHzMG0WJW8hoKmBofvJlbH+
oN0rU7lkOicr/sX4r9MPR1SeVLbP2uYM6GmDB4bdM1XKy6Gfa22WIBObLFLmYCnMt2QeqIRHL1hz
9LKD7Rio8RIPZfcYZmszmPEcYDIS/LYaH2KPlDP35T8NIfWnfJl2+6dTOuuTDmTnx6mBUHXYkCyt
3s4/inuePE1ClFeK1u061IBPqeOZ8jfePmkz/ARND6SMl4XaFZWyZNjOrVNBGz1+mRFkOHKkC/TQ
X9v/PkrqPk5CcSf7rHH8XKKFHu2ionKGGunEjjL8imEnP+UkfwxHdp2V4FxTyXhlLyHLt/+6AjVj
MsFJYn3DaYsrEZMUcpvPd8LreEiwc6gaWv699hj2VW7vna04QKAavp77oavORfJDe6jeDoI3aFDY
CJz/UdrYmRVS98yuewZ5FD3QjT2gFiqlTr2wzc7JU8aYacFV34RuGLpeQtEpFqu0uLzTHB419W6+
kKY9prAdw6Bd19hzg1dy6vFPQCO479QW5KyrpYE7nAsDh3cltzc9bGpw/Il/aXSgIxPYZU3VJE/J
5LoGwrMIvhLZTgR9Spns8Zj8zJyjZburQzkpR/rsK1QJ2laTi7ey/yMGcXGHWbcUsnz5jfwaHNX2
+L4Qd9/ydlih5z79zeRKP81x5WYwq75rIVLJ/7JaJrI8JV3RuCQ1CmsbF3EaXdvbh7oBHeaX7nAN
hxJGA3pHi5Wqw+06Y+CB7VY0kvdiUbBtNZ5nTMb1t5JPXW5sUmSWScBKFwe5LP+4Zz8fWuz4U0jC
EtxDj2q/aA2/5+5gkNolbHB1eJRfhUyyXrVQwV7EyB6YXaseq0UQBiC8L87uJIyV5rnIkBHobnpa
+I8j/BV90FWJqX78oM9arR8undMdo42awPY3rPCisgK4B6JgiHTD5dWm6SYRY9GfUJoeDGiROA9R
gHJtDj7/CDAKo8fAvSwm29bH8DxjwbRTKVUDb8GCQB095UG0K6TKFO1wKQnCDeDdQvoKsxQfHwHk
THMnemmdsAo/aLAK5Wm+7UXTuyonOVZjNdHqaO5z1H/t24bpNdo51ycmoj5Nig1tsaT+/235VvwW
e+b9F9XgHXApU23Q7+qADMAZ3woHeo8KAz+qEiFSozPhgJ30Pneu0YCR26BWprFTiutnOi8r4lng
flVylR8V+hDCz39ACXbPT7mZ6hMpqh2MkH3OFybZLYyR7qeqhQ26b3fPQ7Z1WdRdk5HiGJSv1AG1
xi1bhj2qsmPnVbHESBEwGazVR7d6PkyZKn8TimIpMi9C6y+mC3rQ8t6zRnYW67Uv/sD/5roRAv4k
AgNJrsDgwHjlxU5CI5yoFrlb7iV7mtQgWymu3qjlXF8SwOmKiyJq+x31iSIRPJPqRmYfW2Bn3Zmi
kuCYRp6gSeeUxoKDFlVIOqaIt4nYQjLf2M0rdcu9frbcy/ID/QLRGTH/YY7oM0CGqw34x7MSUi46
i7R1gi5/HVQWdIVBR0hAoEmuDsOhRhNXQAgt3nr6l4XqWrLyifCS+8w1K21kt1sMzPsEDIITRagj
CFmXP1RlRbNvyWjrBM++oMd0h7j1I9Hv26+NaPQ8TNAL0uCMC/tXwxJJPSdrOBphszXV7CLPELG6
taYnUFglNHkrX7ukNMcqAfExcFIwXxndY/Czg+zbRJeE+2x1VC/XoaeafyMm815TwuVa7B7csq3k
QVCA9aZSclInCzBwaoFHyDpjxuZxwPwucZ16+di+a3IIdncZA9CILDGQXMIdPEZZd2DlobFT0s3X
cEdW8j3sCX4xNwaNj+998A+6X3ZJktc2cpmbdPcJ+fO+IMFg3IgNzXiSTcvW81GhMZxNsyhzmRvH
mlV2O/DAlunsvdX2dv0NTtEmYiLUhWbsPLhV3h0DS42jCGYmjujaoF0BgC4lLV1XUQNQtt1LL6Q6
VlK4/7wjKlEPmr0BARGdXXs0Mmjk8fBdqmkq1DsIlHNWmZBITnQKO5Q62fF031GVkkij5BsiHh9i
kCoV5jsWMPpM7v4H9LaLhqUVvTvw2R7KNebFcMj9AD0SHxxmbN/Q2Xz5DuL0xAi87FlU15aRQ+XE
RJ6q+jRw9kQg7rgdwKgHQf0as3n7oXNKlnJcZ88rAay/esDCNkIHxZpCBlEoSCu+e1ZuXguNusQU
vQhSPnhdV5uASkL+JFJ1z3rwPLVJwfMLyyVQtkYLbakwTxJauW7onLVRc0/9tngj2wQ+lWFe90zJ
zZZ4ujobUh9CV1BxaeRC/xjTtECitEvs1HQK+zFo0gT1xY6iA6ijYsSq2YPI50Z8+CT4944PX6BU
4KzWLNGZHZXk3NhJB2PesaOYdOEoGfgnRTlWY30oYiHrYFDtCu12Z/m1wwPOSaTgOEzUlPJu+ED+
IVsvDfLM7/btV4348FoTlphFbkrP++NK8gEuQqNhcS/lcdjDdr3/m2wczQGl7SI2F51rSTsIss4v
2PAmF85DASjhhO5r/amuARaFHDuy92C50fo1zXD8VxMhB0DepORQKjKO84LQGtb4IIssm/9u91IO
zzFfOA4QF0k1l4Xi/JJ4Us4c4cHqUaQ7JV3rXMLUnFL6mjWxTR55xdkkjkiOcNwxvXMf8J8IVc6d
ftt0SXUlBp+nYytKn6q0S/LqPSMc8CoPD0UEsnFanf9dpUQlvMRp3fFmFRYCn0KGsDF40Z7TXNga
23b6CR0pCJfqSNfwKvxzHJ88EXJSdHn3ISq9QvxBGuiaqWjhMWuyDHKicIj14p7nRhQw4GQ05k4I
Bg0AXNFwj0uwr9tB8VCH2MmRuhj3ddcgHemFK91wSM3qdDJ7+WlvdwxjXvyCYLlkl4N1Zon2zfWm
FiYW8/ci/3CVe596Cj0bdBnsM7RWh40AFyrS6X1zk/qB7O3Ou4ixKvmpUczlZcVODShBGn7Qkqob
MPKM0/CzdPmm1L9knrtr+3kRJsgLehz47v60xp432TFXSBUcDoWxezkMeANz6ZO4Ma12eGPYSDFz
skH6xLa0eNnRuQSYp9tqtz1BsCnOVdvyAICuJrJrsTQiYt2ut429mlwhv3jvclWjs+eKL6Y40mfm
zIuR31vKeoFPaLszfTl42Dqyj70W8QabQkpZ0FENViKlm1AsSQ5IRknIT+VxlkRnxZf5S9tHmubk
SnFLkefWdvsgTQVIvrLcMQP7bC1NtQkDQlsvnAZQwwrixC4Xme9Ent3Xcgdr6uC7wDIbWDTyAJ4w
moMbwhfuk8yt85UeZq7KJ1V8xtFth8arXKqjM/qrZOM6KkDzUWypA70qsWk954n8bzg3hDctx4At
WIgDD1oVKY4eAg+Z0/sWVgvYbfdPMKYD3aqvRxBd6zX8LtVhHaS8L2wghe+aGZBqPu3JBWFkD7Ne
rDvLMyNHzjTeHMtU6EfToHrR7QFar4LTZGQUo9ssLxBK/vNM3MZIYp8gyOLfO0pj31C5ewQIHp+H
+aNYmDvb6ulxg9v6OmKHFHdcqbrxFrIMwkRSwsU3UpGLRyMVLBm5/x+epOH2uMEf3AbTeyL8idHg
UiwKxueDsarSTf3NFJCKg3/2KZNgQpi9C5f+NL5bksmqPSQBuYS5bVjQk7Pn7eAQ7y3ST0wgKDNm
fDaZJi07FEgGs0AvVmaW+YW6zzeXehJnAsM124aHQiy3ecEnXvkMFwLQHa9xdyMv54OGvxFgvDWm
yBhoslW/5Amutj70AcVd/ltu0hNraNKsTTC6JH2q93LSKMjER0oPOO620k6yu2vVA4rKrJ5EN6a+
u5gI/giEmViwOgNEXgYpxbbyo/LrEksBn5Zqfb2HzacSrjqFWluY8H85xfm5DKIOnafsxp903iz5
pOkJzstYtSB6acIaC4e8vZ+H5f+8YreiEA8eXLbn7Od/Sj74266JhMFB6INoWy78a79q7ChE+v29
OVcBy0eufrIjY+IRZYM7ElsK0HpVHtP7Xt0s0uzbTG4pM4qZ+023pDFRGO/W8rgmU6pTzpCsQrW8
UuGEfqdtaCPO6l7BVF19PvkQ20hfTBGK2921ZYpfRQNpHsw2+fJJ+884ZwDWdqbIEb5vpooKITG1
iK4BXpYjhw7AixLuMQl9iQc22Wil6IRj33IbzGywVJtzPmKuUDQvdFtg3xCHhgNzXx5jTTuR0EXh
g7SP6EwMjx0BXVQSwDBmv1VYjSn/Qmb1cdGvgpG/wKSdrDQaqDecd90b91esxRMQD6LVdtRcMLaV
HoCxXCZxfKT5i8jPnFX0xqjLLfPkBC33quqh9/ct+/bYYNx3mEfBpFBmrFLbM1OQb1XADBuXdsIJ
yOc+uzl/Pb996Le+D719E2ZkBp6GuwZOIjf+l51h3wjfuWYwyZE7mTtYQLI+7bVQMjNW9rdqSGdk
ncXsvRWkTib5IQHWHccosUFWOrOGDONZFUOSRa5VjEyllk4n+AG8Nwg/cw5hWcRGYKPW3pv2Xo9S
EXHnBwqpjIPn21OiutNvskqlMP/tHmvcabZZ22oCJ/fcEyYsvgigSdsyTompzxHQVWbl1c/I/S1w
YkGsPOWsUgoHE/i8cj/mhWFRcJsPssjO9DEo2AVWAkcIq2uSOqgJ+2vQ6AKkZDyPT5w/TYEywdR/
lqmjs9UOgV+C8U6EodYUdZm3crUHVf7GX6ruRwZOjfKK68XYgYqcc8tJR/OGjUgdHs+q/NbPuFk7
oR/TlVFMSm9Ex1qW+Sw15DXY8W4K719zRh/dVgbUvql5qBbjlEdzYvd3O3N/A9r10IKFpJxdesaF
YyuAcuhdzTW5MI9t3JNTc/u+SYRD/PlSKDsGXO7zQmiTV4kC4NSIRGWoKW+FGhKqwnf0aE8gZuYY
wxFPQ6LGqE109+Ax/rnv6dCqoXXb1puW7WAV1bhacNe8qU2eOsweQ2NS3bQCDZjMflhZknjhbKNF
OuxVKMJ7L/vuCI/eyYPcB4zF9CvRTxJJweDt9PV2/J5hbX+dV3IBrQZsSVvAFZg0BINzM4xOUJ29
drCjK2tIXzebFmeY726V5qhKxICjaEtXizC7hyoPcjvaM6ePXd3UqhamJZZcd0yo84cjGfBTpsmM
aPx6LXpkeMmQz4lFu90ylmYhqTlW0AgWJtm3Lcg3X/p74YiePd/JucI3hLjcxrtWC9SFVsobRnvc
qMEOsblHgnQAxSBksMBEyRU1TCd9spKimWsracAWZM9xB+uosnjbvSCXW3dKmB6FY18epS6FRlYn
RPTsxhb/ycVqxM+RWeefgXcxkITnMld7cwXxzCviaTJqsV73zIQ5btJYwtkEyU1DOzu2sfWtR1or
NIOKNrPeJ4NvSeTRUt2eH7mKpfPAZ1qZe/nlOgyZ6wN9W3hkypREzWhvwLJK3IspNsGKGPcHIYUX
Q4D+qzJ4kH3RTuaEd7VLos63YKzhjpcX6T6rDtFL9wsXrea0MHg2bJ2FQjv0z+0o1FXtsJB+s8Ba
9V/1rVyuEfecGk9E/30TEpsBNXS3aF9fG88ZzCu+iL8dF/UpSeHA7DGL+0stqWd7PA4XttCWMjQS
zT4YJq7TiNnwsb7C/onuC1Rf6qERTK4la4SysIkmRK9lXvAPQZgvH+DkmQd79Ep92EGnYfKrX0vJ
fheYaHnBdYZks2WleLTy3/GP++J/kYt3/cjWnjd1yklmeMB6Iv4Hy4sBxiyMDy+To1wbK+Bra5Ai
B6vQKnoLukmCiGbqeHiBF7CUvyEGKpe6H1ACkj+55XFNaKHt0Ggc4fAdJ6KUkkcu8FvEdtFuRQcm
Qe0j6xzaA5MDebyFxvGduGJwny5Mrnc9+shmOScv+RK0DuEzq1piFCBwXS8T9a1iGYzCEjM8XSW5
FN/SmJH7c4fOgHD4I7Tsyp+Dd8C7/PdOTU4jnM29rLUkZtVxeCiMHCDoM/jW1NTyjo0kVo3jNent
aKDh/LllFXFOBYCa2Hf1wlUAVmsHJOfXiQgTX9B5kisPB+Zkfpi9j3c9MandI7Lp9YtOXjqv3FwD
/qfYXoiKFDVkFreD6rrTrlLSq0qlbGe2GwCT+chDA8LFvf3wfCHA3n9FGdCObJwopKSznj8FSRRQ
ogt4lvcqyarb0Hb7Oanf7d1Nnrwu6hRTP/mUPsT8C1FI1QtfJ2/YKEc5UTHtDsygitNVloScotcT
/mlpRbu6mHJj7sJK3cPTW2hsfZhgkIR1WZ1hk+9HBrUxOjfhp965+EbIyeqrL6/S4K2cEjZiTI/4
6hJKhkG3YOKtIOtf9GHE6h8Xy3q8OcDnQM40JHmiDsDXAIq3Usv2YilTw1IeX0dUSqfDKD27bxs5
a2RDsTvbKDINozHfjvjLRAc6Mu46sYZMi339OYFV/V9TV09JFzuiuEppEVVJw0w9fl+FC9mCKynW
TxeFO48tYoL+Quv16hDGeTfZ5gT3uDOiD6wUfj4NLBZfxUJ9+4CO2m4oKHeVtkCFqnZbjzTXAdkx
ImBMkB6s6J/JpFJUbhgcyHFaz5adiI8Qxb8sfff5oJ1zQJnomXItUYePo60YKpo3aEVomvJVJUyE
jZ2481XCBAa9qckEo9jLGlDulqt8UuGHooHFSCB0oJDFmJ3J4++2gfLhHIe30U7Cjv8sTnnFCxA+
v1jrvKswxR+GI95j+bljYtGj8KFkn+2dfp1XeayqtNWIxGfiVNvu0amLFq2i4kFtY08IuDSwrN8r
Q1gfLS+OocQ3APrkwgvN6AwaGGlvXzgZK5RgRBkHOu/acJwtjeZsfxRAz2TWcD9982y+DE5eBm0K
xWUeoC9IJzxSsYZ+fiM3s9Lce5h4pDI9EWV9H6Ve4Kf9eb7oe9ZTyQSYTtYmETZFA9RM9VRbUmIB
SeHMt5UQftYXLOVr637HINT14mDzCPQ6tlhPh6JRdwmc3MmTpfdLZC1RKd5Bq07zJQmRgVWND7li
wNe8yPRpTAPwe7N2Ae3P2xfiKHkO+TgqNmAN0TxIm9FpzRFUZdKlGSiNk/UT+okUxdK1LEjFuMeL
WMpUCJx81bKLqxIsZqc7PR33bf9WpS0ljuikzzpsVmmGIgAeWqZoBUo90fX5H0Xh30kTVvT0Z06q
jciF+nryDNaVqrJhuF7MCPYyaXYK0hxmlmlACrOvzXBIDOvO8APc7tbSqhPeu0b5k93/Q4Jn/jGF
P5bNGs8lrwXQiYe9Rqv9GmV4IXdwO7C9c2oE0isooXrJO5nWiz/PYVPH+frlsQu2vF8gQ0ADuRps
UVbr+T6qGCp6XnVfRsXCkTWqWryiJxR8NrbQqucNb0x3HAtlTaqy9zreVu6VQHo3ylewRr80H8+h
ehYHfq7u0eHI8vw0GUVYnUhavlpHA9mTMZGv9LJAEWkcf7uVMKN8is7uTrx8nyPa6h8Wzs0ZAO2s
W96gB5+zy7+uCO5jcxF6m+NnrZu4pi9pImpUUdLp5/BzB3PVpeR09yK/28sOw+MWJfRHdXBN4N2U
oVrFfqswSZdOR6EOlsEF306pLE4iei94yfEx8lYphDaYRD6gOmxTF+VgIXvRTBVN3cmACw7oiZtV
GnV3ar5lp1FuW1XEoPqOpPgLrGm89IBIPPdjqkjo3vtlwdkaF+LZjpLdkIBM2lLS14jrNqvuwYR+
N9VKb+/8VIKS7/pLYYH8G03uaBcp+VLsUNNt3t+lMfVylidO25OY5szEh3CIyZvpMtDszGn5BEHD
NkYrtFitDfDqmLL8hyO0oHnLOftZuwodM2VF9ukxDjLwqnzhvXRNJNvliz204VxAONnuUGQJRzJ9
4TcfKy8BxxiZc7nkBmk3RmCgudP4AuZO19RDSNodLKKw/aee1kE0QE21orBceHxrA+2Qy/M6OVOu
kAo9/i4przUcv2rZCGDHwnUEb839sHCxFZ/rsjixxrYCvt9qOV64dLx9uqinBicjOMzG4kehV+5m
sDQ3y/Az21dimY6HJqq00HurXM8V2FkSrb+lkGgi9KH7pm6Xp/eVFX0nmOYARHM9vOaiAoH0lQQ7
W4EVybfakK01Gl2bqE8SpfSRa13FAy5l9eUAQytQyT+wWbHxkDuldalLETd2NTiRkVk5OWGn17Ix
9n2VZkJzjMerAyag7c+7NLVmrDH7OnKXtKcAkSXpCJFf4MDNJbz0esa9F+lCS0tgrq0h8bsRrK3A
57JsIHEK9rKk5ZSZ3t2U/UyzGdFvnag4T1U0A4p9dazu5hVnaAwB7CTtuO9Z54OC0qIjbyAdyqse
sjBFZn6d6gXFvonvCSL5kJb+ntx57du9XYZsfiHYynALWkEEeonJhe7l1GZOlSwfZwaF/L2GwGE7
IDxn+ork6sJOvMU76pef0pWe5RT4P7hGUk0iOjHPaEo6GqxBwwz8Q1TgCR/0b+Qnqsvpws16UBlw
/JcAJP1E3y9u9ysa0TXBMrLrJ7hJE6Y5742Fk83tBsMnIwPBlDY7vefkOXQXK/VrWO5fa8yO7Xyb
m0+HTDx/Rzwar/PU+/fMgBBVkUO3dw3JNYoE0ZcLAZgQJSZ+dVxn+SlXKqw70sYjbLzEejsl7FT7
uPk2gSYu7hUQBiOC5hBCu0Cu8yqKIs4EAFHzfGPeAuUxx2dfI2kqHvo2LRDQ0bHIpvPLVuzM52KN
hpRwPkQSg+S/vtjKQY657u3Z9J0yeKkcIStvJaVhPF+guViAoj/8CgtSversKunmbdO5NyiaMFWd
bYgNsQsDg8wV4mBcJtNdPqzvnzy4e7ZKlHgRvgBDMsS13st90Jx0GKm9D1gyonWtbZ6YA1Ptzx7x
Q64QN7J+VEWXeTs8CMXoBg4GX8y2xT9hEHH9SItSZvfCEqP0CfFD6O4aH/Xt5JkIHZFYBIiEYMek
gDIKPdfABWd/qX6pAlCB1Xkp4Q95PhPOQEoe9WqBhlb3F92EHKMq2uIbmfSXmbpDs9VCpFyuisjd
e+y7BCQPEkb9nZtdroR1iRHtfiImWL8XwK/2GBlq7FOzzT00oRiG4HLJCqIt7O5j4zViXXTofiO1
xwXgt5m5au7Vt5O/b8BsGhf0oHkV5Od6KLfJvhsfAvR2rOmxLd8Y/igSXrkL8sfRddEMs3iJ3Cgr
I0t04DXXOXgHxlRvUwUpu+4I3TFOJJ5b2/xN0j3lTMAeOUBi6IFhcd8plpXKbzx7CEdKg7TCt7jQ
mQELYRWMhiK6GE8RbGy6AVLIdygH11LWqMoEyjvpMG+muoNPgDABEw6MGy+3fzzzky8BtAhc2fTI
/q0cfviEebhVTyMeROz4f/WaTxTsgaJYXefPLTNxhrjweyRZIPa6tF6YlxSnRQMFnucshbLE2TOX
6ajGI60LBsYTIAfqaia7iL0WayYS+yGCZ83SYLa01ul1E0hvwcto+8p4q2emoygv5Vg23vWidyL+
q4GIjXE8pkBouXhrtkHzcFGOoFAD9Vo3/p/8R5eD5kimIYlqKKDcxcwcI7qr6koC65455RudkuhQ
iVv6DERM9A+bIWVtQofq4hwfGAI7jbqdqrdeoF+s2+MHV2wsg1eI1EaQCHzub9GZtbIWv3a5pULy
DklS2kdkY+WzqgT0NoFvWz/JbCEiwvylxHbdD4zyUrPIrob8IvSkwpfz2CZLjkK75z+RVY3AMKpP
peQLH52wEChLGH2qgimP0XASQjYZdLUKj6VWJOE9DeRD9n4swvPuFvXnTzJ41bvHsyafCCDSqDen
uTPSj+sr2sG+XcLwNMqfmPMxqE3qUu2FmlFc4cK4rTN3/loj4RQcw0d7lwwMWPj8N8KJlRqnSuIl
rg0AU/yxdNsYQi4CS67wpiUwlTBpXroubGjqu+tTG33b071SRxSW6AiYIWFwbi94WcynwtLyhkZS
Ds/fPfnIK5ez9+nzkCD+U0mIGZGqTYeIvKVG6PmxO48HFnYmaNjnEyyCVD8yYatxDi9Sp2QOMvdM
MuTfTgFu3VbZY0IAA24NFDLfDSY6xaTRdgk3AYFI6hoIb4W0Bya4ZqgRPIv66MxdeCcizPunWQYs
1SDD840kMFOFfZ3v6KWHXcyDKbwUcNnfQr/Cdrm7Lx/hiLab0i2l4D1k9o/5O8lLSB3qv1YxMgOI
8UyStSBlzP9WiOUhX4jmdhJPLy+yqZBTWWJY1Ty6Qn7f60M22UhRHWTEwT9Kb2XTLlZZNa05Stts
rPhEvtsG+MxC7EO44lsKZiEKUv/FYtiuB3JaMkhUX6E9RAfGfOLEoeQlDBymgx78il4g+Tw01TlD
SCwSYgFzmiQrqFuXzyhlfSRLI5gUI5l4cPTpKx2vbOJ378FxaAzUg0gY8zhi4qXw4+Dc9i7cQ+7/
on0IJBd3tDmDLlNa11JDm/tSZf9ANdMWKzmlNCRe9zp40/upOaeWVr9nyebTBjLWAmRj+uhxS72T
HvHNTCdgfVnfGZStSdnhZca41xt3cjg+BtIJTRxtFvG8rMWU0x4oJ/23EEZJmHSRFKfja2jlgzQB
47WaabzkrsQirUzMkNnASl8DGuH5+EDFJeTiEQVp1mxqNrMk+zR7uRIFmFIP/rySLEjYOvM49EBR
qb60TAlPnu5c+FnWUUrBtLjbb+AW64UmhxHrxiSqlWSKbBK+iWAC9ByWz6ODqqFTrJCMsXd/URsY
mUGmhkhMAfi9PQsGefOAb10aFzxhbWWR1kMfuwODbeQ0TLDxz490Ub6FUWd3wo1181vEKzx3qtM5
Fn9CqzRvDIOS2cKoUABnpxbQVtYh+RLJ5s96MdLQhukm/17lHBf/d6iE0jYOCfX2nZHwjSw28dV0
GAri/V0AvLCEKw2mZwWpOWC6PFrZN0Jr5xe89Ka4H2pZk82sijEGsZtVrlrVDZewaCiW2c6d895a
n+PZxKsndM8p1SjVvdWz9gnYQ76pZ1iEJuUKn1lIexv6vkHRBSOuxWAoDgE6rV6yXnsobyEkHv7i
62GbGdgyosmZBRC25svuKg+XcBjW/VgjKe9UXWZeDP+xUY039HlmGrItxNZ5hNORoDmvCbiZOkZB
3qFwBuz7fI5v4IeL54KzvOJRQ8+07SPgqz1ccHyrBcM0qy0C2nnYni8x/0AL/07uNdor6aJ9njoi
Fc1fYVN+b97t0dZXreYNjocv9wOIvwQx7qfxVvMyOeZqfTGulpnlP1agn3MQuRWN4rQAy4gayiDf
XLDQpJLeB/BURTU+PBknxP22Pg3bcm+iYCVeVA5OVxxqD/4XwOSiHraA3xE1yGXn7TiSlbI7hySF
SCM0TH8Bjf/DViFMu4SypM7cFGQfLfr0HdE5ygNQTeA114xejatKTVsrnv0sKRuLK2fOVSNEDMIY
2cfV8TdINSOHouGh/3hjl36XGuaBqy/BE6Aw0FMzZCfOnxlXxFww6j8f0qTWEDIkM7VTDH4VXPiK
nhNrNe9K+t6kKnoBKu/fzr3aHAXAA1H6srQp7EG3+f6Dw+uppkLsdAk4IYQuKc3ncufRY8X1Fhjo
sVwX/PBr1GreaDExCNuCx6V92ep45GxhklF0ypjszytopukWvAvp70chErJE7c+JLfwXV2I2Oem9
dQwpKgpFprTiDS97z428UnmrmhDy4ztK90EPR2eWAP3ZDOKzhNOfYXKe0kAJC6TZcY+14Go4ryvN
IMgV6j2gNdpIcr1/s3PMSlSvCUscvSR/QUNTUUkAuMy7Mu7btxAGAnknZTrXoEdBmr2zbrknImY5
Q9s2QccFZKIaK/x7HtG/8DMApIPb2GxEFSjeBjSOp5VmDQzf02ulj1SfiTvc1UCYDw0f3Gv4EkAx
1Q5Vl6RJuJZxmnZZkbdHyVijmYQYOAqkU4RXOEM5eVYT23I49Ufi9Apkrip93uEtX32/uDkhACk4
jIn8YO/Oxp46Z7PMBH6q1UUm9b+DI8TteQ6Dha3ZkBDIeEeeVZT52k5g1atVuMOSUUKj1qatQWQg
45K0UFSz/Ga7aSyeM4M4Fs88qDJ/+5WhtUn4FoVB+bNT4NhOEqwQzXyDm+Hll8VSJxrqwLLdwXG0
tdctw0T5rBQw7vqEnSr1yggJFPMQT4hIV/hsEX8xmusFziRItp0v/uTEpG83wHyJgVSUu6ZalhdQ
EbZ6q5muMxrNZUrZVAwxyl4zYB+Lbof27FJd4LjLQwiQNikd5gkaoT+JPjBeV6TSk4vMtFDoeMCb
D1+VhvdBPgFn4mxKyNOLExEyvVKFqzdnvG/gIMOAvW4urtYRnzktOj3ZdVmBMAfCIHPQHE5gnxPk
WJc87xedaACm+mboqDMHXd6VW6+/tqGf0K2jvDNUkqaliUFnUJHEM/YWzykZGYutcslUwUAL+lv2
hU7IiTE5us6pdhS8Hy+fHhQhPWR23pdepmBjoXxunSNlVBQJQjoimz3/OUHEMa0WKFCr4EJClI8L
n4WeRbyK7UO5MLc1cV9fKjJD8liPNgHnAZXeao0c7uqjLRq2NTcI9YeF5OiqX2ZJlNzLJD+c2m3A
gua2jsu2w5fvOveftT23U9U3R+8dQ9Y3K9Oov7qA4D/E7z8RnBY4xGcGPkq0mVQ9xvBOC4vFm8Wq
VeF8V0E3IYegwM+5A3uCMFGa6T7UySw7RDmkQUU8YFjMw+JTuuGXKWWa7NmKPTXflGnSdEpYR7vQ
WrVhvkAopVpNIvvv78DGQsooWStZKKzlquZMKqSawPJ4v66fNKyEzdaAcGzuQbyB4Gkc30aVR53o
FdY2Hn8+8Lm30WJqZ2DsStJdXvVQB/Eoi19OJVp72T0wxw4vXlmCWkI8loTsD+oa83Ng2ZmBO1Wo
I9t7LuBwpeCrHy7lpTlzWEk/RvqEaXBdwavBVX9tDiGUuBWFqzsEpvWNc5QjFtwH/OA2jycXHaU+
HHIThtTvw39M+UIXShyrIG6p5G/5RLTpDOR4uF0z52k9maHV8mmRLrwMZ8zi7/XEc+OlERItfKga
F5lcXxPHIB6ChB4a8pXg9xi43HgwwHOn2uZMY0hHhFWPmtGkTyS1LFs31+JtRFDHHxO+gknY0gli
+7VYDwiQJsS4Ng4AqV8m1KajCEPkZ9ksJJU1OxFOD5B/mWBrsn+5VQ2AamC5oBtSB5ACZ8rISkXm
SUr9ng30nEqyqKoHvTTAtx/ug7paVX3olkLW0bc9GQT3Kezijgw7heGYPekX5+lMpLHw/Qr4+1zu
bqoHOZGMWEqijKUyXW8NwecZgDpF3u5QSIpUyviuEUVINJrqf6Oudv3tshHoST2Tu28JM+SEROTU
iczHC3cxrdtrJwWbsRoUA/F51DafQYUak4kIlZVQdPgkICwXD7DHH4QyHwVCcfq6vETjBNer6B4Z
VvhyaZ8BOWk7h+VT2Wg1mz/qo8R7i5g23+tLXEgwX92O5jRPibX++5+DqNQkWtMpHIgwnCmP1zKt
Qb3zuUAARCph7i1+E0bfpY344d9wnFzqtkmW1viBNGfanbeVCIp1XX3ojLW3xuO4le83MocQ4LIK
ieQ+2uiieQosyNFSOouC2k7xhpQ+2Fave1qFn+I9bHOoIHTEQcShbv5oK2Ae0JbL/fyafyBnO+iX
b3b6VqJ16+hew+Klw17eevPEqhMk6oNjLdJAVgjQ3+5eaVSH4yy/TtkmVgyow1VsGW88Bqsz3VqE
o7GnXHeHOPoTgvHWViiWB0HFmHU5XXgtjGHJ89tm06yRPrTpEE3m1noqGyziu9ZkKWOkKBU4MiKw
7oK4OQ66RByO5GB9KylVRK3eIgBujXDNsCOzqXZvlkW9TR5FBNoH9A1zLpIj4OVP9nB9MbaB4jJh
RRukh6kCekwPNu6igtEw6y2hOShiOFkfHHzfyB0kR6lsuzyYaS9cXo8OZmJMFAUFxgALqAHkDw7j
K/rV9b/zkHmuqD9FccZppPiijILThLZ+airMtVS5DeRyz46JaIeBspUqYOT9V2HFmZpFxqhSG46R
f7dxxnlm8PqoJfzY8PqmV0rzqnEXcg3zVVv32sE8IsROIEC4y8DFokhz7FEWr6myU63LzS05AyyL
mkTAii72HCqo5CzUp8ALy9FpYaHdWrjXVwLpQjPV6ZSEW5t3IMo1Pw5t+jlrRG4qevXnBB5SfriC
WoVPP7r6fk3M2efufF1qRCxX4WPHKhg2xvgzMXUMmfSBEwFCyMGzuMYDKGRu7SVPmebxzKWRFCDl
5MCIZBf7otI+1NfWdA5GB++4jKkxT7NL5eDRgdKmXq5S7PuA8snZ7jQbI/in/eJ/getTyfIEEvwC
H/o1Alf506xvB1InvnUy52ltHXGjVzulnw72uxom70k/lolRa2Nl/X7cZ7m3c02YdFq6Qaafha84
D1KlW+vS1A98+IEOWOKAEpmqr0Xp0BSdwJU4RbMG3KldO5XepTVfviNiaZM2j14bJn/PQASOumhC
r5Vhkys5k5CHy/818tZO2A+V0HwYVueTGMGaY7/kVYmRu+8qPnz85julRDfjORVHMi/1c+4OlqJ/
BHOJIUxwMui45WkhuN8gRMrkQoxGYdRfJVE7wKRVKN7QcRVExotV8Jted6iRscDQfzr9+JPd0AFY
soRFEjDInJRtZxkVpAUsyMa/bArnYa1yHbSuaMjfc8ymgbEZbgmCrfGmXc4EqGPrcrWsQnRmlXrX
Y09LRmbIbJBwP/D09FsrXFFuDDlNLxhvot+m0naadqxlizn02kI5IFKJOswJA0O/nLgZbQaZ3g1x
y0xvYtZmCu1+XgThL9iByBee674PFWz0Plz2C8zeAZ7xrV9f9imLj3X2/l09CvM0BuF5cby9TQGo
mt/5DK+EsWspv9c7HKU4I63XQAlfpFOxp+g5kKxCeXo3XWHAgf8uB2NfjlMftgTl4kEH+uq/jvH7
0eMZO7cYAVJcCwFSi/B2FfZHf/45zO15XamHt+JWz2QFTzde0l5k1s0QhrodtQ1k+zrgG5+1klUM
Q4GbEX8IW9+WgFKdSWN6qWcNyztMJw9BhIg44e4LWBNrPjJkAss3bUsX9mgyKDf0/n8EXNdVhvdx
bDhSgpfhOk4IbswKRvnAAX9AQNVfhhWbwKdfBM9t3kn/vlRd2hRuDcEgCWwz5DI+7ehw8W25ycOp
tOsURWYF48BOp1tB5E+jR9SsBYvgzRk8RBbaVxXnMWdR1JBd216ZgmAc//VNHciG7pfJNFSKhiPt
KjJ7uWKUV41GFe+X/2TvIPtVYb5eKs0ZyBqwqB2Uc14D5LcD+KLh99bn9J9g6H3WFxuLrBG3J1Z9
gbaV5sfvdnzVTxooU3BfStd2c0IiGI4BjRiEiDcLoYE1ViyTagMkBL+HvnOjN0ASDC2qNn/cMQtx
iVAL1k7GuMEhkOwxifh73KBfyiumvIzoqJMQO4dVRd5Uvp2zOc7IhdtvbNrDu2XyR/QUuGej2XyF
UHMKUCRO6O7Hz/OgVfm3yvUkodE2R185gsrq6ZtZVuZUPxenVCZ4CIFwY4mBXkxlSSYiq9cGexXr
as6iJ6E+v8bSDe+jT0C/ChPkrL9mpAs03AsdmeQfVEBjfRnd9ExqXQ9zUUWD2uFccGGaVTVpQk95
gYOILkInQWtVn6jBR7nh+QUUMQeNBSoTMS/FnlRjo108oV7inxhMcknkfwe6UmAdpP3Elthfh9CI
yT32kaXCmKCHMQXGvLle7EDNoPcoNPPdkrh8ZXajqHwm2yxHKKj+vxqLHnfrCpGczo4LuOBp5EPd
XtqKgIZ6RZ7/98xytD0V5AYRImVrzSJLBpw2x2OAoS9Acz7+4p6WZdHxOG1RsCzBSRCLnja/nYPd
1vtzPKS5rv8AaUjhzsTenTnuHj8utrLi+XgllnqLm25AL5v0Cxh+R73+dYjkFtQGAUYKqrxegfp8
nEf1Avc+J19UqH0JROQVJsaUkNLYCgRjYOffhtC4P5qy/jK31b2K4UmncRj+GAXDxPF5e05EuD7l
qm0hHf9ZPjoZAuaO+fcfqROhf77LjprRh91vCaDixhDhXDW3sLIp83Bj7ZO8Tt6olOWIQzlCCoLt
YInAEZkJSlkDoR+JHOb42anXhJKF1yG8GZg3KE2fCoBhL+uFR24DE7l9HKCwajG7O7c7HRlL742d
q3KkbftiJV6u2mBNHcZN08dxCPA3UZtF7NPBzZ8aW1Kxax5P+U1oEBRXsraRk7OqQl7oH5Ae0E0h
bc2hHduYfzJjs8cikVsmIn2gg/eLLg1ZrJxaG8krqZI23LGm5O+kV91oKP8AgknaZZJICrr+K+En
Nr7AS9B+GruCovUUsVvyBCeWrlnEu1QEC7U9DORbWs1c3iGRgcZxW0StcPiK/mcnMaNN7Cxiu/3q
ReHAe977qgH9aZRoN767zqky0Tw3Ywc21GZbp8D2m/5uVpefdcwo7tiJoZdllOK/YKTE2jIZoI7T
mx4+aRwwWb7FWTH9Bl8Xk5VuJEWoVGMqei8SFcyMS/qJKwCjEZdgmusERypB3MqzgBh0u9N8pzlE
8oBN6UK/ygF9lR/kznlROpVOncA4yBS8Wc4KELgYB4GlkKccywhBFbt3wkZecMzqNDDQDjeywoIy
LzT6odp7roE38sY//UDBQlUPCkV48JL+9UOXBVQMlUII8rTALaD3dmOUYGSZhddtIm1JKcL1CBdg
Ezo7d8H2pKw+TRx3Hs5qkCJehIqRSMCy2rtc841BMzA0dEOg4LYPku69KtQ4foLeMg2SRw+9k2W4
/3uhLQpoX9xmWCptrJplftRO2fZHMBB4jdSOImgIEghR1+uOxKXpSrEbZfh0iVTYP+uaRg/TDbrX
5/D7HAxkJZnWOLgO1/D6qagSESSJNsozk7+PLPYFB0kEwxjNBxpSi/H2kPCBqLsWerYwBhd4Py9n
G8rSZUAeYlhasIMhOm7JtQRDbqTO2uH8rC729DdlyuIJ00/FN0pacs/Z9ca9kd8Iqcj941W2cYEG
GVYbltwSOY1v3A1/jHUCfr+FTfM/wYB1/MsicdkfFuzNDmt4j7tkV+O8NHPKSDGmlAw4w9A1uwO+
1XmCE3M1ZXFABKWq/fPUGUgNpaaH6EDa4HPyDJ0u0Sx0ho/7e/lLdZ5ws0oh7i+AHaADQxNIJ9oR
xEwUvgx6IeptNu63NW61alkKpCyx2K1K3RvfRh/o+PVNh9Jp8qNLE1w5HhlKR6nlG7NCkQoRyD68
Kn1uyfUbuM47Q933vLcF1h7THY25oh/aTiZ3vbs1LFQkVCtMeZwvIPcUBLQ/4GRpOExAj3AG9z+m
Se7oPNuQNteMlf1YEeVjmk99dxWGj6NYj+814ua0wXE6FMJFe5/E8Dethptgq22aUlcFbGBBAJeH
6k7CLuWfmfbTYw45qcw8TQCRfgkadyHN6f33MZNdaz0b4vSuRif/4DHdkTGo8WTETdFbtXXlfWdG
jR1kBgEcyubygOBMyM3bQ7K5mIe5xKGISt+c8MCe+qWUr5HRDvaLokihHJbJH9eBfrvRGlgvtwdl
VYLaoVEg7EeJn+97gHIjrdavbMMF+kY64/13eGcsDSzJdCr/cQXFuWbW1IumInHNqpgAdt4PJhX5
fHNVf7on4tc3r9cIKgRw5MlV92XuSdlfNiWdNps8I4Dvc9DD7gcxUG3qdk6m1CpNxS1u3RXluFG3
GU6BfalH+3MuqtjB4Lwgw2bP2mxaSyN2pvlWWQfh2/QdMpahZR/6fIxuvydtrJTtgTYtLeMTXmeA
ZUPPMBNdUSP0HW4Qj64dtM/nSpX2JUSEkQTR2VZ0vq44IbgQjsxVaUh+1bZNDf/3QzM8l5KTrSCf
tkmhskANE2A4lP2CuwtXrjbezKMqt5zfqjH4znAWsrsRQdrw6Urd7zD/IniiHQSHNp3WdxK4iCvN
u/g4BzGYEyFyia3+MSSJT92Hfv/kXaxXYe+YbNDTS+CzQaRp54VPR0ZvXbBs29zCGwSMEQTkxKSR
SabzqvYAfA2x5zUFBkYrCmNXQQIcvFoD0C4VJZolG2VbBLcx8Z1H0PuEsDgpgthRRfiilInOXzTi
ZejA69yhNpU71t3vzZsYU8QSDU3JEFI0irXrPHbnmgddNCjIBDWMoZQ+qnmTly5DrGrpQwtJ2c8u
sWb5/jzEvgTpG5Cmx1dZ7NGNbAys3DvV/t4+FlCWiPsJz99saR+e0UktM71eO3lA/OHu/cJOOZNz
RbNI9j4D/Bs4YEBrFl+dHj2W1MPYWAtz4JzdG95UeaIHlU7NG7tSRuCgyKt3t9qFRDgRygLsbaxC
CprLK4cuss3ml1Zwk/n79Enuny4cyNAps1ZiKzMrGF8oSccXSlIh0xK7jQj3WQBLUJPwqY83ZdJb
MLhIO6NRfBBz3Bd6stO2JCVqlabnoltDKx5df2PRmeF4cZeoT0wweHyrvW3UFeNaorL44QSKbHpi
Ad2ZYj3WsXIOLTlLLxkydtBNNSDwJEYS3QoY32qZ3F7ycm0sMmHJ/QJsKAq8OfRLKxOZ64WwE6NT
euXlt4botSBjzCmlat8BDqsY2qQrfdnpcr5GUoYYU0UQ8k+idpSJNlY9Ct1YLfqNBV+TA4GYDwGz
QZZ7SiZ3GK58e2CYQQz1Xixdvz7cCD9r5rvs4+laAqrVMbF9B7MJgHTO+EXex7Rgv/p/D/ixVOwJ
aODiNw1bWEQM1Hl1SZy8ET7DbVUTHId541g9McnIX0u8XqQBP6Mb0N3dVkGkM80fvXpcJcInEOmt
4C/QUHwLoPHI1KEuhlFwnNRm7Ej23tKO5yQ5Qpz3RqaZDPVVsEFzj4xoHfe2Hk+aNTFxCFnc4SP6
TjChLPhYmOeXohxhUp6n5x0yGR9iQtYE3g1rOcRF2uu095yqYG4EFmvH4Vs6/VfP6u+iTtcjcVnc
Sl18zy5Vpf3AaoMB9OCWL7Yne2usvaEAvbe0CRjnDOlZFY7F7JYwZASVI5AjpUHBCbGoWSP3J3rw
aN4ZlruRTaybg38+6xTpJ9BLZ19r+YKHI3PnnxfVWrWa7EbMofNI9QarRcdH5Abl9Sb9e2OSaYtd
UgfvxDhYOqnjXJp3EqP6MldNAV0+swTyX5Uq/dS32k6L1quamvcXE+2me9gIZJRRcaXLDDtBYO9B
b+25IOu9IEuN+H9j8+fJS/FXMQqSem7tCSXa+VRQYWpb9+QwIsNjskOJrD8aV7tSlVLbkLH78xHj
Z+cNZsEB5MsKA3Nv0JghgaCIWHWpwfv9sUp5zc5Ug0k3B5bDKJaJdS1XC0lqzg0VykBUNnndXO49
95Nb3XdPdjupHk7ppM61BZ8LEgljQfM93g81mt9XzLsfoEUZ+p4u44CtgKvcfZOFHxSfkXM93rI4
QewgrKLexMRhGccX85A5+7zEgv55JyFD8SE0tx+gkc+DoPrjhtG7i2HLBiu/6y4VilKYYTrjylDA
nmguIPFXgmAuvqrG+UnX+IzO2NUi0X+urD5UiEC9DVfR3F+SMtJ8Kxahsys8xkUnMalxw1KONZxp
a8WyUJEqJxidQkI0C0c69Zo8qPikyHU7XbeLR4SLvmwQwPDpa3gfVW2GC+A/wSNgBukllmOnZWyQ
SBT2qTVMk/f118VI2wgrx1FnW/EAfuADcAOEKSsCvE/QtNWVOTxm4xzU1Va2C1YGmJ0mCjebgqke
MxGMiQu7o8Dcu7TxP+WktSgSHop+DAr+uc0DDymvRc2iypwDDsSc3Immdb+DVhyWzpxIBCbf8aVc
tkw5b5fVV1tihJip6tPuugmwb1u6oLQrMsnXtF3nLLUs3KsFdDXylwrJt0ouuqZfOO5tVk82LdMn
dPAE5Wo+/lK3z7C43lIWroCKuuTpwMGJurwOaqyVBFdiq9gRsw62WpYuYnumh3qJ0SIz2kUEjwSt
DktyOyI+dU9jo1wp6fhwFFz+KTyXY+BCSiM6kHFCf59ueZp+arBfXMjSEjQme5FNXX7Kpo/pD/8W
lIVLXT+ZEo2JcJ9IsK6BCTQRFcJcub/5dA/AHa59T1iRRJfMdGj1nDdl0GoyYXAv+iRIGDnrKl8R
zJ0+T0f3oH6WSDQ9FcLW6uTsq6pPokyvjVVJ6euNogbqo24ufgXywaXHOYkVwbhMmaAx3qfQwZKs
+UakI9aUTEYU7Jo0C09ZFJproOMGbj+mu1e22ryjTWvmFIwtFsy/pca5ZgF0hoDIum73jpk0/Kkw
lwKCVLR5B38u+pJ750EwXL/SlqE/BhrF9mu9VQZ0PYXVA49q4CmoKFwcgvZrMb22vyRAiHSgNZyg
8fqaW8mr10YZzKtTUVDk8rm37WkJ7rUW3F4ywknGUGzUqu3G6mClzymJPfi8KyTRGn9mZyMmutr8
ZXBh4Uld6rUSI8VSSqb5MYsVN5vJiHZzRMKlGU5uZnXTZ+zIj9vNz3oVClruwC3bQwU8owr+IPjp
XtUzNMwyEh0z4h6EsP1mB+TliW6+Sn81OuCaKNsG1jQargcCsICwnycDXHIKv1BPTX9CzILAyW+E
eHwhI7VAQPhkgew/QVEGN/lg0On2XDvkVvCS3+j1UH8dzVNLC9BlR6ndqPCfI5TOfjRtcAhkNA3/
/W3dyDPGUO5Eb9VJMiCgu2ussmGW4mY98caO83rO/2JNZhBgjlWDzjgD8t37NqQZPJla3G/6Npne
H03TWT66j8kR/MyIYTymAjau2j5gtwX2xC4avth1wxTa1R7IqgjIMi/s8jRZ+F2VPYD7Tp1TtEYB
9ySD+l5dJjvWDpE81wOOS3iwR4UFTTokNNqcTg/bFI48aMhan0/HCoGact/ejv4wDOdmqoskCLM4
eFtRHfZjBECxOA6kNJZ2++0fRS4XinIlrqF1o2P24wak3n+CpaTCfqQD5JPYr1YUq9HIWHkxAULV
pw17DJmWiLTIhZAuejUSsc5W8MksCof7ik+41lQF6TcmbQo9AVTK9g2kzLHoFyUPTkwkoBHbfGrD
0pssio0HKebW7+/rPjbHGTr2Vzkbrn8QI+L6/k19BaHLOT4LgJxoGIJuSufhc2vlvLzfsNuXb/NV
e932Ovfn7keIhiYKCQJL0Hq9fdbaMyaDKSvwSoOh55GTccptCP9RUCcvdcCaVnFy+9kz+V88atNB
andhJxFrjIV6M/MrBIl/JY1p4rwO2i4zleeZbg+zSNRLTHdE+RNP9bgW3r19tGPnQUPr5olvjuAR
CBbE6hZ1UkAWm/fXh7qSbqUqCDjMasfjggYwBm+Qr1PihG1XThHvH1hmH/eRMq181ui3LJsiQvCw
TUS8715toh+kZFbfq7+oKFk0ehpetateqsM8hZODofmGJ9ZUIuoO6bGU3vG6MdT3TEoWbiTYoWLT
30oJKg14IhBbw9xosnVLrDTiAwUa9z3lASM2dYrcNBNdNRa4xlAOI5a0VtFEPygQ2S+b0b7UxkKJ
Sf74EePuEnl9NIEDAYTl2Sfq9OPVZrciuC9KSsvrexhSEQ+rBHfq9Ik16BuvfYnt2xVcc9/tJUdx
0o0a+/p6OReOPIs0CIK2bHWn4jfg82zicQIxkz+/9B0vbck+ftXO08+ll6nWdwup0pSKc8CDxGJ3
e9rz4eGfFrXeJeYbg1jfYDx1TWCD9b3wwFdg8qs7SeLzl8Tsbd0aJLTB+r9vn9nOLeKfodYpk9zl
sogxD538unnhOPpMRSdsaQHLeSVBmrAedMtB2539csXW7cbfJfv4W70hHvW/YNNvWSUDznb67p0T
d0hObbiVLZ+PM3yhWSYc/NirJFnXpTruNbvyhulM2I84sIPCdxvy7oOS7rSCX8mHGl2sfr18q6Lj
NYsX1W4Gui/FbMZRS2+WMFWqmHbX4/ytBriO/0ukSHoALXvBQ6THBYAECj3y64abZK3sglEDSpl/
3vK+l0DXWckR6ODlwn6SMdAEKyl3bwoN8k680qYmfZjy4gLcdeDsXW33BQcdpNB9O3vt8iIjOC94
7YehUnmf6rvJ4QKJuLwt/eHdWmI7HilaA/xH64ROXHfO0Gp7SdZYNwqlOts9zJM50q3yOGy4gGbe
hjXZXSUSqGIdlC+9AocDEzKQ555bgWKmV62SHYk49gGrbLonVvgda6eb6TyyDTOMLXeTVHSRc9my
5Fr3Y+paSyVDhOWHPi2zZCi4GyLMvRKF9NEIG4p222i3z82IKrjMF8E5lZXyxnnhiXSyMs3ytrog
qG2B7w0AwcqqRfwQ9x1PJs8PhIWo49l93PVxT2OvAm4ccPRXQcYLNLBlFojUprlyWykbGzRkU/hb
ZOgK5NY77OWChr+D1QAKe1/8I/sQch5K967CFzwKD21/JoaOvvWyzYkpXviFQwcNYmVu6hQTtKcf
9i2ZfwfTiqVEWsddWjcwm9zPtE/xUki+u/PQgbUe/e79Vx6Scr56RvI1cYss1hdJBZFD7qpyYHDm
G4p1Z+WtKqaYDgmbhs+orFQFCXiHJmwmjW4j0pn/ZRZ7XhvFMgRVADHUBzaCNxdx0NgH6BhJSTxU
cwzjzB8Yqyt6uVLM2g9Xu8FzoUWUAjtvRESv6nwR3j/69AmMfYP76RYoyoz/fwq9JaY2bXVpsV/D
ezE7/K4bb4mRNARBQQ1/7iDaL/T4EbJLw0Eut5P9kS2e5EdeF4LoB9AR3WeFUudjKXQh/oJRtN8p
gFU1uXegS5ktKRMrOKU+qT0NNCrcnr6qTWT6fu5Pu5zH4gBDI5HFTDC9JoIkyX6k7M8XNEjH/Iw1
P7xaMKhL0T3uW5+CUpNy1nKs3NhNsTaoCgGw4sYtEtr4raiBPr7LtCc2FUKyMPVqCmqN2Ey/eA7p
/kxrR7Oeox7vWdu8YQeflEiQqII9RlWa5ykvyQ+FJQLJjGOzUa5vMk9UTNDn1C6JmzPMqV9HD1yC
yATJg1o9SLgEDo4bpD5i3HxlYeL82j7zb5McGEIkAyWAsFuYoC+wz6UF+uYERkHK323UB5oVQ7AY
mLEwNp2jzuGYknlILRxhob3byjHx3xMJnm86f5mxvzoRccukL2UNWnf4MzX5xFYSoaU2HXY3UdP+
D7iZO664UnVHtdfyn4SPvdlWrDCuXgPQ6gQZKj9XeY8gQwiTP/ZXPqoZOJtD35WyRI8oBxXEv2dz
dL2V/g9kpp99bN8aREz51bY8x5gM9i525fnB86HtgZI+c+4GD0JJejz+i2YBX/FlNyAAllfxHzPC
Q0/yi/L1VH3BPpiUtazdCK5NslUWYWjybhZNUXO9CRIsWw+AujoZNTZfxBSMxRdQhXm/u/DOCis9
WNXkLcM/4y3xADqTPeGm9PCBxGu0wdszMYm6NbsxwGjhndO8n5yEq51O0rsTcbEzBvZRvOOAQsOM
/4xmx8X0HN/t0/fqJ2J8flUs3asVxeMP+diZGVwbRC+qoiMJs2sOLRXg7nwTi88NEaGyeQsUusEH
giO1aJ2s+HpfMWQhjxl31oa6hKgdQe9jY9J++EEgCcZAJvQ9U5YDRPE3tm7rjd0BJz+LCT7nagRu
K96iSlF3SFAMM8rl0hwYhDF7mxqhuIt3hcM919BtKvJoy9hcorxzfMiIvYTrWnZz4NLCWwnMz4eU
sptxq3R6yhGwpE0ywcUC5enhc5TaLj4yuzBXy/LZY3dHdNTgIOEIUylBitJJZggeKP77HrZNQoVv
bs/HcjD9hNbDvwgP/VTzutBKJkX24EahwDWOrPQHyBjxexLtrrpE7DDBAIcwiVjc3hAcfsOGADz5
hBgYAfnPn6N2h5UG/IyiI/VA360UVzDuHpLFuaQcy4CXJofpkEGMfaHJvBbSkBuYntTzXSKD91DO
/DPS2WjoBnfsMqGoKtZT0QBCJf21jaNLehbGjJZS8UynSfdAVPul0AEdf2y7dCPkfM0Brnc4GYcA
aknw4GATBDBHTw/4NntGSyRqB8pKe90+BskThmmv7n7mlTG7LVe0GBgDgl5HfWswS31Nsd4e8jPH
PjFtEoCq0NbB96oliNeeeVooBIw+qOWPGsY4paQmCav3LuEZL66tawI7baxgClo8lgRqQezzYVY9
8LgSnaGPV4nX5+iIh45X4P89QVhg02Teya0/+NLvhh2kTZcRY4ZfE0t+HnH5X1rw2OIzLamLU41g
0wwPO6fJKmBn8bYhuC0ze6nouaeo6bXZKY+rxonppPxQ1HG41sU1vJMMEfKvT8XdSszui+U5EfMJ
WdJDMXFyDMrXUXszops9LV1spINeRoxHgaASQqFtGTu0XuD4Fo5E6t0aWLG0WLoUjdAbOTUP3hWL
KrstEh5KO+xKVKEXppnzYnFdXkFlbB3DahHt/MHmoW3vG6bt9XoM+L41XFvcv7zWGQCEqbqCn5oy
SO+HewDQSp28SLsIpoYqAEh3Y/UHVMUESQLa39ner6JvZLQbe/PPC6DDj5oi5T8yxYfHqWC3xjUr
wAEOjR0HrFOfvSlFD/Ampy3TSlAoguIsztI4f3ltW4ygj6F8lfjJTx5uOj4pzFay1tRQOi0bt3Wb
yPGKKvmW+o8iIH/w64g2hJ5ymIh11FU8YPRTwAaH7HeSJljCjvTQsHUX+enywxjE8ZJr3LsWSIcJ
DZmEVxLnpYkvXqYACtUZKEK1aV2pKrKy+rk22QEA4uGKIKe1yEzkWfyb9C3F8TYJNWPxkiI8jnfN
H+5gec2sMlPgUJmIQX55BRkBPd/Jrxq0r4y4FG0vJYQ2KUetUYEIwnaOb3ADW6N7tjTZqtrg8fzg
OeYcBvPA57oaMyGhwYVID/NYUg4mtEg10U+FZMcAqM0RSaUetMatMzMuuQ5Xd5Wq61+g9PkNPjw+
APv5gxO80lD9dknk4GorOQf09uXofFl9CMMlBxDqip/H0pLvQftT2XQA3ttboh9v4VLM7gCeOT32
ZzPXh9K0htH3id2WXuR9bCO2ExBiHz8Atsprk1mT0S9PVTOL97mRvO6llSXkLJe/g89kYeNUmeQG
+b9RVrB5vQn7M13nBs1u7ZhWxHXDJWZFs1LknmIID2Vs11bRo12kPrhXL7B+ji5zN7blg1ZSyb0B
6wh8/Ke+KyqtinOYO3lRKBjNe9bn6yuiCHtRzta8sZ4nOTK90Aj5Pr0v4DWKjvOja4M0KVlLifSl
Jl7MWMUlqGkl84aO6peXmmp735PybYNJ2z3OQthoyZR3sl889770/Tf3dq1BehN4QT4Zl/hrgXt0
NKLJ1WsykzT11YRtwp545m/PHCC4F3YTLcgiKdvPcZ94j6TS7U6m3nA8MToF1MT/zO6Lwt0gVaaT
agHiHdZKh9Qaltp+ZJ8gwIdm8mM+o2PWhvOXA7Ca4ojn9J7oaJqCULNk/eTKGo0xqIQJQR5NAXOJ
QjAeKuDwXnD09qVe3BPlq0cr9E0RAu9w0DZt7Gz0VCf0ojDbgv2igTSi7VbSbg9MqYw4zD/AkM7U
gsy/LvfuqHlcdlnao8VU/MIu9s1nVLk6/EJVRiNdgm0WHzrOjDwyinMTaKR93bd54liqPcOzK7V9
/9f1VvedOqbI6Z4SCSXytaXSJLt47VYjiqkVvZP1EjyBnAa5HYqYyaEUb4N4Fe9D2FGEfCMyDg0v
StQGe42VoulgVh5MNP4N2Visdt+7tccSF7f3wwzRe0MiJdLPbUqQTmMy6hpahErFuv9w/gGmKQLm
h+IL+2d/dous9yb5HS0c8ZB7zyanl1JZ6YeUgFr3Em5mNB5/qbRwgmuEEDmU5GOlIZ+a3xO6U6AD
P/KEeKFOHdo3TNvEKiCaC3CWaKxDhMOZcdYgx+eu18cEt9Z1fDRUk6jywTu0P8r2P29nzPM3SCgJ
Q4T6tBKhVWEcmSumPzmnTkYAct24k1ww3WGoqrD4nCgYt92G+HdsmGp/EyiuVleFEmuztLfTaSi1
z8BLlwgiTy5ARLVDWPRF9G8dPWN2Pn9Po+AeGGpoXPpBFAJh3YL+HhTVNh52Pk3tXhy4zxCi/CJW
l6+06W8cNP6bvXImP+Ajk4D2aKCA65o26vPdL/ZWvs6fHtDPJR7zsgWF1mxIdCMbCXDT1CAppfJA
rxTziSyXWWosmLEF9GhvvetgIZhoDApMkduqq5zjke2Cw1PU1u3XcbgVA3c4+0MhLkpAAgHnYDM5
0RV8/hyayhNvhKp5c1EiHHtV0nZGpJYooLfb44pnryuq8FP2LHjueUKv75O2aECrfg7NWVHGa5If
YxBkQVqmNBN0JIBhtEDhEq9PbrOT8tiEW/Z1RyM7j51Pq2EGg60LVfwbc7JqCyiVCBt4j8plolq6
O7f3AGRLU9lraMUULAZeBMZPf1rREdHjSCvTY2uzj6DxNW++Hy6PhOrY16Xm7mIA9VcFnG9Nl2qh
pqfd8bL81wSia6x2S1DBy/tI5sn39HhPKgmWZZjN+Tvf7zcI5kSTcfokFV37AwRrySXpuxyqXHVF
eBYHNw6KL0pkmqyyDf4ognFBW3VIJjIBO7cBZj0gRyY5qyceAIrp7300ew80jag+rMS6NSANOO0B
/5vIKynFxmA78AWEA43LjKnMV3rh0pNppAW7QfyMSIfrAqglTF99FfrfTkVPmC/aKxNJ3kSXXOUL
YjibLltWTmlHz7yzArJjPkKGqH0kfLyznpeT2LrwuRTwV1LsLIl++HK+4NapugbjdELpUIwPc6fU
mFljg4Q6zhJCsRoxVEqx3OCGJ9cas0BnA6TXrIhv9mu+co3f2soNUteM09Ssl9nnCfMd+fqP+51V
sUKFFPyWnPwUjxIT04HsSlS/WmlKeOYtw3MAOtKrZzodZeEM3UnxXCpVNVIOQm4FML12SEgdzNdD
3igcKZ6C9giT5DLOw5YdpLYrCtkeQRjSMoQ2846g8DOT2AHVogLIlAs+jtuuMrR96wSzXjDMEfFZ
vfYPfV58oNpEeftgjLNenixUxsrcCKqkjTQG85hsrBNHyj4vX9VvkZzPnVmqYbH7pu6v+EYEs3V1
96N0ZfdAqRCZ+m9c7jQeILJCjR+QXv42sfHo9EGi3Esh52KgcecpcjBOVbpFS0yA9HgISTyFYF3/
cuy/mKh9arno3a8hUdpMQgxXOZAXVlKrnY8O9N1JG+rpY9vBW8svOkkMasftQ1OGVSGCk4OORAom
7X3b9EFSldkUrQj/z5joJZkKxLBnVD6kwr83Q0KPjJetdqvJw/dJqz/2JuJ2EXJnstpQE49ljzEh
2HUhsvIsTDBwdrAhi0uL3ccC3XcVkpGRdywd/ITyNOAU48s/LMuzNUWcbKQLe4Ex6CmNVtJUnYbY
FJdm5SaVw8Nbg9UwctT9Qs7HhgLzpitCvhrDH36grhU7mYfYfyMntBcgMHFq9jU4MWARPorpSoue
0jPZFwi4/mL7wjzjEewhk5KEAj1yvkn0s15787L2V/KoPEnj22tP/uDAc088Su1L9k8PUN70nYgJ
5b2FBOYSeDnUyW61geFw6Aco7FNCUr166u67wtR0bVCNDmOoxnxceI7E+Xp6sLniPe2k86Ril2Q2
fkvqwN5K2nnJf8L+LYc7PyURghnHP8qJ5lyN9V7Cw1tN2fTNzQXo4eA0orbNpZ5ShBv0jOOTlJuB
xDcbCSKAmyOEUK0q+KWdWWDU535Y35pdJciiY1JAepan1x/kQgK/0p5bd2dNj3JyXqPE/UspSx24
OnIeIyBr5aLHV44b5qRc/jCM7plv7OGVO0kYGJAyz6yiTfLQVYwExOnKrP+Qpm+WYJ+IVkocim69
uY+xHuxkr2R3gDBf/tXy68Qmw5t9HwPSskvaWBYf/tFwcNB/eBXqe13rfx4nOcMGi09mXc5HMmMc
Bi+//JcDefPNviy7pDlCUdU8o9YXhe+gVsm9Hqbh9ARvrm0MMAFeK9jkbi9rEMtCzGKfK82LrwXJ
QJ8ds5SDGDqwL3ewAn17jJeuPksXGVM3WOdODYuOyVXaHILV8NW54HZagsdKKR7bboTQ8IBlQdZ2
Vcrbyhp4XQ0VnRK3e6A2w8MTHtP/PCNmKYUHuxeA4z+qcUFL/uo3VIVJheBoabxQwCL1IsyLJIJJ
sCattQ6UBVsMj9GOleLik5y+jdxhVP6iZgNaAD7dqyxfkUb+iZkktDlY63JgY6yZNeRkv24fpd+g
gLESLGPa/4ZLgXMWtUZxgHLJCdtqZVwFNLHMZ8hU63t9KxiWo6Tn4nGZPKWaKaKXtqiVFlgONWD6
k2G1MUCrW8o2KPiPK0dUi4ya6wVsgKMFI/dyKoA7BeOMGwZkpS5QpmotzZdt1ZgsL/3PbeMaufCk
L2weNrYBCr6ov4tzmz2qXCGgvyc0rkLpzJXDFJBlw/WpUb7S96/iwGI8PeCApdat4mQrwC9nF6XB
WWzisxXybhu5PB6rJlaFzQxqv9rneKzzGLFBQ/t3tm58fQIjvIo7fj7ADfDwDfO/sdsIPW8lVHn4
rhajiW32PTmRNo3lOptnTyPBgBtkoWfS8nasVaX7/ZiQrPWRgqmCKBzZPIhlhJf5z5ihXp0/wStA
Ks5L3CdgBEy1AuV0NUaIO2XHUJHhTR/6CgQw2Xoxrb2YjH+QUQ0qCdS2Y08lo8AIUXekmTGFH1vv
1oOMpEQu5/KRIn83L+clOZ4j5FI9rZjqA0bvVh8w0oGXQvmHxpG6Ld38f0pF98db182FzPp7M4qo
T5P5/0ZW+gaW0Rk5ulu/IJrtMMTJDFixXRLr3lm6ocwYICaQvaEqVR/zRAuEZmK/Tp60bn5H2yh7
8Qo4coMEOyO3cYZ9S7pww0pSOo1X+TL8CHxYLt1/qcTA25x9Nzpk5BtNag1K4AD2HeB45395CK+/
YBw82l3AmQEWdDRFyJEabUVzQa/lmFZEVE1ddiYe/eRCgS314uKiZNzCABqAS5Ym7b1Z9H/+IGx/
pPQxdMC9vA9+HJN0e05gP0q1Iu28GaOEH+qYL8cPDKVWkinoeADKlqqCBDsxrDvaqyx4KPI//O6T
YS+S8TrU+nUr2VeCIOwp69y6TyZxOpIQ3tJAqu6E9woQ73KxNhkYAevs4GXAHA7oLyMsNsrhTP4B
cncNCamHC17mvUw0xUncXI3MCXC+z5WTs/QScRUr6TE2mP1sTkKungHQAswWFxU9fGxHatHeTjO9
XnZTtUpTmk2ljV+oWx+nyOBopNudRf9CGiFeAJ8qx7FsdeinhwThj9yilu8TLPYCeJ9SIoU/LqTt
EQMj14hxMDEKEzDVOvL782Projq87ua8ToPGbv0P7/bpXOToB61hxI55H+OVkDDdNlGffjpjm7v2
IiO0xV4IxvTCRViYwag+4+XoSJ0cb7yMji29I5JjoCH4LyZjxnRqXNdqQO8akEXrmg1W0A2ThRgd
bzof7O7rkvupYDfVF/CckLPp5Ghz+evopSyc0VH0Dl3ksSkcEVUK1bMlAR7K91UCQpKvsLQxRyfo
jVpdWa3/g41hQlnssZh7rie6rA3G7b1qo1Dks5V4WAxvxWQl0yz9eFOPuArkiaGsKMYBnJDg5gYd
TfQG/bBrvrBeJf4DWZ6/pk1XpOAbEcnE0dHA8n0rVO3N+5SxoUC7URX/I2TTVYTVKvM7+zc7jlmS
pXYct78/QBItAgx06tGNvum7x7BJrPFS0D4OhQya4AFMmKs5bKEWZ3fkMnrt7m5VyjB6qgMzRnpN
cE2v/kDVKE/RWboF648wwlEnB/3Pnz5B40EjcoPlkKrRE8ZdaLrwl4NNBzECGm5dzM5BMAYMPIfo
lroFOkUT3KvExogIjNO5oD+FPe9QO0PJRA1JxlM8xEYLngQ8m2CM4o/Ak0EBEmezKEoHYryHI0Lx
+7Ww8blS5IGMgPXJL0PZjX201Zx9jJUCFDIgjgR1bM/KU3YG5greFDIabtOKukJir48H+4OVWYeg
z/V2Qu3n9Rlfj+D79Z74AGXEUlYClYaocdsZHqzXg6T0MWBUbNB9vwEKfFZFU0C9KXwJunfHNXkG
AVO/dPRD1uLO/F0nA50l4Srk1oLagAp3qnhQk04p6upcBi2XewZrzcZJZTAnfWmXwqDmICJwFnb9
pHw79yCIhR5FqtPTlcc6sHN78FPKijgl7wyatC17Py/Ts01ONd03zC0uyWpRBb9obYHpAWXU/O8J
0oUTlAObMXHipjofGgbmtIJzS9hWp8KsvarrFmmy0XWjmpVxbiGQeKmWGCyEQvWElM2aOQ0TmGii
q8XNS2fpvXL25HvMmTt+CA0YxQ9vguKBHN3V8KCo7rzQip66lNMcxfVK+Z6TEs0UaJOawL8fTdwg
oM62CxcSs+s9KkiWzvSvn6YqBJzqARS6Fov7xBCgxsv8ApAUPoo3QNTDKiNKPWSsKmx5Qt7F/YMa
COxXLiUTXzMJ5IXzzQiB7qhRDa/kDEj161W0NtGNlUuKTClqrW+0u6dd+zKR6S4L0ze0ZFsqdH8C
BvfBxe1eHHFPS5+uVb7qmSbM0E28m4mR9ycUo82XuNOMZbBe/SMuESyREgHS7gvJiLgoYRG5ANpf
yGitC0IE3gaMnEnhxSvJzJdDkJXnWRPditzkzz5jDyrvaDJnMItEKaRKprrCVz527mp6oUTbpKBM
2FnWNpNxWHEkUqR6eIFfYhgN5gAzmd5eyINQa61Y0LavYHhcPyowPUcVTFEwXSTuEakcR5JFSNpw
Ndjr/yYOzmfN5jo7BdeTIsNcYh8g8/MWRxARTkKMDkMQ/H8D0q3y9qoscC5YWj1xqUIPMc4Bnh/I
/Ws3GXRa3cBVcfyL87wpQ8Ip99cYIaudM8JApcm91ikmchBw/HgdH0HLW01WzA1WT28IlSJauV26
XF+4IDQe46MGxQ4G9li/y+OGF0HSN6Bkr5JAaC+HhuRjvY/yEpJAl1W5AMpPUgpgPSmRIxoYIc+J
EEBoqjEbNprPPZHJ3oUnjjET2TyEXg4ci6QshDpFo9Wcs9dyDFF8dEufg9wsCGGR20ZNeZQA3l9Y
LalGIHIUW6zejUoo0JZdECoyeM57yieFYd8Nw/PeQpyYBqjndya5A8JJQa0G/7yW02nD64uJEpRB
uwzm96aga4RDcqKP1D6Pxm5e6DdiVO4Lip/s+gru3Q3bWeNIQNUoOLdjaPWmtYXtb4SwvzhAryQL
8fp1PRPIe0bZJyl+UyhOpJjmu9i0vtlmlncJKAaulNP1awCtnbVFLRugMtOTBkE7Hj3G8jF6IVPz
r9oMU4amzWk9loZvkTyw5VQcdMNZ8fBahPXcBqhVI883f/sJYMm7VXhrVEE6ODQSY9HtOdF+grCs
WFHi7qEsRtpLepRPGEcRt7qlKhbdgmKJcKXAonXD2WK6bDe9/o0i403T5rwdcA9npyVAESzN/6sW
fpSvRpDhNkf3rGAhII7SkcaFABkPgWqFtPZocvlcyvlHjLeGfU81uoSihu0EUiDY7zaIJJjESjWh
oG6trlT+QWybJl6vNbJTArV9UxDm4Vq6LUV6oB7uq29jgIyPp0yGHVQ+F7fOFk+Ybum6X8AHL9wZ
6rYC1rvZ/o7ZqeiRS7nxlCUn7pwhvYc3S9nBgO3N9/Sm/d62IrkPyYWHGyATdRe6+i+dLzVw2Dvc
kt5TAR3t1vF6aVK7tHpLa+FFr1hBOZMKGCGkCm2mxLkkWwMrTtNcxG5v5a3JrdkzPgj6DgAwcpK0
e3jbClE/D5OnBaqaBDcHB4ypBpL6PhUYFOuTW16IHISXnh33ibu+ulZYJ5W/ft9JInAij/2GhCbe
u9CHRK0hfPy+6HoxdQKK4rMLOQ8nNLXlRSsEj/9S1RWrs1gtmMG/63tbN/yyXDeC/Ow78Y6JLmLZ
zhVatN1TuJnEeTFlpLkpnT3QP84OpoyvrAr8iCu2am2UGm/uT0NcqzrckrMovg980HzJTh1HM/2V
Zx//Mf3UxaeCXf3+DJwb/4OIjGpexxNb55BsBc7K60Kr317GT5VULlmveYRmmnTqKaGg8CYUIFDV
UVum/VnKJRFMdaAAfNUMemCGAS8urBV9f1spty5HB+WZCWe+NpeDNZhYNJGH6aMD4G23kAouRLiz
mqioH+evihv3vV6PIr9APq598mjtabSLmyglvaRXqrEDw8+J8D9VWR0sSoqV9Jteg/RhX4fFXRy3
RJXFixI6/fqPUTKeMpcuniumQbsFMd3Obq7No929Rs5EaERRNgZ7dNaUywP7e6iviVzFT56faBcy
rdxZqkFOzNgOpAuFogyqnfj5VZ8W6LLWVEDK2z0Tszwvn8Fep8mZoF4NU40TqcJiAWp6+7/4q6lJ
qEuqVHM9VhIf2mC1R/RQcJJxDhhWz1GH0j3BjsozmDU2KxAF7S/Nhte37C1VA/j2wcy3UioZCHkg
bw20QIqj8UJCE/YwORx71op1ZRcWE2/GS58xj4IbLu+uzVZfI5ytgiUFwsKGegNibHngtZOaIp6o
xVFGfXxtEeY4ODfzXJPwYdMdA1vGJmhI2X4THCkp8HayurLD5jA/36vEwVyymYZT8H0cvGXLFRsI
+H3BOxJ5x647cVLYJ7foHyMg4UNrcTmldfjtVf+q8iL6hKEa04qawOQI1x3zYf8OXOxkQhVYZ4ri
oATVlW+ch8/3V1PxoK+5WiBqXhXNwj7vu3+qdy5VoZAh/YFCJ6Qovv437IY4quP2nEK8oLYWXUw3
yvIe9YGy3qKAjvNaO6e7tuIKF6+LMmIKN/mENBfNO9VWPzVifHDlIdB0YUrf+xyehUJtgzqVOA26
cz5U71J0syK7RGdz8LCi9WM1y3NNwD4dbH8zp5bdGMNd3zOK1SYDwfEta33dENgUhXPc3MB/7sB5
hUZc3KLGZFMIC7SNGdeqNB5XxWnNlHXgZWZ7vTigSazais7iHUFFnKSHzGfzXmwcDZJKjiDUM2kB
B5EaAAGFEvNEBxLDQ2VaHtJchqPJnQA1FNW3V7NU4y/tvyUR+6NH/BtTYE8Dtu1YpL+RGa48cfTs
Wpa34A7WTSxIJaEFGtyMSdz30595+h3h5LWmoJnvCcldOXOesXlazdYm/+dINnxLypuD2fqSELnW
lW56O8s9JON4SR7dPtL53ZnEiYb5DK75p6D3RZQ1lhj5GzBhBevE9g7R5ywLXXumNGqq+OSkN5xG
YsrG5svAyWH2Nq/s1OjEA1rnMlRDaoSz5p0cIGftd02YJ8DuuQti/fw5FMhQb8150zJLRonE5DYl
lgPTgwLGIfqCQimvtpIT5uQhMH+0x6vW9zj9RhELxavbdkLrgFn28PuILljvKtP1WmDa7FblR5R5
qIYkFlU3j3HJAmJyCYQ3ikQnWNY2SN6szBj/BkyNRxynuQ0sX1TFVWphxgUsiPxZSlsZcOquaSze
pLVqCcUFEJYQEPEHSgyaVZ+f5+9g/G1AVW/PjdlUzQ1m6AJLT0rNDDCET6T+QsZ3ebfC30YglERC
rE7zCPov+9oDtEASQGMrS8rZs3GD51ET8dKUbd6kU+T/5jagGI1qiNTtTabh9Z1NixCFtlMp/MLu
4bSdVcYMrTUcVbNPEyCzRMBCXAywMxqEVGj6uTqDLPGyjI3DnO7XqGHHdGHDabo4UCV4X2EidtJ3
JoeDWeVnOVG2/kKlVeaRrflhrzAaZk2lOQMhhYYUeItk2eAfbxYkFomhC49y9xiaV9mdVUCvdrph
p1q92b5iRKJ/WLkwk6ppQTPtPr3GgOoCSFv8vleyHu8YXwFBzPMfRDu3fUPHoMzo04dU34G+nlwu
V1ckdmVaPN2V32uHZn/kA2lhjsBjkNpZurskWph5+3/KamjWo2qmBdHRd0mfYcvJeL+U9NBJLdK1
DMcLDefDKDhV3zqFTC++iGJ1lK4Bat3EDnIKNtNi1DqgAW9VgILf2d8RVp3JMLaHcFqKWq9qb0Kx
FqoV3YkVy+dhVrzQBUClLAtw/pJ4YD2R0lNdtOTxmVEQEx2woDt5Vs/jthdvhwtGETVXJ7UrUFOS
aT6lIlZS2z/qBPVQ/P3j782S0PLc2W5OpGTmMfgMjsBhfOlvXu5TbxU1FQjErbyv349QiOMRwOit
co78Oikp5Vw9tV/AC13hFvZO7qWDnw8zAUpeF/6ikdpUEsbXM/Qfaj/nQKDUd9BRHrAurXt5db5f
C0cxB9EFPe1VInoBAB7++W5KyrRS+y5rPPAINYnIT73uTgGA3XnAcmzOVZ1JXXAeSNg3i5sX+t32
NW/2kx0AdAst28hfJNecOiJe57uCAwHelmZkht52TxQyfqioXzVkM4Db6pbK81aCjhIvFoqL56y8
U9f7PSIXzyQDTz6IkiGa3rjTGe0fFa9a+tbm5J+DWLDGve2fCOD7sC7Fk1om3OOUAgAc0NrJ6nEF
6sE2o6CCeUdeLNgBI3yN9IRQZgM7G60V6KOTRKvB1LQFqfHgoJO7TE8YGGLPyD40WJnbVVqKjifi
DW+hwpkasQLKznNfxCY+gieOk0fZIIpty7RWevdS0MczdN8Lv00vzSmz5rdperZ17WWDzpRHFNfl
LGdO9yVgu8wWHyXKm9frbSjk/uY9TX7aUi/opVEi0cbCICQB2zOYNy79JrA+mqkPSqOTcjcZmu03
GY6wUejzQk5R+1h5HpqQ04M1TB2nFpTxbw/TFcqc/fKTJ/se/7gjmWWxRignzbBe5Uc8A9rPqFt5
n2E4OGfPVwGWsMtQrFMq2RNOTjn4KZ+65TEmQERguyl+jvS4B2JuiRARyi52+vfkNzzszINujAH8
9/EX4g4s4T/1pOwzvGxZpRbld7J81O6JlqdSPIybtg0/jJTFN3mQt4z7siIhZ2Iza6iACWcGcOje
WhnXjtcv1ACZkVVj+4T+GBnlpWtPoULF8uUovjgAncLms2MQnuGggGa2J04fCx6pzO7BUMOVHS1p
UZH4k7QB4A70+Ud8Lpzy9ccvUGt8QYTHcAA1otgYzdmL9klbMCzGUBCQNWQIZyreL1xST4UKudRs
ppDv+9KWGWZvyMnzYUSA3dWjJAx7X4SJlKQg6Ojdz5w4vYP9dqdfxgo9ubCx6RheUEQVXACYEECf
wwH+lvZ5mjEunm6acU3w+iz0KEmQgeev+w1p1ONy3j5xSrd6B/6QB40VdSApBYEmXw+7V02wgrkz
mQaEylvXcRoxbF6eSp5uHnBzXA58X84EXz5aeDkHD9n2eQVOdUS5QPFXl2N3Qu6X9NJE4GwLPOt+
raMzHSYFIVhoAE8cYDC/jpLfcxS9srZWf4pX+9tAhf1ZFhtS5Fs8PzJRGWbUv0t51cKzXLAgucdy
UfG8X3Xend9mY90/p0dCQyAz6QRArehxfjQiaNY60gYBWociJrqOBsCfRPpGezNByz7LYbZUJ6iV
NlcjxFJntZ4Zhm/IHM49RZ6CBglR8JDp/gCTRbAjHiEvgZFJuLg7jVGpdxY5/Se05gO90iM3smHU
NqE3g9n3Fo8qWu8Ofe1+WOCRzdtn1AZLp6DyPcIDWkG6MmCwtENZqDcg15b2G3M4ombcmpdvLWaT
67lSyIOGkw3dNCNdM3qCvnDoxDZq8fNolPY00mXuCdNucbQAEM1OMVKNvnnOHlJZRO4I6OMla7YG
KVEuRJqFDN68jbyVZ3YWerH67DQ9T6lWKu+Vu9CdG6k6Rpz67iv5h55bzmTKpVnI21uxA42ybR2k
52EcyibRM2Ljfkr+v2gRDsHLWFpkttQiZAoycKITQEJQ7aspyGuJEKrobSVlonkdjFjUQeR+GfxV
KNmNgC3qegyOIQ4fu0H6y7/2owNP4h8hKYXUam8yyjgtrjTRwfKvNkpzQs+YG6RzGMlpkENqcX7c
4mo/ygvi5m5dth2iCwKGCgPQO2WRcMV36hR53gUM7gS9axLVjIVlB56zM40OAFfvWPc7SyONKeRh
G0j2taY/qc51yMZo1v32QOkl77iyCJYshzB0RYtppwY4dpBc1+vMHgMqqXDT7NsLv6ejWliGfsWD
3zpkUNl9mDbIyUSx9ftHY4zizM9y99D5uLVr2r/Qa0+EgsYqj1Q5ONO9ZPMylT1j1gv5M8mnJkMQ
b47CdeOQ0bSkDTOlsY0oMXuISFo9vtkkV5PClvF/T4LW/1Cy8O09gZsIrK+QHIObBr4WVpeT415C
EL+ySjsIF3kNdBySb9DfbjCMm59wGATK2CkeRE9qMqs1ORO0HkaUL3gbxfe9Uoaa2Hkmv7Tq9qj0
2JY4+Kn6JG8d8pNxgKKSTar2fMKoNd4GOpXUGL52ybxKGazqTHYUIUxbvmJ0rEXBs61ZQ6Z7+zdr
g5infpRVx3TRxBQxpIWWXRllCD+33ryMeJm8fC9KW8EAywnOiX/S5IJxn/sOVeE+3Fkb5Lox3ytj
IW2bzh2S74yUuLPCDzbrbd+JLZp9eD9ipxPwiFblxM/FhvRJcEnWdtNgKSUS9kZKlLB/cuc5dd/H
ErA81j/USHRQVZ9WnUQmUlab4QMcdeLIILZWLT9WBZXkx1GhlKzFxnEg2egQlhuxxJ+2cVJa6Bj7
xtQRaQrnSNE2kFh2IGcX+wPC++o6yikSqjMZCxnxJKKBBZ5H3bvpdEjsSJ37FRaaGkw9ybTb6vcR
2HdpO7N2o7eq6xb7E9ust77vkDg3hWChFWXs5ZGiODrEiLevulOLPwFf5aNYqlNweLPPEsqtiFwc
teQPiWbfWyRzO1gPQq5kQMK+wynBQwsFSWF/VC6iYZgdrNxYH1FJZgkR7McH0q5l7t5ia5FjqoT9
GEfRrlnruQ86jyHrYzOj6Wdslxz7UpWJvETbRqN23Ymnb6fzOn8FLeCAfKsg6lpBxDI0l0y9d3Q0
31t/GOFqZtumb0pVWRRCZBkDm0yL20G2ia2ICtOtL5u1fscUW1P+IJdlSJ5kZU4CYCit7qVynX1v
jXaujIT1NZuprr4sC3Q7pPckwShH+C6zsSn5qYaPPN1GfMXq7dTlRAfdGS0tONBURjYBI1PsRVVK
hxnA8saFtVw04CFVXM4yXBwVPOVKFvnPvsT2yIphNOycfKei8AezFFFw5CCXZ5L6KhExTCfQoXDd
rrC2JhGWUFHZkPl4c8isWPwUeQj/rZzYWu6EAZSGfA67ckVpKkSCooCkdIaxTFgRqsVotPBCtGVD
rCvdGVRnhDbsywLQTETwZFZ101RivMiunSd4E2nRxlW8AT5Z6YJ70C1HyvRy2Otb9DQBSBYh9/wj
+RG/QCDYISv5L/ku5zcnk+CRsKgw136xqZjEQCeC1L3a7uCjPfOzlVoSqVaMNNWFBgSF4TZVbzPu
hng6Hpcw6FsKuVIk6ZbQ2SBrqIAyUmIJhKfrFET1VDIX0937j+jle+GMjXTR0MhGkJAOqh9rEKVr
VCbTVBXZG0oy3Hd1Qpjt1LrEtq1djX1dtWIfCnlJHeD6MGEYgrAcrmWB72886VUKC3tbztBpLqYo
HPh9RGR6QJhIp4UtYIXtkaYD4gn5Oc7gBmq3ZkUABqG4M8nOHGSAIH406TnB7gPmhLnEdjoRYJ/n
K/n2k3g9nr/Xh7JkS+TscO//HSTH+5GbzLgWfNHUUdsjvvfMYBp6ghQJsulpSK+ktYNnbRiOZFuk
18Lni+LdCF2yiuLcty5pcRsJDE0ri3C+HZf0IyhLnbBRSqehvv1GYtlv0RiFDXj+jPbCDPhMpTs+
owgArO3nIK1UfQgrq2jUnt2uO17dZJaxgaMgrYL3Tmmmcom7aPJu+1SxtXcaLBy58S5sGa/HGRJO
+OBGOjIz0SnuSdlbxe9rIfMAp+sBHU1Knk9UltwoZHZ+xUagwcF9DrwJHlPL1sVMA6m5e+2T1cQ8
q81W3E93Gpzx7fvmDckwpXsj6h0HQg4cJqIShKdKzmji7/BohOwQdwgdYB8k12Khxl2tpXJ0qMQt
B73papma7DWZQE1nbkxa2ID3wEk+jqkltcE3Yv9t2tV1QO1wOcxR74VxhC+6ezlhsNoJDNwxbIN+
n7yrnavujA7+1JP9tFDaAYWz2fcZGwszj6wTEZUj5rmfKpOvFvxWG7CZ6St5/0EmQoyU6Q+dkQyf
xy1kpp1vst4YG+HxOc74sJijcA0DmYGJYxOTsHA9jjTEm1VKZpjVoHnbkTnK2gfgyO3RfXOm8yZU
IT3rNhynoanmZaMTQLJjMCSF+KFksQrf+ahUMGd2KJPPrT+3b5nnleqa4rZW8KAQYLUgDIVIAGVX
qk59wgDznq11Ib79HbF26/XKunoOleNn64ggeVEdNVLD2EV9wrEw1HUoG+Aa9/5WC9qUql5VlZ9E
vmzjSyQb97tOIkgC8AqctZ9DcSdCigTMuUW8x+PUzQ+/ueOE8lvRTYNspNDZzcVxruHp0AWAur7V
0f5/Q2fl65Evx/DM/26M8PVY+dZFYVJ0IuyACNtldS/hy9xJ/5e8kfEcOgq2g/jG6UtkhdZhrgjF
0ZtK9kd8TyP0C3CCmHm062SYGDBttybBsMyAYmUHFK2VsKwT6IQsc0BiAswwEtogJIOTl21ki+4t
4Ihmy1cFBsppIWG2RgAReDWXIONlqzSN4HyBym+ApsUdg9jbpoJKVPjdmrgxThTDHp2Bew3uY+qo
BfvBsh9Bkf7QGo/040xkI22KdhuAekzGgd7m2MkmRQrMtquHiDwd8BTRtzByOYdw8qe9lMlTVQNZ
9nyb3adyAa0cpeldYCmQcX9IfVX7FxJJ0hNUHlBB+yOVB50aJ6cERzGGwK1m5fT4SQaC1B5Vhbxn
OOlyJ4+mfiSKWWGjysRzuYDH76ZaMGajNg4ZFTuAFNM/NTQlJCAuMoeHxXAqBqpgia7ZtkIvU5AT
qAeQ9Jf/p3CYTe2Cb6VvBTEQPD7XvM+XOL8Y+F1Sd/CL2VZZU+WJA217pCILDuhsJ1e1j4O9nBfz
EAtD0HwWl7DOLpop7nllG8K+eIJiVZ1yOqLDOmpAPxf8pE6nymfmrwLxK+xf3AKPoHm8s2syNuhh
HYqsBm67O3x1huWYz08G9v80p4KBb0IPHMTYjh3L3r7lcfYu4sYxqsIAgj2MaUjTpNxLpy8SrfSc
6JPLgkYVg13m3+RaWNUmoshSqbir7NrLAx7BM9erOD+4x7NZH5zXxpxKXJ3pKOdA+m03Rcc7ObVT
wXVOunNZtLl3lfF+QxlxSVY4puvIux/bl8NcUk10eaF/61j1SL+5zPz9rcnYYwGuQWiucvIY4Olr
HRV9FbLxU+Xf55Cho09Aey9kUVtn+WInO/ONXSrmAEebnZQjaEWlH+TFf4+0KuYTs01b7Lume1DU
5SU1g3lEsmmRFA9uZ8gT5hTrwyCsmjQtIynzUzyCN1ZAUoRvcaWOBd98HSgWPM+Dbc9QB2EeuWsI
DTGBZZpXU846YRVr6zYEXgEFrgEuS2+acG0sVFULeS/ZGA9vqUeNdoDFWBihE2ngOnM9Kfe3bgm5
nTMfk/sBW10AABmX6IHagyyiul8UfX3egDyRaqFZM1sFBLlSPqI1KyV8foP5bhp0SXDUHKhRl9PQ
SwJsJBcK6TFWW0Opnf1SCfRajY/wUus0aTkhOPygpYxVGO6zuJmedXdMqI/4Uaj+HiXZxojLqDuW
QDFqGy/byc/eIrnwGaHtM7NWsuWe+OZ4lC62QGbl6OwFcJ0dSlvCj2mFeKaSOobBLAooaWqR0Idx
VgVcJoR/W75TJL/BtQU0dmAz5o/hcYOuZEKFZRbfmenKoC7ix21kqgVA7kgUtSoHzdbY6dgSBk4I
EBoh3vpcS+u4qyPsENijGsCQMJyGfeRQ3QEU2hfActc7pspfgHRq+dSd014MYMVcDkujzHCAjdQl
YEy6HqDlHwrtw3d9uDrvytsLpgxL3g/8Ip1669TDC0aHT+h7frD0iVfk6oH8gI+UBwNW527b4Ilz
QaDvGsN9cVmpFS9eYJXrrEFIYaMHYeKtKFv+ozTKk1ZQ/XSI8ih51KUE8wzi3AP7n+AiReVkt/F1
JqMoEsnEmXKQyKOsOFsaLeLZuJpCQC2Afoxv124rVYzsGo4RmavfzthD7M4XuQxD5QTNAcSi0kmH
64YyBOUvg9VAlQ8SlRpYMNU1k26SqAuKlQp9ZT4SXy4Ff828veVuJt7ImlwKNW6frmUIfTNiZjOX
aae4/JATIWJhmSPjxRHJ0lGa765zLdCa7R5HR6T4Viyz5AHK9GAS1IXs/Oexg29ImE0PzCIK/rhJ
96extWnG0ONjan6n/jILaINt7X0Zgh49DWVPJdCTKsIzvU5tSNBjiO/VqQ/EmDaiL9GOWF+3Ca2f
2cezjqoklb49P/jYRK19iPE4+bwtoXJjGBauQa3m/gFpn7uzRUeyvtpgZwDneJaStATXXSspHPSq
+DlxwDaz0xmb6FZNEDMBdOc0YShT+/zF8Fw+WYtRDGms2HIYmpeBgnrwe1BXFfS4GHbHfak7K6/l
Zc/GK9HZGc+a3Y/FLi3jhbKJQQOMq++sluGMiD1/H9stqejoy/IjdngF3SwGfm2qTw+eYcnfUJGf
nZHiB5iLS58SIo4WrTxvSySNmS/0Ep2AjI4P1Pj42GI4unkGiooihcr5zRnXEg4lApQbwaK9DQIN
dm4Ul8xfMdUMERxpltam8RKZ0+pU6WN1O3LWZbUfYQraqC1QK9z5KyB9NZ9bCwXBgbC7SYvpd2UM
CP0LuW1zMcL/N41jN8ZwvGpVG1jGIjdPkv9lh+nZ/MNP5OzXwZ7xnDvGY2DQJiUrT+AkoeWDxilw
rJvp1u/igFEZVH9XmE0zW+vPzUDDi0cb4TjSBAcoO7IW2mJHtN1SnPdfmJlxNd5TpxgKzAfy3cjJ
XIeFca06wKHj0kiQPaofhC9yW0Q0nHVMUGlWl5BkHEhUNJ1DYtnUnTm8sedF5WxpPJahIBPfxAF+
jZbWAe3GKFEmRZf5c5akGLThlsUm41vZAQQ3kctWAZKZ+M3h6e50CCSLN2uEM9SLjHhHednCfmS/
1DKsHNis8/e++41inx30DkfOQ4LSgoqOBxJib0+luFRf4AeWyaXcf0jw8/ofggWslm/4rhVrK5QW
odkqIvdl5IXtq0nzryXN8ELGpSPW8ssMBcCU///ZLf1Ml0svmU7GCgGfndAbp80h2jalvlwU/xW0
qwAjoxf8Tlm6ruIofpRopH3gVSb4LTVxtdf0vf686yggxYCYPXFOPnZy6+OmbV+oZqirw3h/yW1V
9VfOTCrEhoXO5+CrBY9ISqrNp3UChzhIMDM9fCpluPVaTEfICQLjMF5A4bDDXJqnKZcdJahIZBYP
8wqwoYlJrYEWH1f51fi46b1jZ9PdufSptAnXgqWcWXAT8CKQwxESLN9Thd37C0OU3RN6Y+7XUCqS
r2Sc9C75G9QvSH1KIsZJNKV1D3kru2xD7TIly9QtOO8aG2wd+sTOYJxeN9Wbr+Q+LyjukGzQNYfI
z95DnwiGvQD8l8cCbyGKntcFHTVzXdE4c97yW+SThDoRTE/JrSxkfV4ILMOa2912PNtsUIwmx8Am
Z43U2J8etM+Txb0p0HIDe1pYFDcDbffGjhjDJ5XmiFpCuqZbVmZjwmkJz14/moO1Qw0Lwot9oc54
PL7bKEm0veBpF4Tm9BSu95jr3Zkwod9VmzJ3tElUc6CLgmWpupnOWGAh9XXh9BTfDq5uUC3kJ8Xh
cBG5XEydbSAvjPartXGI1L3y5ce5a8l+vuzENPlM7njhjk1P3tfFHH3QpELGQhRLApZDeBVYPqWR
Pjd7B2pzjVu8AgVvvhr1wFoCSTBbpaAhghE+w9l0p4owYkRTLHdm+LjfVIK1GXTnmldIEo5b1wr1
L4F/jBP5P/HdoHtPHDGcMwkwZB7lM1dN3HyPj/YioQaBxjOzp/rh1PbsxYSZJ3dNcWtsHI8edihX
S9+am8XPgsPhDCGYm2XLbJuxbBWHyR4soL89vSey+hcqL5TnhXy6/YmE/hwDyOKE3An6F9W0kYby
o7qooakX5GsyLAYU4yk6DvqEiG3VHA5KTEYULTgYV0LP0Q9yYHelIBRewBjAHKp+pwJsscIhHQtD
UiM1nyf3qzCE+z4Y2cm6B3XvemQX6bqfr81xOVtyzdvbc9du0GOGjAxA1HoPCQIvTNxcbHkSPhFK
o392DI9B5I/WtnKV+al5/fOKF5fg40784x96PMpG6U5igGOFjfOkMYUPomOiej9VjQYrSXLfZQJW
xEvM035CBMTgb/NdIuzzSMNA+4KgK5+eDcH72r6u2Gw9HkS/uB23au+DNGst7+f4d/6OAcQdBjdq
1Raxyj7Fg42lSPNhMwPLaIoJN9GDRcOkW3cmaC+qFqzkLQs21GjRqCGxG0lRNzEL3TODOn8o1LLJ
sn2r8qfX4TJYKnk1guZTXbDtGOiuUmCr1/GlN8tX96QtZW3RkT+BwOhL0nuI+hSCZym34uRcaXzZ
zN8HzYgG3LD84ZNHoZb3PqFk+KhaZFRYPRCVwqanPhxJuGBt9cZGfDUWS+d7mJe7luGMbtYn9PoX
i7cFFsIF1I7YHhfRPbTTepnx72b/HqgZUnj7rf5ch+8w5itAkxHNMsXgQxwOjJwv6QO9holgbH8n
Vap/6eyACLrob+2nJJfIi01S3EYBm5UKHScxmIqSzIasF60Nz+R7DFatKWyBSDqtlYvbcVopmLYw
oRRe7WAL8TnwbJV89gs3Lp+oIGVN/Ti/mbW24lFbqtNJErw3JSSG0ANpPd39blQsKx7CDWB/TFUJ
tnMuksg6rojjW/YBk4dC0eLx/rfCeRmGaKwUpgaMLFC+pi6n+bmsD+I649lw5xM7lUiYqE3gAoL5
VOuN52GgP/gXTTDGy7fafRjlY/W+HEAs9tSPdDhIrgebGhzSZ07bI9JJ91BigjGLrTCuZtJ1yRzE
/5sBG0xnUaobTnW8FHKOgVsJlr+zfWkSjHdRDinE0I/e8LRNH1xxDhoCntEqemnXnC2TO9z3sjn8
e8PMoSvuNxNk1tDnjkgtJPdDMPaXoo1iVfBIFfQnaxqEVIWDYCvAIOj7YWAGdX58LVN9orTbkRum
6sU7ep7OxQq/KvhprW8gnuxktIg7b1zXBqkqcWT6M4ptPcB9fwu6Fa+5rYacPCQS4yg7KfdbtBEc
O8nGj1UBkmgZiwsiUPzagn/jsDZTYiPPT5VnyYXddCIsQmMKRaT4CgFYiMQUqotEW34zsIiYfmoJ
qeAHfSPie3qjJbxp/4V0Bc89PSjhows9rifCSAhIvZKbB7L41SrDgeVarys+8sXDl0X26i6wAbbA
JQiEd3Ku8h5RESzJ2E26GmvIjH9HQaYFbDELkYEJXeOZa2fQwp8Y00J5SBh0aOTuNTusn11zMvgd
lkW6yr4NGU6HVyfXf3zCiQAeoAYijDAJpm5KTuX46fewWrZMbDwG35LMlL3hNUWCDQeA1a5Y9Icx
PLQ3vu4/yrDeLQLwaTQH+wumsbfgQapdYonLnM/42PxcyhwQrLuwZULRDilmnakRYTEoXIe7H48B
G5/Xo3x3NYmLJPB+l6DiLUFmdnJdvYG4uLr0OKlhtkQGUvIQ/5tgISCT5PT6lpRYQG7NiPNm3XML
gzvEt6005JqQoDelfHP1zjFWaE23FAnsXjieXvrDiIZgi1Jldna09YFt+j/nSKyXUSkQlZ4B2ZyX
eEjcCSgsA2Q7WqSs52RgCuqgdNi8+7NWmuuB3HYVaHs9ir72UvuBYyr460JOkEf3QmSajiHdHZvi
+T01Ei73oTku6D/1pv0rM0EHG1wHQdSARiZM9Xnsim/u3aompn0XZjfMdCfzZNDmxCwlC959S0lL
bGnGC/uJ49RCJGstY4NiBt6IdOB1+Y6m5sIesKwWhorvTlkvifSmDU1uX0vp47gAxPrMOw81APqG
pQXnisJC6WZ2hjL7grXL94JRceb0xBzC6PfGLk3+Y/V4DcwwP4gyYoLX8uI4hDsN5r/j7PazKiPo
7LCisHmhJaIIUehNewWvMuVszfrF5rvh1IARw6rljgGnn3ite1f/GujsUgcG1yGXMmRr6UKjtiL1
Pcq8wA6G3HTx6iKszzJ/GTLTKkfMQnuYS4fEQShVQgRyITCVp1+gzkYjOAQBhWcCDuWcjN+HDrEr
NV8xvWSLQI3nXm6HFOm9WjJbeyfLOexCqt4N6r+D97fGIpFiVFPtctTonQJ9IIIPN8sjtUOhz7Q8
OU0+28bco/pSICJO+g0DpBnig/dwTEXVQXmMyYkuRntgLk8oUfeF3VLMPTOqZcE8MKBmMO5/ROEJ
7kqc/1pKzGVCY6Z6h3zG3cI2ZkFjh3fmFyXwd1t/tK/P/5aouqimbGMoLHsMnuRXFaw3zBQrC4AZ
sErYMWYUOfc0VKbPIWHqwHyzs4dvlnBJv73TiKdgc17gC4Y+Lg3jTy+C3zNw9KwYPTq92QeoZKgc
3kjFn/wbmndLz6wQWdns+aladX054jN0eXyVCkjLDFerKmyND/37ELqMydhJou78Eua2nkhRdyPJ
K1u2RLMTEPuGNW0kWBf8nhYfMzML3vPn5ecjTT65fLt1vLqdmA9xcka9+tMFIluvSLdghX+QuBhU
LFEAxrqumoYlrk3APonMmTGBGApdXfro+n/xMtTEKOSQhbqLtFG0FBl5SK7ZphMdydGwMvLmN/Pb
cZklnsa/AXd5PA7as/xEhndgC4iLfMR827kbn+ESvV6QKM3dlsqMAo9cH6V12ViTRVLSZH0inaoy
q6mMcsTSOF5gMs+qU5GpCW5xQ4p4QLFZ6XiozTwMydDOVrA6hNJitC8V/4WLgZB9GRrHGlbEEtSh
U/NCwUh/ILFlraNAw+9s5YdboApVeG/ddALhccGcrfx2KbXESB2yA1nXMXI/u6v7GhwGoBD9Q7cq
DsXRXnvN1pE2h+J98VLKB7MzmmurngFs+vtVu4Kvtby801ehuch5J9AIKaV8ZG9Gc4eq7FrnW9fb
LkEsrXcblcM76VVIaQeuBfR0W0Z+x7NYUxgVxzjnmuDu9bjElgZ8bYdInAgMduWEx0UG36AfOPkD
bUUNEjRiwJ5HqUl4tOVe9rcLv1gelyEWwvF6lP4Fd/x5NBhuq/oqqB3AsO697n3ucZKjOUkLhSoO
QeL5pMU+SYja7WF/Gs2JzuwDuUVHCmpXhjM9/PDJeW+y/39l0kimdLY2QBj9qfDdtZUVjn0pO/9y
TrRbKZnCN6MWrYmzQprAblvilS60MsnA99du2sc7/RvcYyV1M/KVT8QnjwiNs6qihsgo3b1K6qgl
/Yyw8JmirecQ/OIV9AJDO/OJzeYyIfzQeocpWOoLu620jQU8oCqeNaMxS+U3wrmOpYTqRLTSUhCU
1jyQ+jjgmtPUcx5ib8i7KuTUgKblBUUFnmzE+ywHcj4zQihdFKXdQKXNIXl5WNoIBpR8jqt8WlAk
RaUz2EQcxXIgpB1D9jWvdIlwnQVXN20C+MLkOx3Cq3BGNVMfvHabZkdK42fJQ2Ss3k7OK1mGmDwm
lGB/1fOC2JIMd4q8SX8kv5g8FnGeL8IhnacpDZ+I+9hmEyaFY6cEoLb7+6R/wGygWho7N/DfyZdR
Uh/pC+Lbjq6DHqdDdMzAqUTkLrECSXZEoojzinQwUVsok9Jn+i1BcAE4Pto/UkNC3sflDUQ9rQey
4BOjRsXvcXev7V7WuYmww4WATa2sKp6U94FqkWQfExZPM+3QymcSztZF8ZVHK7TDOWPa27/sAsD6
TijGkq5D8bCrou6Sc3s+jG03hwIJSkE0s1DtYIajejJ6Nl3wV3gh9YL0oUvQt871jxrd8DiVq1Tj
lwejnerzmoZyhrIdXEicWME8h9s2IcmMbhzHmNRW1UwZm7M8mGVng5ZsGoOGrnt2Xz2F3pNUsvJ2
Erwjk6bUkJ9mLjOAS7JaE+2yZroqTyLWqqzuxQIIBaudrNYJB8xU7XnQ3dBg1Z22xRu5UYCXXTKS
0KzEDNyo391G2UN39HYeoGkxPwbcC8dvxDTfL8gSQQDO9SJaSw1CrqEiXZJhPT97fOKTGnDjarzi
iN+Tv3A3JjGHWtbK1E0eEEbL7qthFukoAlFNn7N96jAqweTDSgPEJDNvBkYrOtiQiYHVUJcVJQZ1
q68XQ25Y57Z1vWDdSCUVyFuvaVEgk6raCMcQL2D3ne/lElVrvkyaOg30XIGg9iYqBYzSYxqqRB0z
2cPfeCC6rLxRkO9LdR8hKh+9LSYeeSHmA5zMNpDT2xrz1YUt5sxJIGtQbSzwuSTbj99UMOlkTTvs
DQQF/XvAcJBgloQaW6kPGyk4CR73UaBsMitTyPKL51AZb8fOBQ0dlxO4nBrOcyxbqC5Crmx0Q5Ut
QLHV9Nj9NgMOVp/IQspsOjnT/kZieWqacvvtWiB+rr605S++6Kl89SAUAF1IFxd0Dhzd3xT8Gr4N
Ua/brlpJq0/d/Ejy2VDZbKYTV06HAXVMR/E61mWk2TxpzeAZvlqxvlUnuT9GarVqDDt6U44riQm3
dKQd0L4Xp3904R4B4jv7q3bnPJYaNHzfIfLAebND/uAnEEpFSG08SsvD9HUbLSrtK50UN0qe3i/H
BsrKs5KZ6SNUaL2u8rrHrSkIPCmIO2vWgpKdX4ZfRbyytyQUCdoBFISZ7MDaNvVcAXAqFD4xnvFZ
jhzMMYOCVUVeKXqsZHe8Lmv/qyKsbjNKe7lOPN6GDyhhOaGu4Jc9H+L3jZ4U4YCb1Vj8+QgWaflO
2LtAStWFdyG0xz5UQOQFrrsd/qMY5u0ite+K9L7CdH/Jyt6grwR3o/U/xUXWyldzEBaaSnFSA2NS
4wl3hvM9RI8i+nGAjsM550Ct7ZfziaE4DEIqytEYzcxJZwi2QpbP6nDL9W/1RhoV9U6ioX1bNgZP
IgEZ7RB2zwWQM6kh7QJxTzeIPZcmJZ86165JDtU3dpw2rIeSis6BnRUPBL7Se5nyMddRPPvQREW2
kDTQ7w8CsJBDm6l/K7E+7RAiKEA87L04kB4/tksl/pjkYTyA8UgQrVESpIEYwkRyFJkFPPE0R7GF
EebYO/Oz3zjLv/Si/Vxv2kK1mwy0rbY0gtCDzwVBWmb/qNreAu/TvnfSM8yytGJXmpcQTTnJuzfr
B4bz6pSb0MKjWjLTfqrvk78QLiMJcMB40AzbijqvEr07dAbrcavSohBXQASE5qDSuFWsOAQGAAyv
eOQxtV89ZXvndy1WxPRX0B8wOwyQgQEO/LLkh92pCZQ7qnHTZsBY22P8f0CjVWLDmvjKE2L9plhZ
I3YjgbLMhOQ6HwxU3HDZAJkhCWrm9jdteGPQVcximnF1TYT5ckZgvYxsQE5uLptk6Zjp649GDh5h
sOwg5Hx9FgjvbU+UYEhpx0HkPWk6GDTHDO7eev3cQVDgamNX0b2q2RR2ymdDktPgrDhSD0Autv3P
rwVCzUUdXc5d/klw3LapqvxnlrHK3DjhmyndmSdNZ5IUMxrwuIaLexrM4tI+ivNKfV4gwtnr19SJ
nvgf/uFElaXhgPmBOyA/9IiRw0DFDgt7jNtiQYSNPT+GL+alKHtuWTzKBF0s5YuuiOy2jkYrmODy
WyFn7AHQ7xMUtAwzug8q25MMpCj0uDs8TMMfVDpVZftlgs+vqaOKqk1K8/vonB0bhglmOteJPF1M
t4PY0HPHJZgsbaeEpSYNcTpJv828hQInBG6nnuWxPArEh24qR+3U7EZHSyWQ1jN0OeCdyGP2W4Qh
3cMdoat2kSMSPrXodzgnmno++A70nN0zTNq5V719PfHBHxd2mHPad/FXjeqM89PxnfpwO9QwXKFR
IWoNkM1cB/aKjTyi4vRhlNvoVFTXJnrMywmSxu1VOwwVHUXx9AUU3/jFP548/hzTe68ZEA7CPG2b
4/2alahWBSYrEx7bByGoule7mPFVATp95PcewXOrZntrIGr4fsN8JANe4+8wrW87Ru+6jndejxD6
svOrHyDoCB5dnky7psUw08VW2hH4Z5Ay1hYZcO8kx5sGmoTZm2qCJ+XrzkBbTwR5dGoZQbtdwxNy
j0jYGVUGBkO3sZvwhEPA2PjIXohZdsE46baxFBMxm0P/IXhocu6EOHMohAqpSAFZALTKWrLEnvY+
mlHgk4JU0sjNymL0B1T3S+VSxSpl8nTyHwfy+tWMKczdldWisCdHhPf6RRCQnKm8xrgQAwcilVSC
PdDdoypOZd8x86TEVBi9G8V1wvPjmSt3d4E5BAMT7Qs0qTjym0e0FOCFfNy8SBsNO8x/PL46gkYb
Npzjw3+lr3rH5w058viyIseQ1ima4Z55V8nCWerGfmiXFAcG/wn+x+PgVoQWSvG0mR1Tt5mLuzMt
AtQT+nEmvvDO0tOtIMXwbFwdClGi3yolw2vUKkjPvHQtwYLID3Q15fcTCbbTiKI7Dn6qP2Oj6BWY
31mHQarUd3tWj1PDRO7uEiVT/5ryBBimcYE3BICYGhDscWFHX5DCmQjql5mz0XnFg0IhhO+IvzgG
+mS0bX66n4GQZ+9zsb70GRksWmVz9lsJPzIYU1Oxp+cUpC80AUtrzD1l8w2mKYO0pdQ3Q1SovKlx
mQ4C2Sp2F8mtynghZs1cbdM7xLzZrYm4e349CTs/UERcj7At/k8caPznit122QKSyk7v4OHynfJu
Ffn6CoyQe3DF8Qxke9QVGOo7xbgw2Um2zeAnmh6bkkuwxBDhVGLQPLmDGZ/oa5XJgv2avyTFQAB7
qu1hzG1PJTAFE7EtSPjp65Ehx5qp4j9WmM8sCTBqDjFyG34X5z72nTatnBQm59zoCWQijGyjRMpg
4AIpMT2duUJM+71jnB13AiYYpwvRUCQ6JX2RAM8Oe6VRq9MfrL0BIfPiFVb/4JeNP6ZbJPRKv04X
rFwSveAgLcXHRnD9DDAtoE0ajMWRYv5MSkNFDPG8Qyy3oyNhLPe4gUAnhUS6qERdO6xALg5R7LPK
VB/NiW9d0BEGniZJ4yPUKoWLiKdUg1cx5DoRB2y0teieoxhdngbE3yMGs8zsyYhmRKPOCGegMKq8
p+jPfx7uJsw6BIzRMR4bMhxfq+t8gcCeWQoqsaZr9+QRMPK+zgfT6oXJojmUd2gySXAc2YdXtKID
969asNOKHnmDF1AvQS32Odlet7z2phSw9Uc7qbNJWejDibe3vBrun+862TTPFQ0cMA/HzjJ2lb7X
eP5Q1/G3ZEu9AKMnpu6Uzp6oqDyIUJjcYSFr2CNkEzu9K90ntWxp7GJC33fCdpcaYn9pRcW+BDi8
U/2DiU2Gg94sDaTb0NQEx1k8ELBKHIq+iXnHCOi8dRvaK+KLAs/kj6UjREtbqnXGktwWzwt2Mn5v
antXFHnJ1P//H+8f7BdU+RqfXKs7Il+iKjvx9Hb3fnl6Hr0du36Q6bx3pFDIbk/vMwJJk3v675Kd
04s2jdOEXLYYzWQemNDTGYOm6rO03zVq7n0mMtbWxwc2XVzKRwu4LQS2zoipTm7Q5tDOBsEM+hBm
mNM/1ZEtL8JBpwyoF3DT4BTy1Ho2d1JGndQXOmmsMKXmIn5wVXGnBf+p4MfyjCwR3qWndI83X9XO
mi7Gg6HXCFw080gIGbuvsUbz/i34kLkbM8m/F2cOdNwUYrzqy6lzUGKehTqRTuj3n77sLTm2khSA
q9/PAKHo8cyjPcyRiaeZpOb/KdQEJ+30ihdYnzHSF/7FDUqWhkZdtzlnuwBQ789L0z7YIywHtXC9
5Ur/v5GC+92KIMg/LIyGZ9TIva6gJfpYY8bemrTYjCX9OJJ72lmhwbPuvrNdTnxwf7Nf/+yTR1FW
FnRKD/EZlDexgnga8fDO1P4nvTn+Ti4tP45olWN7ynUAYVumjTw+i0NW9A5BbLx922kjpjBFE2DG
o0dOh1LTlBLP7cP9oa/dZ9BjwlS800jd5nw8AuDeZPLfQv7x5csQMAyzALcil5bzufKFT7VRisxM
vlGtoj/37NCsLw44IxmKlZlQiwDY3++sZPbygCDmpDVdqAwxPgpGbdFlJ/SeZCzsehicVi78qDQ0
dcIzwF5YZVegqitiCYhibKvXz3nWn/hXxP6Zx7HUlN2MA/wE+TcVFVHfntT947dkSvI7Bvf0NxsL
+GwKn95jt6tOwrQcFkYglCLThCSNqSIV7b1D9fT9rzoLGeCWbH2boGSgZziS5VaU0ty8M7mpedto
OSSWMv7lbCijonati6G1JRIBPNPaPEMjtkmL2kLANZKu0ZrX3XFswnT0cP6/YMcNvuTiiDgSzIjx
eJ1Aq0H4hMouDUIrbOOETt0ohstt+Y5M56HvU3S7KzjvocYdakMCcK70l7gDMhuE6oYR4lHfdUC0
WF4y0bP7bKbz1ulb7YwkWiHR/nryt2xu7cAPLDLO2haPqd3u1W7NTaH8xRemstLpTV1HnWbnhDFt
w2q1etHkUafGmB8+EjYN+9LXmMjUD4HSXLehfDuIax4pj34eTNreNyucXHhIyjNrvFSraU/D/PhP
Ra7vcpsqagTJ3fs5LyMTmo8cjGoL5Fjefhkzc0tUUvuwgryymFD93FM+sN77lRCK5WT8QlhESRfv
FueMHCC8NI+XdMmlU/pEkNkSTiLQ1MHBmZIGbFo6xlS5aJJfRK9qoGYRVV2ZepkrjR+day8jsNpV
qswn2QlFdPNRsziCDH2W3oWODBulLQT9Y8IVSIO4I0nZ9pCQH1vq/90DDvBNoKW1r7DaIea3aoMf
Wv3VGHwqDbFNXgYu2OYHaZZN7J7Y+DI7nkJG58lQHHHTdZFrfhAfcqX7G0X0dYWLFoNwHAQ3aI5W
juUNZlTKsliQ6niPwV47NFJW1ViDa3xfki2jtHMXKw8lNik/aNPIXarfF4XrqDBLeRq32/8Z0EZw
13SMU/YZyJ4AF/wJwbtSw3cmmZY1OXewrIfdRmGx4s8bSXM3m6ZC2mNYz53S2nFY1mqUsOVXmnUV
aGjhHZjr/q9FVSfZ0fLt8frBUloD8pIqC+7OaiB7LiRG38Pkh51nfQKEmq84khIJS3MTvxtdNz68
EM4dc/gOme+iepfbkiNS1q/oR0eKEjkZvdCk3sU3t83oWlj8420kQ7q3S9GlpdA9kGFemNFWgKpU
NYvw6wgsfstZTeFXvj+EA+p0CSb1VuV7aNeDASDM/e5nYLM3NG7Ny3NmMHd89GlivwW0yfRTDXcb
zlnQDJ3289ZYOvKYpjzM5lDe5tn+pV5Oy50M3ABCwMF+isuJ9o/XY0yAbcB/0M0HyHHiP+nEb52X
ywgDLCDWAucoT7INafuOar2WnYlZ17Dj9CsPigpIIv2QwJxoOihJh1uRykEdu8nIwWwlwALolytF
UZCCHJX059b59FLU9mMrxzEbMAitqemSexWwYCNDAZQmEFiYa02Ypo8jbrVfzZFDOJOgNsOuHbD4
L3QKp/3RCx4MtSqgEeSxkCYh/nl56mpHVlYR9lY1KdCO/xCA8ONhf7UmeyvwnySeRzzmftGnP55H
av2PJvuEL5kTyyQtzT56JZmDvhdZ/gaI1MCBjykAzvxOepZAcbdGHo/pOz1YlOH9Aprk5BMIfEf6
GFtZwInU0m0ul6J9LOcn7rEy7FLGCYlF8anOotiC0D+ZX7JBMqaEfrkhmQCK/LGJXwaQ5A/lwt6Y
C8/8VLNNdNiv6tZwboul8oWR8UKai0QKlOtm7TVx7PTKLkIdBNt/aRPfy91btTrBQmBuUN22fpno
y8kW5rE3dyu+2HW19RNF+WQIBuL93yx/o2H7qU2zpyVkQ7XBMzETw1t0j2KZAFRs0ffM/pI0kWM6
irwtCeG37gfwPXSdoLLiVXU8p6QNAeGVKkanJwlfeniCMtCwkcUCexHRVFiCPs202+BBjfRloEpl
2PmDOwl+gMJIRBOvKD2tH2tv7/4S1qe9WYxhpgdJQa6DO5zntZbquXL/yVg3jGe0S/+CUDBz2EVb
rggTKgIxnN2Dh6LoUEuRBuH70lH/4QfZONnb9Ntk+DeP07erTFeQlnoA0YD3rY5XsC9MJSov8jBN
Axq6/Umv+hjbHFtBJJ6Yjs5KuYanGhYELqMX0lZdm/c4/wU6tQWcc23uThmwZiu/jWqTLsD9fgQ+
RxSzxRdstwT8f8oBXo9JFQGobhhd+ZArEHkNEmOxd/JII8BAmjRuhjwfAUeptTosaPTJF7mP52Fw
uK84PtD1Cb5A8NJVVOEZNJoSdH25Bt6SIm56L9qu4HphazI5XgkJP+XH9hnFki+8e6AQxzIAuWco
kYCBnWYZ432ItMJ+s5R889tQsGvnL8DoQSiH23xY4fUZHvMUvyyhtC2GD5FOF89aLX11v6xFBrBc
Z5Z+kNtagWwsjq+7v+ABJwqGihMdC+Y7PjrfAenrTHqPphU63PqkAFbzt49em+I7CGd7J69QPAjF
2UuSthvx4d3i8cdpjdAuG71G7ltXRr8LUl4oN252OSqrhyrdjBL6fhvzkb97/Fa6zk7L2koKrOhc
PIgiz28ifWDEjz1yJlHkQfRhCOZe0dIBcx2YvHW0nUBhk2m06tHz20a9uq+YELHkdPajDRMxwApg
58Gza7eKESqdZNEp1mmPowV88WydhU45k7BFClFLWDm5tM7izxOVqUicwtx6yA8+XQyFhLqCJv+D
uUmYvHbHJrBnPu7PwjbrM+2tT5ibRTHK8vvTlcpIr19y0qKk6e74+fU/4ZhR7iGlJ/emXaUz38Dk
JscN8KYxEgyIt9I9bjoCxSEqfD72TkMhmIpmetfYF4a6+yfistCiqf7yJe4dEfht3sWODITyVetd
m35Mf92vuPzMFStObz2b67gMClkEaTqEQnmvDj6cI5SenJveSF87VyTjyWBXQ8rNZ9OHImXxWW7f
mINTO0MwJkoqkZgxSGzRm3r3myeyD0G27Qt5H1kOMD2oermIdkWrvhVFprpDwJ9BQOkywD4+KHrH
QmJcr3jZQqgxDaKdJzmB/C0ncH/qYw18cR56ozj+Xfqrnnz5pLy/MvFudvrqIrUVBj0bZbZK+dAH
roKMycsZ0ote2cCwjBu3wNbzpDNZjL/HPrH0P6k5kQEK4Ml7O4Y37O1bSCMA50gwGRN47ZGtmI7q
p8ZdgHjrVy/AiwC/tHxbY8IVM3CE77UWil5Wawgsjm+mth760ozogkyWd3mBmOSBEyBADUHfwNPR
5gicrTthE1lNj7uwRWknQcoOd5ogezejBNhhCPkv5KWBahmsOQBCWZJcGDtbXalIzINai70a7jyb
vQioQ15G0Wj6m1v79cYH4XKIsI04gJkW41pUYEp61fJsdxiIEfRrUkm7HaK5kwT8kwb7kgmS8zl0
kqXXsviUKDqURKxDUnLn6XOlsFZFVla2U7YNQPPREKBcOn9bDnysR5uZr3AQardgtsr9ggKMaiI9
srCKZnf/XBmamQTRJyIXM7SH6RSdbrA3m6+96O/F7iHHTUfV/Y1KoTBbxhSmmOURe0qwWBvf9Car
U/2z0sDBMbwGTZdPNl6fHA8M0XNxrXrNo9bRHmmZQTU1DeGPfSvsxS8r7VfjqmfJH86jjz/uyT8c
wmD5SFIH4fFvjJGfRbsPR6Zc9uN2rhZhxWMhXokBD3Iy/V4YQAOmlVrKxtUu9K4fAZkTu2ZyRoSR
fYYQweGYJIrsE+oELhU11JxzhQS1VwTgAw29q824KdBFzlvVlOuLo9kE+O1oVnpmd98Xe6GNMBNs
iZSj+2g6RJg9upeojT9DQI5/aljpigqG4Jbg8i1aBQM/tQt3UoJOncQinXVnubyXZgqtyET0SQ5S
HK4vx79BXjOTmYKQf+xJZCMgo2YWjtp0xdj9CRbaplssGLjjk8PZelA6hIxXga4EPQ3hL+u4UOBT
UI5mpOs+KGRYM/V0DGk9TzIC18+MQs7OahdpfRsBHRT/K3WdEXxeym43JusUqeLFB+gr6kctUze1
y52Uua2uKmhYYP7G3jhVu57f2coD0rM/R9umyKpseqJ/QLQUamDs2eLxUHDrxT2fxj5s1LKNBjEP
TKpQ2DP4H0/mccQiHUdZwKHKWgwa0W4fp2Q2fFyOGrZWxWlGsim+XQTZhNwN0XIc9prPdO3In3zl
Telml2mfljSW0kycrgw24yT2kPsFglWxdHJKEQZ1wAb5dm5S0k5iFyZhNaWt7qh2P8a6IJCqAnTn
dOxQv5/YPn7SEAh4ZR+34xnEajHj7Xf8jAqPHslHKoSne6spGhUId7jTqU38VwRFIMXcSTHUBOsW
XB7LsOHn+BraG1H7rkMlTVxLah4HpmaDy2axou9fDtjxVBSMkdMbnZL1PfdlG8zEPlq8nIY0UBJT
Hi5d6u13EJyqEQ5f61iEHHayjxBhfdBKbtjPtHVe7Uhs2QsgXKbk28d8Mz1sAZ1pmUjKlhVHgKFx
Giktx2RWkKZamIbrR2EuqrSH5qKKSV69zSXHxIrd+eXElIzCqq/wXShhy59qkf5oC1ytsUKr3QPS
MfJ1WqQQhejtD9Cv2rLh9IgPJgS8U9/zES4XP1gp4VWaOrMi7YbyEDFGJx49qaF9YwH9RCC5EQUP
kMH7Gaoa/+ICHb/Qr4JfUD+d3L2QpV7+KwhFv1jnChEcZQ42olEwVj770YAOxw6HKdqzNbHmyn4J
Jn1jrHXVoLknSX8wqFnVSRw7bs0/D8AUUTffLDcX+Lr+ox2JeMv5FhXZNwgUujAM1sLEoj2NMKS5
DadrYwLPNxcGyofoYTzGvSIQjPI4yYuRTcbheHa8D4u3TlwnW0BNy2eu+7jQGjPTp4wPWXQGDh09
E/jBXFA412d+leqUzH7X8yf5Q5OwOBtJlxS1kWl1IgdVjsTamAiokQLAEQi+6GcfHy9pFZ5XWXSW
9tm/rX9A8bM3Ma9onphsftHjOLSjakUPPDf2pTh6w9rRKZucKnd1Rv/kcFq+s/0mUNJZB39xuBLR
hco/vYKza9SuOgkLReMMnYlRsbqRuu9V8odGhVK64ELHUQ27x9rU5j48uoEYxr59KAOszPRY5j0i
NdGv1TXDfsI1CCbqfXk0vXNFZVfCGXBIwh+f0dkipZh1KZHwr8DkUozzi/2ok1/+xXXWlPcH+yd7
yeJic74QMLRH9CwYJMI8eZeW/4sCu7OZtmzjQP7xPVTWw68wgb7I1Nfnws8OCRjaLvkMXjzye305
6itjWTXO8xOwj/C/omEZ2/+cfqmpODQl6tGPGz6zsHSumPMVj923LJZziO9HBwSrGWoeeNsNOY1B
UnU2xP3GGdGAXSxjfldy3GLmwmmqD06trdI+yeoWXaCaNlhu5G/3bt8E3FXie39zsI4r9W+RBj1N
Gyn5A6z6+OzFumebbsu1y4ROI9gEcM6e+pCTdqgVmM24EWTyp+zHZC+NflNbYX35VC9pSBvpqcSH
tz0iO4mpCpwFpvu/HUxFoppgpD8S50qM+FTxPN2aciSrGvT52AOHKul5qiXn3TFNu5IHuokSbA7M
nLEjg8+gy4zIpYmN9sqS1CGa1nEHigyG7O2y/VKuazgGYT5mjn17aV8+pGkpdl4I1LWYDqSXsEZg
GT/QgytbeSJ4G7yU9bCjBA/34tjiwCo1IMsl1jr1YnEG2zU+3NEUrNrFkM9u0R2mXMDbJ5cY+Abg
uusw7Vw9nYaodEF+1Z69lOw1Swd+292KhUXLhXkXSlNTxtjxiJ2z5Rer7aa7igOTX9nghGNjuxXi
Wv66YidqZHgX5kg3Pg4TUi2gbVOfgml6Mu7s0x8ARRzKnfmG2lXtOMeHb+JRZVQoLU9N0W4w0TCn
JTJ45r4Mm7hVKH9YeOkOPCc4Ebtjb4qbw63cFsDdxt6IfSsnjxUwz1gEi3QhyKGFhc77jrh23g2y
d4pS2frpxQMjvK43CN8FOZ+PBC0CoWmHS9PgCXKvViC8Alpn7WWfEUm03dxdcXhcD1w4G4T+1i3G
eCRg2tqjbPkR6+xoJuQ6Atm02NsLLyAjPcBuKRKEECdTjMYFA75pOhqkFILlD3AiTiVMPaBNxZZl
e8WnKVouwWZCMmiMy6hols+IGm1MHkxsaoamcyqLQLkOrI6JmPjce27Cp1ua9yNtsorZBeUn+zaE
4u1ZD6fjF7N6YVikVpB9OQuQUz+oaw0rqxTacoGjrNAus1O40Hv4S31mBTOil3GqnuMwLMCgzlx7
3Vkq58IBaQyS2Ty3whA2I2msdMA1p1QOON6mJpRyhtT5wOlahulJ8QnAl597ujxQmRuJOGdJ9B/k
g2ydXfAPCLhlhLP1My/4JVJTn80/Dp3cqBPL7tFvJ6KljPiaK42Q43tnrgGtLEC9jhO9vQCDZK7t
tK1TFDCy7w0AAabnPmdasvuYv7b+Bo6X6cpT7Z+TF6M2G5vt/FJhLYVdE30x1IRlD2U3kIEFUxRr
5Qok9aJeL/E24vO0JufjbsrHWhnl1wDF9t09j0q7hr+I9R+4lSXd3FJZ/n2pSRBJeW6dopKMbQS6
lO4TDXs03BqF8Qa+60Tl8Alpvehf/KifGlI+sUReVXdz55NcrV+83AJ3nbTRTfDxvAf/2sIOFF1Y
wAzRv+NCzJs0yHAtv+P+82f9oMFtLrLfIb3N5ffzDAcqPCpwooWAhC+zaVd62yS1EiLBrPt/TcB4
HsXqjUc8uD26zcbwqI6v8fOKN88Tfn3M1fKn56PPF4fsKuKQqnpGj8wr8IZ/yFZef3WYvW6F4nSf
zFbzPecKcM2gcdsNU3f4dF9aRV35Kc2ZEb7udUtMRDxGuF/w9gaM8AZ/wXs8VhwPkBQlRgURLvXZ
TfJEbKlmuiqFD4QWCq00WF11+XR/Kq3aSYslhuQUuYzDbBME0FvC7v35NFJF/8w/9/fYh0CPP6H2
74v5T/MAe7ZOjQhRpMNz7+4+n+vIpZ2VCws7bEqZDz7gWcNg/XfRnQ4soGMm08U8qmK/eZs/OXC0
4OLG+OB+N3UTeaQ6d/OlSfTMo7Jbxk57d7aZucNNDpKcItticQ+3VBu0OHzsz24YPFILyc/2wsrw
tpLNbOL0wETC7klxlxO9QFa1eI+lcPcmxu6p2gLtPN0vFGlPibtF/QQ/BE2ruB1ESc1Ms8Xjg59i
cfjlcvxD5NrgZi/jjOUmRfr3RPk1Sn90kbEU7Knp9rW4qdVVif+WHwKMV3pl3zxxkoG0WXM+Eu5o
hkliWr2d2lAc5wY4+M67B+wxjE6kj66jEz/Crh/9GvKzpq2UxXKS40SL+HSHg2lmeODTMCUdAwsn
hq18D0+PLZo8mAYNvnQPhmKmVzWjiYaqEXCzHZ0OaWI1xldTCZ26NLPZE9M/5Gj99E0iWP2/C5l6
vNIDpYQuatxN7A0DaZeV2DGnmDNsdNnIUsVepigSK1LEtOS0SZq2dFlI16dMMwwddfASMFeUVloc
0zpZUd0ia5LnyLs4Rd2GwpPr50BBT27Qmvqg9dUR49fi/u+s0fwhlS7p+GACaJNg+IVZM+xIq+nZ
OwYPX0tw4hrqdUExi4m1QE6cYbkw/gu0q4sj+x6iKIHsazFQe57TgTZdh05Y5zab2kJsWqfppJMx
LzrJW+9i1baqYeutF6PFqR7gC+6qAIYDrX1WHPmYzRUuT0MphfaxxVF019DipTOJd8tmgJRD0sYO
fWGQsLYnNCkemk5jMzNZcmdS5AXpbUpJdqVnsXYsKN1YlrfCk6yM+hQ3MCrG2050FE4JRKs3w5wz
83t7EvwHdz7Z2gTnpgfwmCbB/TWl74+5o5ex8jS99G+2ugY7PhCSzffc+t/x90urKMphQfbGGnfk
hul6Y8xcCiFbdz27/JqFMSGoz4keMKZuAcIGXdYut6HrCNC22gDJusmwIJQke+H9Fo8ZETigk1g8
PX8CI1w7pGG7tErxtcH8sIbxrtSsa9BOAE/SXimwpRx/zbJ5pwZPuJFId6TZi/LK5OLnVfYuwtsb
uDK6gQessh75vxeNJsNubxVX1weicDwWIsaWmiaO5FXVW2B+yBKc+xP9OKwt7OuvRteyGXr/I1l1
RvmOrbQRLxpPeXRC4qGGtNQU0mK2j7qCS++Plfsbr2bf7t/x3cysWjB5ff4173TPbKqKtuxCxlti
MK7+KgpuwvMTAbN+RszQtVOIUZsSgJhxCMrb+lqqapUaCZhHGVxSGkrp7gjXpCwnpSlWkBJg9MtL
WO4JmBsRTfrVZQveplEdzIP4o3AbdLo/DLg26fRDWioRR415US4MSO5bkgdU8mf0fGQVKdrgGkdQ
ioEsYTH71B22GDtZEQbcWKTZp0JJbJCNxFX67oppDRCJPIR6MCuzQjbAMGlTokQe1qJEMWVTDggh
7o4KyzJ3a4ERNm3VCfDWDBbQD6VJAxEVOgF1qfYS0+cg0vnuTkgkKF0BvkLzYvE8aX0vRahYAKx9
z1oyjTBubhWAtpKwFWpalceXDYJZdmrpGVGL7rETyP4j+htn4aUmK2N1xx1+odY+pWcVsyJS+Zq0
bAzoyK4fxd+m2zfWUVmcj+b0cpUGTrsfzOzeF2PiV5HaxAdWsdPrG0Bd9BjL1dPPbKp9duHM4rx0
8kWtvXcrJBlWocb04PbHx0q7pqmI8A6GbscY8xhb6rFgOjVIR5e9LGChLahgbduVL4dnqXfk2Rz7
bRH0U9YedaJ5GHupCkua1weP/2+LtXZwUR97Q/gMTA6+xNBIHMg2azsTBNskeZR/g0YnKgxoxZ7f
3ntAz5yzSdijedmWn6QOJnlgKWB7DqMyK2oP/Gfh+VbR6mqxMGCnh2PDxR7ALE+0Eg8QYvl8Lr+c
8s42nGxLHrsYnnsNFDCNUtVUkTzpap6T+4KQkFZCKzsnm5gDjT0oc5CF0c9rU1g7M/B0jrDLPxTx
Xcb5wvbRbjkmDugd/RsA4zhGbXThl6hmnGs6sgCK2csNRAH7PHPRUuDSNL3orugS9/QJyzwvbDJ4
XyWBBqYH3TXO0iRxFpIOcSSYoKC11E75GQU7nXvBAg4U/0O7NflyKQvdLq5Ud0PYmWD0fL1VFqwc
7bjDZ1HtDlu0WZqLEncfxSqk+PoCGFa56lXSMj79g57HzTe4GNgCs1CkSmcsNMomrTRWmy59HJQe
dhqhfseZtJgJH8hd1pMmjSfrfUtp5GxD7FWFX3KkT0L+yZ6A8lJMHqyG7gqcr+2PueKZY9v7EIdh
EIlm6W+XLERbtN0zPz7hWGf/CtvHMb7pCkb3Zso+7+wqLykNYGIvsAT0PIVt6cPlb+Zs/70pxZ6t
gzSCazzbo72Fmbi+SfaCzCeESYIfGBMtcx+YMS4PZkrciEq4R+KQAb7G9qkthZUid4wc0fjuQl3S
XJ3cw3KTuh6gi8BKhsdBGfEhtl+2ByZwR8reHIyvnl2qwdDHKWINuzt6uegDy4rKQ6Mc4zMfeEw/
CztwMCLocEMEKMuGXY83oV432UcWw4Ek7HFGDcBJwCcOS/VARSt9AP1ZXclBshtuIcnrvpzjd2nm
8I5pc9yo4kpCK1d7bj9j+jLL1wtRYTXOERtNxskQBKWVwp2tPckTZbtSHKlKHL1mpewUvS42u4WK
woOfXXUTs2KUV6ZfFGJ+sk6S3sgETKGdxT3KTuhu1D+m1y9uoriOemiYSKsgCQDRlQkRlr11uTAr
8QVcU34PITplZijThuMBV3KcYW3dI1WoX3HF8FthM38L6yRktEkB/niQmeSPt4x9oPpKUTylF6Hs
YXt4WdUOvm2k8pBNB4j51diUgoodS4M9+ecO5UhOLgeLaPCGzWX5Z+Cyb/aI1Rcz9VnKL+PhKfwI
Z9NO8Sl45in8f7bHnQ6bfRyp9a58jMNE2IYJSf3r0oz3wJjUoMsO0d9KZMobOXA0xczZDdboHN95
hOf4ZTTXrQ2VFLHbWAcxHhWPLxl+ynKVRmKiisg3n7dWodmvXTa1Ulex97xc81vBpE7MMyr+R3OT
ZP9seWdbZQqGWypCxz6cBvr9rcgQcH+DU3neE5yTbanVfak6LW613imLWoimp5X7QtEmmtmAjXer
pbA5Vr513nTom+oTzAiWdlYkrNrGikaJzLYI0ekXbZ+mxCmXaM1ICEN8guTEA9XthwAjY1vF2I0X
r5iONaD687FXPFjhtZuWILdSwou5xy7Ms902PimexA8VzqGaj5qDGZVI2wjMl86+b5F3OEQcOzkY
cEv8CPAQbrxW9liEsIOfPFtony6VKkiTj+qBIxNoeWIENNQFzzjloA1XWvovvzq19NGDy7MaSImC
sAu3t7sa2RxUjKaD1o4PIiGyMNZYNJq4VMr859gjf32cVBSW/pxN78n6/VV1+jHpI2+x4b3aQEv8
XuhjLQ5bHt3GIDeBD31WVcq82kQYDrkYnNAybL9Lh7yDrYAwOjebiBmC1ldvWheAo8BsGBOtaIr+
02hbMZxLJkJYQqvDkcxEI1n/54v7V/TUvB/o5aD15dVLYT2ooZNBiWqFoBLCc7lnib4BJT6Ak5Ct
AtGLWhysE3kWirkhbe+bkSFtuRz96cDqIUWxzozuMsfA7RzRg6aZMXBj1vkN8MPY9ikWSvh0a9y1
wM4L1AObv2RGdbwU0s5MipGxuwWTrX7VaIj6RikRfmfa4cIzHtQlhkZWsacpVWzPYekiQIwLUHjF
12WcXesA1uNy5nnVl+0pQmWwuYe7SJbZhtB4pGvji3BJdP2atmEPfvE3C9TTQRwCzje/ZDl1Z8zN
2arRQHP3gTjdC7zUcUEnuue1oF6bojt4dlnQtJqli3g1yttei1UiGlRHe6eqKH1MDPdka7G1hVxf
HDftAJQF9yqUK3fnLDQX9Z81z5ecAe74RLK0Xt8pqbsvBZpGyQyRthqkKKSeEsmGhPsp/gyAOE7X
lhTaYTx8mj/x6Bdd0LstlDVY9HnjZogUKj9+kcqszI8QHvSNC2StK0GxsETRN1xX/LimI8xSBkeT
UveIrr+Wu6s0yHstnTkYI+i6VvUWJFSSe3EdvlF91G15xtIz5MSbMa58md6Y7i6pLm3UHi2bAQ7+
w9mQnwaXTXIdlbGAv9gk4vO53tGQFMUHWphBQedBZDbOAohWxzQxykdp5iqQ4jDcYPy12t2D8r8o
j/honF0um8T2MOTsEvjxrrnhIx4Kf4ZcQYaB0xTzYsdTl8g8tlrVvuQFucHrPKryyqsCMJaKACjL
jf6VO5gj2IJC+gCQ9lXnc5ZZkcjX1DjrCfuoJyzV3xgASLBY7nIDyVDYBRi7DAGdC5lKj1bihkZ0
tBz2QjkvYx/vStHA6pzvfl6dfTNAKieT0iYd7dsVfFUiUZsrBgpNnPxcU5RbmNJIuX5V/NThe+fm
mwXti+NevfYdLcR6mh17VVnxNf17pypA2ZovfCVV3LxjoeS0w00ZprOqdf4ShprCgUaGJ/vYBHVd
Il8d6lpSwkU0Y2XWXDUFkmDCrBfAexJfIjYs5Jqasi/sbplwK1/CO5HkrxHNBSKKkIWit9OGiM39
x6B16jfB8klT6gvEWgXWRyclNK2rnM88WpfDSqRmhN3YusvSMcM5/+zkUJESRHgJ1MCzIZZwgfay
Yidv83v0HAlVBERrl0V6ulE5sb3qo+7vMR7tGkRBgHOYX2kR6uc7TSPdu5CaCnlzk2dIAFGprQuh
iNpf2KAcHEU2WNsxxwjRUD8sCDHA4OcDUC67gzfk8ynaln+qreh1Pm6eON2icufbJbAJflgOcCNw
tDjetnv5dzKIcTGpUpu1d32wCCQM2N+d3eWAFltdiSgF1yidZzhBKkdBtb1Ela5rLJFH8xgE6nog
hxk/RiXcgYzXkagFevDaTqzNelQ/7d4ad1Wvecm3z+Q38VfIt8yceCvFl0YxuVCm0nijs+Vw8nM5
SiJchcyYkEBk7FUoOw29ljm58TAxWmf2ssR+L6JdCNjdPmHvOjQ1jl2/XjjsfVXRUInUyp9pgtdH
7Riq0OpGQiJVLtqglrSfA7JyCCKPCmC7cbSh8CpRVQgPSnR86zI+BqJPR0MfC8WG5xEeOGWbEG7a
ueLbMZ2wnd2tK4Cd87JsP2bEzqF17qwEKVIBXQENW/UCRus7QPFTh2oMOiPWgAUJjv+Jj+87hV3v
3dcwDLneY9ch8aiy/NxAkhGS6NgbQzLTSr9onPENi2wSETDwIV4wOGurH2G+ysYYpp4slkJe0mZ2
73eHZDg9QiTd9FWJ1OBQGD+C2VhbwGnlLoA3FjmhBcFXU0i+4JR+SyZOJChqjaoQnW5JO+ABrq5q
3hn8pIrc3itbQ94puuRZ0UJXBrxWVJ6wS/6+ERh8x347uQS6kyrLJ2mUFI7mF5tjrTOaEEZdwB6p
qQmEA3V2B0KIBrteXw8Glr7PnjFTBV+2ylSBxTkr26Nb0CwsaJotxsG+bXxQN9WCmdJEL9QTMhYw
i6QUC0ywnuRDaZ4MVpENx6YXcrhGvcX61a4vzrpNNQ7C7na3EbAVClTQXZKwpXTfogI1KGSBHpk6
iNp9d5Td1TTKwltZD4nhXloc5fnSgcGKloMrUAJMh2m4dMPw9eqy5FUAzHz+ELq5txBLw6sqATiE
rhj1ou8l7Ue5zIG7yxnkKaGjjVG3pczTSwH0p9Vq9LrrlAiuQFauWl0s+9NMzmn7yoXFSqle1i34
btRe5uYxwFGWY/kaBRCsMZP7wzMdvUftTFKgk9M0lWMZhCd9sUJO3Rv8RPqmmfmDkHZiyRkfthpr
Ohf83ryb/EkmLit+GHmELQq6GIRywiMOFlyHNu3UkOc8lfq2M5VmtA55r2uh2Vsj5PB0q1SYgizB
XwOwNFRSw/exeJJvFXIOmJtP2udjsJn+akumf62+bVG50CYiZZ0oMOW2ZyFO77rbsu/GE5laVUNK
/lxHBK3uYmDzO62UZCczWYy5OoTU2zyaIUvRxryF+U6cvx0kmiMHiiytK2ZW8FQ4oRMwFFC6gNzz
9naStF3nJVTjNXVUx31fE1VTwcam/IpCBN7D82JT3U/KbYU1ygpOQ6tBoFnafVoAPYxdw1lVJ0KD
S4QOjqOtT/BC0ZF5/PF3wHhVIII7oKrUsdRhmPAvQGHVTX614XCGM5EX6k/hrlj5V4dAgV06PP5N
yyPH3gB3aau+fR8k0qoqmtZuSdPAsZaxq74X6mYoxE5zyXAnj3kiWl8Lrhj5NyDundpRhxB2EzrR
BHaxVCMhA0cMPW9eQeWa+22nHqgOB3vL0ct4NYj2oKd8ZHcNIgmvOL43CbSHNcjmJcD//Qy/Pby7
ub9ij1uZYBVQakLMk669j7d0yohdTjO5tZM6p4znrd9Kx7MzxZeu3tiejnJ8A+HFjSl+9L6254dA
kYE9GmYsyBNA4dS/nEvctyRBM0JoPd1ij/6+4Qvqii8YveK74O6srva9Q++xF/6KB2jj67/KwOs4
inbid5dphcTOGK8aYh56uZwaM2BNYO8g3bmK7xImrIruOA09AHScTW2DbSNvnwaegoFOa2ufWcRr
8KpBH1SF6bB/+VwAdhQJQ4be9UNKyeCLx2FTOepIF1Y2cY3CzNdUOQcxCPNqUXcU7VHR4OHe9FSb
Lo/sZPhUYGjxjJbSAKIdc9SOCoYZ12lBts/OmlKMw3a+WX2dOtBo1Uj8rSE6Cd2Ov1GdrBydbU24
M/+iwAPzuXTvmskSO2iW2DSE+la8Z+zeWMrvanEjuzAUmrjEfv9HSD9KsnkIg7TSCPgVw0gDb6r0
i/5iIVkId/UA3wHtUHgWd+wnbQ0weKmxWRGpIcIT5XdwRK7BkaQKvyV8+xZU3R/n//mea8JpDMWI
FLwY1TEbl4709FVi+b5lF4aCT5Speyr5oVZ+zVpK5YZHDei2KJC2BPnm/jmlXx2ATvsoCcf7JQAa
ruF0uYR+jNLR4cJ/gXIyWyROTvETW3biDWT2bza4fhEvizwJ5FNzQk/aMclZTvNuSEg9YxkbQLol
7UOzkBlX2iBueUSPyCRbgGg5l0xmxNLuzC9PRE9Oulgc+nkPo0KXCwRekHJcfbSZqMR3bnn6ShHS
RGmSBV2a3cDkI6rbtDjuep5TTUIKig6WBhiYKuILsncKzxj6jvU1j+Viji80lOTdromWgYGoBXNW
/0WHj/uZwA7giQq720dCRrvMbmkghzaKEZIx8RWbArVtCEomotcjVycjJ6gTs15/7vZnln6yaz6o
8nk1VkWazDSS+sAsg5NwTx+OUm5FoGEu9FIR3eut0F7snhP9wrfAi28ytrRgZ8x3pCTvuLjBYuR6
Wa5c0wrXolR/b8uSeox7O23HepAQuVeoLQTrqXpSUb78lvKsq/T/kXEvpRypqWIeZvc24lapyt7N
Lto3kb5f2uzJLZlgjzLrdMZuuTDPv1SUf7DMPNojg6kYZP0M07V6AD61b7t3NL8jbAj9Un4H4rvR
yagtd/+0GrnAYKJTTbd4Qhk+VWWeqE7t86vwjA8L3E5H13Sf8VhVkjMYXfe4zB+ysITtjovbIVtt
+oDNNIl5CPaWfltlFgnrWr7WqtjevwRKOGMyWz5h/TVUcLs0jhvuCvggZqGWKZAjpzOTB5UpFXJC
JCiC40iABwKp6B0lKjDI9oNfNUL0VAnZhjGuTQ9rvD0gmJPv1kupU0jyBGEwlAedQDhZUEfAZIue
9St4xwO4P9znzJ2hlv8tky48VJ9uyhN5LPZtb87sQN78KfahAGhF+3mF0/5wSdr8Nu4u5HpUTwv8
0HXlPq5Km9EjL7I55PxvN/v3pRnHqe0UPAotswvDZntRY1t4qaDV7AW5vnhwmjOwUXDLxa+Rtz8T
5GqY+cfK0JcejUrE9UlUfWCJv7Pgu5cFyStJCEkcM+iSKIEMcSf13My7aXU4QGy6jVVwBFs4f1ZJ
CLNK6ALaN5Ii9oGMt1QwU3hjhivUoUSIkPYEU7oFATQPCJon1+Ssaxp4h8GyLI3TbVgicWvj4CfL
Xn7LbIMNvyZNPZBuZugy8imMk4W5PPZnWC7kf1qQtpziQe1V0JLVddoyeJ7tgUv7rQVse1rgCvqI
Tea0knj6/siWpSnSHLDaFH3H93lGWtjCll3qy/wKXU205ywOlour1ZvCv9RVR2C2NW161nWyutVB
AJ35/DmKki6Nu4PBkJmEx+FB8DLuEW4JIkvvUG3vWf1/fZWV093Tu9nyji4JRsjvAouPURy0aX3C
G50qhMHU6HWsbJ4Jaro2YVo3rBkdtwWoYgb7VkfgtzKDHGrCF7KGHlBtx65m/PL9USgMgiiohYZO
vb60+YjXgKEigBNKtX2gXAwt+msJoPX5quUiXwT2nrhGfrdcNymPL6pFryNIWGkJ00E7bd1v3A0b
yBt+838c6EVcgnE9WNgAjIfEiMWjB9FIZ/q8M6IBwqgx3/m4XUm5HKnGcEPgduo10fctxut6+H9D
u1RlXhvXQz4AGMWZR+sTsK8eMiDB0HOT9D1JShlCOG4qoOod6ehujf1MSRDU4YZmi9t39RBHHBZu
LgNcC/s7iXsFBdXl0SGSY17dsuEgrAszxtjt/OW8/Nm5OfefsZ/nmtmRx1leTqC7fQMmBYJ0rLGt
eLzd6NSLqAPkjJ/Dplk+hQoXx+qYrXDRHirj6jVVMv/jIvx8/Ks6QGi/BrJjwH5OYcMQvg85DQEE
ZDNAV5j/FYOhTFZzrP9IFIhG1+cLa2WGnb5NYL5kz4bq+Ja5ihDMGGZq3/MAMuluN0uheKE+POaa
9Pub06EXww0vyfWookv+80baO9QqVnjdhhlieGIP+XYvtb+QuHxt4m/dJTH1WOwO4tmqI/5zYngk
n5wIkaUz+ekUHoGrVrw7vdPx6B+TZfi98KJp7whpOt9mRJWuCsj9njqfMyyGc588vsCaFRSknYD+
pu9O97Xy+Lei/kW2PmqXVznAQuwrMklWR7EYW5L6FwHwWTMlKZQTe9XMzekrQ3Hrj/1iB/nSjf1/
zhBzprDpv3683+Z2a4rXLHyRL5Lh9jajSGX2SLTxo+EGKMBzYQe+KqmjpsKqLVKCYPpw48FyuQRD
LnSynhg3rgZp+Oq35USi1e5+MlSRikADZgQpEIZfIZFNJ9PuoekXPE+fX/d8tB5KtqlU8BGwh2au
RK2ZdqkyStJwDPlXEfFNl09IYjqE88qVcmryqxwrDNEOyZrV6PhDnBRSB60puCRcT/jq9lyYjt2W
0xvlA4cGRuvWgHDrpgJQ+Ti7GO/BCTpmcX02wzFwyp8gu+7dWwU4agVOYoaJmnYCt/fbcvDtBNQm
avCCMFSenNd820//8Pom639QdI/UZre8BPWH/fKG6wlyq3ClDn7AKxUZe8Mly0f9QExWyyXjJvXt
AQqn4zsX7VPJ9CeZlpxBlOvmnFgW9/RyHWRMtVS+svgdU3c7hXddf0OJa2pL1qZvbJD0tQXSs+EC
Vft4m6HrQ1ruI6DQdZKaeB33YADr1tM0cSHN+2GXLAL4P5KQ+1638FcFfXAH/Eg/zjF0vogV+Nzn
/M4/v2+dj/I2z25sh+PqyDJ9eKitf9KJAUh1QOQgP+KfOVp3uWaVKVuvccuor54hCPX4OVppk0hj
rhdcY5iVq5l2jaAHJASE75DIQBN5HYquu0rQgsZPfvB00dJ3VH0xNyhVX51y4N9juC2Qe1rVkbtm
W3Sm/599cDSQ55nmm9KwJ21dZ/6vxu+P+38Od/eFsuD8pwFKbsZPbQdIuU8Xp9VfqLqJZ/K0+gyh
YyfrKjpNsFNUt0NUoQ+5RgXWrgC6odcx2R/nCZP4EhA+76zm+jxDmLXhBjmNqC8pJ67Bfdo97IWr
nTrZeEQNbcFp9cyF0tpXfjPNNyAIN5RtjJ4JgHkeTju5RQHqhzOicvGpl9Ys0A8iX8i7CyJD4Ae5
yo5JAtE1kxzdp4I3FmTa5x9AGfVKJLyIMUiYIDBVoLlr02LorlG+iSbZOJLRkNxffGTakWP4tKsC
1+J1qRQ8LerOEgziu0aWUUJp7xxj07af51rcAy2uzhYmhEExcXMQF1JouYwsYsT1yHs75IPwUu4y
lsdNqgP2+2FRDte5ep5zTk/crmibuHuaPGye3+LjXXYe8vtPAWG1HW+WB4iU14GCc6qHAr8Cj08s
WMxPonrLK7+H2sI6nPyxpGTNF4zSl+xLd8dZ70atA8jWBvGjcELFcCe1IxLNEXCv/o1y9qwgkUNs
fGoJEBHalPc7EeXA21IakkbVlpin65JHB4s6xO8VRLimXx5kEzhzsnkSjlKWi9w1e1SMIZMsaBRJ
JM1s3GgF5TeZ62BL6yRnDBgt2JQNGo41BDeXQ+/ySDQPsk8E8MzLI37yb/L9h8H0dRCYQvcsGy+w
d/L89U+Aeejldz6OkVFP+GqH9KrddAmWXF7NecuVepIMHXKgT2h1wDXVjbw5pnHsbjXmo416Xw4o
2uFpUyOos/q0E70H4MHCfcCNHcy2bopHbgmhvN207ieLyAuOKNrl9kb3txEsHOk6wDu+hjqsOw08
Yadwtwrh9j96et4x5n/0QtryJPqJRGIbdOzUy5F4fDpCERRi+eAxs9F+ddlwxNPpzV2Y+0NBV0/A
6Xrouf0aoWK7pqNJo1E3sfJ5IsDmYkEhZ23/Aj38fWHlqL667V5dW0hPzX3rVZ4hdK9/7iZBW4sy
X5+Kq/qw0ykX/37lO6tgpccaqimIPyLy+XKCmyVyzKgoqgwcfIXDAemj1AXRy7kDkkXbQ+A8ohnQ
pxkjwmsCOwwggEKqQadR8TTaiuvSNSiTDTmi6uaWfuVPFBvqnBzM5cTJKCzZwR7SKYei5QTHEC0N
UgMgwNoxsE2j0gGHY4TSRe4VyTpMxVPAmOL5ukXxONChPRFi4N3zGX1O12SjlmjoQUOCLtpHQheC
p/jBNY7UGOQA9CQseHb86GpEq3KChM+450+Ob+kVTM6pKrykEIEosGhDIOKiCA41cYlzOmVG4drG
6JSUAC8Y8NSthWcDrODpkrC0A4TbDsJuzqxm2SyiXEjApZKdOjpHVIzhXOQCi6WlJ4L7TZyHXuBI
BR9AqVaQcMu4pVEg4jqAkEl3mm2EenL5QUNHodYm6s1ipkPocn2EwROQ9qEkOeyhUVV0ojptirgK
LzCzQmqrr7jRhAphssZ0AiMZOaVpoGieFxN35zZh1fLPAHvsl78IFlPQbkAcHdgncXLVYZ6+mohi
IIU3b+KWtf8D+y1qK2suWa4plyVV+/mCil5dB1QvuLaXy83dz/T6J7LL6lYalIbqbR2/sfg/tTWx
UGDbML3jKTske6uhJy0mBVjHmjhY5RfqXyl/Z4SgpCeLC4G4GJU/dD34ZB5eO1cvs88R7M6lUqmJ
DtDvRhpRxPwMIDGQUERM8HK4VJQiPWGUax9Fv+4eSROd4YWFdSUV2OLFMjHry1JZvYQTAaNxo4rm
i8ogye9x6maweZtmXtNhqn1wyIY3dCQTRCWC0Q8zpitXbVBKIXSxq03/5fS+Y/8BaQLVJgm+zzzj
jKdxv0IZ2H2GuNPxwEHPeHUmY1R+OUxmWaAlX7PmUmyjK4MBi5T1lBS4mZDcJIriD070Vo1YTFaR
ABOolhhEpmH2kzmA3rFWWbw6MgPYLH2UhtV28knVqnrWCsWPRmqUuc8Nz3OX8xpJWhWxNQNrxo2k
v+wb1KrUDHKYwH13zFCxu55KVrBN/WZwmE+SXviDQ47N+lqe3lxKU6vPyrq0OwKSEhD6khsiTgSq
4MwVkM8QlqcNnpZ8sKnoT5eEyBR89Rx+8ZSVMYmjoU1RvP5YSpoWjGixsNkuTiMIaKlySjPZ9hXb
wwA8rzXhJCPoM9H1MfY/U4amOZO+iQcdKnayTKLwoobq9sNJ2WR009VsRJl0MG+Zzl/rFFWu8BGs
m5Wd1lpkO4sQsmZqDP/Cqs3bgVVSMv+ew8gWz9NGscnLyWyhbXoojQceVj27ZPJMhY+6S9u8qitj
bWvfECw65v/XrlEL9xYp8kCxNs1oi3E/pZiNYS2m5SYviAabjQSEmCfe3UjmM7m9vOVK3OBNES5Z
YZp6W2W5PVlSCzVvHgt0QjEtWbRd7vTcBxnw9pv6r/24b4er87N+O1z+vo5h2UKiFgnKFGBqySDq
E4zQ+pWXx5g/CLd6oJc9bHFfp4OJKczH+nbw4yK/1PWQ74RWGr3c7NZwitECHmCUDVDkk4HiM/VH
ts6wzmsqStrLVHZ3IAXw4BIkqb6oat6Ag2BjBR2bdrB5ofphb+EGhLMXdjlLOOpJhjqWsDN24qj4
FfcKwNOf2pdChGj5abeFLqeMmm39KgmIxgSEEMxZOxN2JqA0uQW6H2pAHgEr1KakvKSDdf/cooWE
xsE+R6czCAm0GFZGBhRQeWXm2R1bFL/PaNinvanM0nOO+dXEQd2356gvY1El+k1aGwkLUkh+e8Yk
zihpwzDzO1Ls7lPsAo/N1ffyvwJ66Dj3BX/aWoPJEtVKVgc3kdJGMidmTeqb0lOUanbHtpEUenNR
ssKW+KbtFCDIwO4snY+J7MbuOOGwMKI3iutXHeToVFJ3KcUb/YsQmn7dMyO+jB/nrZNsCBoLzcw4
JngQeMMSjkFisOCbLdiBvkEDCDSESl3zR9+jv6P3IxSRTlapt4fHkyaa6Jbrpf58R9GbUvel/TSu
lAmwC/zKiF9U5CLxhRU9vY4sNie2VSur3R7qBAuL3zVvENiRlvNhxepCxQxRc4VP+w9yMavlxKMu
Hzwk4ZqSgMaIee50d2P+0H38mKvKRSa4cMzT1G8ObNeOxoyWK2cxvYBxu6rsfjtuBsxdNn2hwE+u
x8O7dcvwqHtTih4nK0vECcCUfShT1zgA7B1XLPRzwvGkIUXZP4Zf420YY+JqvPvGWfi5UlceSbMO
6/PiqIcJbQJQ71zWVnfDy5Ff3Kd6XID02pVYruCWjqJk2PJX71Ka0nOXhpWkNvZspr+H53+BfDC5
/73+IPIfLiq525yCo1iwdBdkLO7DobsWwyOyfdtbOS6NEuxBvTuA48o82TiluSVHtBgIX8KIHPGg
amFZJrj78laTibdEhCHabx/GLh110KK+bYiBsaByop8xsPDPqbJYl3zynLvDirNdlvN6b58vMFsv
7jr68I1ZXOwGIsczB4mNmOBpumJMlC9slB7TZS+02hvDNTfWKSH1vf6hHfXe4aZXk7l+D2cnA1zH
b4yy2FB1awK0dWhiOdxPHFJFiKlN1dueBuI5c81eQNCasPbH009AY3szPpDv0kykY6LIGHBtxPt6
kLUXbJHVwT1Nn+Xxsksumtiaws9nK0a2uCij46rkO6q1H6nYB+ZDcIiihHghwafrjLOU4tLxjQQw
HqGx+z4uJPqabZmpQKnqfJm5sMje4FXrgM0u2fHrBsEYXHDrrdGflmMkyPtZo//qcS66L/EOeucX
1caDsleir7k9uK9R44fTyZkcP2l9O+34T1Asx3XiEBz+AA8OeKbsXgtRfX12cN9pp5xnA2z+GMUZ
3LLkmO6GnsZoApme8ZFkYrwZnNBMXlqEe4tpqN0KWMHGRwxSJZAOxnGyBfTl4ZizORyaJYor68mm
9vktCOc0UufsaAc0vqtZlSI7tHkG3PIoKojODN6hnsHwTvB0/OfU6kG7JKtxg7cBfgQfvU9ttfoz
g0xBP8UqWECPn5mv+rbjANcw11uX5yqZd7wBzW8G4RGIecMqTXCiEUk/3hFbPNrm5kjEgk3v7/m5
Mt4hCQINT1bsK5tsI+t5jwyjXtVsIbD6v3pW/lh41wM1Kqt8itU9zmciukKodgKa8erT9TI+mrxE
SJKy8958+eF3oqB3yn28+zcb+m/IyhYs1o0najOTU52sTiB+AkZpp6yJfD9yEl+8esrg8VOuhj3q
G/PAPKk85crwOBtRa3zbjnmVb7slYuNOZK4vcbTO1sYnJWj5FrANS6tnhj0TqYk7dNyKCatHCxkg
Q4fjMiXzL+Zv+iy2K3vbCX84iq+H1aru4CjhQx6vtqp0qcNM0Z1m439ApqDtk05lWuQ3HmQoj5m6
aM5EXJvQynYJ6QjA+tvzNtIHHfMnBfrdTNwCB0TNW3KtTaEoWV6vf7XuHtIlq1bgoytvqTIK96nh
UJMVuelkPmohNDDOqV5UpWLq63t9+kFtjHQT+lE7iCxDHGFhguzNCKZ+kiw+zRTGOGOsdiHSm978
bz8J6uieogDvTyPieaRbUvN3Uj1jzzjUTWndyUcWy+aQklRxNLfdqpLjSi8kgjj0GeeuN6kQLaw7
8g0M4+R7sp8lyfodqbH/ey4CYCuRVTR1DJbwajwGfTdp2dhnwO1nVgmGyeM9Q9BeLW2M9RPCqtiH
LD5GfyG9r2EehTW0TeU6RMgiTD1N92ZI42krLvgURR8ILQrz6G+k3lDOgxpjnjaOvGx5mkVMwgDx
ah9+vltpHDjSVhF88yeFm9kbBdHuuzRv2M5bo7bCWGSvjJdafrIHrBlqeWULIoPtC3Ek7WqXkQkf
NSdJTRvfYsOwn1Vun7f0euX36p97/Nlj5WyD7ES3IpEICiXCM/yQJlXU+MuWNIEjnUhFe+v+DjyB
taIolO9H3RR0jBDhrwnmIWhmyPR5VxMX4nlBQMduLlMEakrGY91l20p5pgJXLMQn7UZQbUc4K59F
0KogfzPzFG9lSdNlMeEVidO5bTjM3V/ZpU/E867JTk6ZFsm++uny5CZZTlkgy95388j/29ODszzs
itTLGnLtl6lXXE/4B+r8PoPOTvVsDZ/7WIPoD8Ar74xEq+qEDCW4VUWfXEO93vFL9ZDBN5wJm3m+
eu6Yzfw4q0jMlb719d2xXHORtdcA0Gnfx/lKZKHnPDz5x24Ojvz2rYxfUsbY2S6lHMSricgP6SgU
36jd5oKG12q50tZtF2yBvE/djVifAEnEWA4Rfdx+c+2EPXKJ3FV8za8UWr3665RbnPpQqYler8iH
LEjOB66iGVdhWm7YDJPfQAvh3UqTIOv2yivPEok3JFdm/rm0s3YRzom8mGLqL7gvOQjwC6Xz/dvT
E0Wtf7pL7HuTlitk2wqdNbmXPjsp11dBEfYPZgvegIS/U5J3X1Wam8u+RVeSq5kv/q/o0A5F8jP6
lUDmvpgwWTUSL/ceXicZ/vMHeVGC4nV0iezjx4TkxZd5GjctNju/HolWmIA0ygnHeOO+VdniMnRs
YVtWb4AlE37Cipiplqxbdm2WsehAedhEkUwAZeD2gc9HnpZNhuiCn7MaNzjwErrpYOF0gy3cgOWD
MXhkyvcqhs17SHnO+cwXWUwwGssJhAeaBv8RrXz4V/usXBVMwSciY1ni9njbYZGraiAn0onsGZbS
3HSzYoXBu9/swH6RUdcGKaB63p77dd146X9Inq1drRW1piksAVyRslSEnNleSy5pdcfygibyrBQj
hBKOdlceOfXNpQ4r/kBKv2P5qa1G6QhrWUAeuDVeLdyycuc/kPJqlxET75cKpNq/bMMm0M5+j/e9
eTlBHx5BXJbyrPO5wa01LnZorz9kuWp54K5Uva9NWfEhF9PNInqvk/SFpFdO7r1koFtW+sk4rI7X
xKCVMT9DBuWPrrZ9u6rt2lxX/51tHM+iCiL5VvK/4ZUkSCW4Pe/919fizVJhw4aZS1Lfy7REsTHc
WmV/rFgCJxZWakVbC1/OmpjGhN3HI9yCL2VtzQvxILvwuh3FGYlaPiGMA8QPTiLQLZ0pPyB/hXbD
8nHGKkCZWNYoQ813x7/SA2rAMk5W/uSNfzJOtIMIOJfqYd16hwU5zMk6XaOPJtA/18L8r0JbOtqm
gZMqjcJPn/7wT975rxckoclFzZPf8S8p89zgHvQnY5eWa5HX2xhBiM+lNt6IYBFoCYBy2l0AOshC
SsbEfrqmHJpWvHFjmsYNR/B/3rMrL21kQcygGI5WluAjLifmF0eDKRgttDxCRZ9PRO/gkl6SAmTg
HfaoxLdDMJYYvB6OLT9TXg5oy0BaRBqVQcxhGlJJUgVHRjWwL1ycOUUJr6NnANoqbAwIoBMfbfmM
phDkVQj5oIreScxt+A8MwDvalTCnZRfi5gPkF2Bwr4ADF5iMYk5vYpPhbN7Dfd7MqcuoL8wBrux0
gRAHKcBwZ2bXx0gm29Zq1P2Soaggyjjy2SukuRWGWugJs3ZYK+PyxRZyv42tZPQB+mvKwmXlLrfa
FL79ZEHs8rF5YrHLyLB1/CEwVBmW/IkffcMUbaDErMJ1dZ/fI33x4c5SZwIyXK/ZwPDFxrm7oe0i
zD1k/V3cD+4tzB8zUiNQnV0AEX7bh4sjm2NLr6eypk2nQ0k6TSYMjlzYKO6ttCohlmOwyXWly+Xw
UxdC9I2mwBBKpLkovNig3ydKMuBCpJw9HpkCqpzl4YmkkQbepf2Onp+xxDy6xlaDXBpgqEPU5w4b
exADpr5Y1vgQYEkMXiZLpEof81gWRrgdo0l8qcibT41zyvVO/qKILj4YhZLeq8TTD1tG0xmSDe++
jRFYCAfAYqL+acUh6LROA0RjBHtMdmuzrn8iygLBvfCXv/uIXcu/A4XfuKNT9i4m51K9bYrXX9ie
b/v5vhtF0AJkT1G0/pMtHJmDQdPAgN5Ijv6W1foxk5pLdzugNgz8wLyP1UVhXX9tXEqSRmQggix7
rvVKZOrI930e02tDniy2DsB4DrTakrXL0VF5f50cR0BovVXvLjgHkGa2EwSaAdIUOngzc+SamTv1
olMapJjGoB4+spr7vYDXS2xGaCy8nfGj1VNoRuBXP6N1VFGYQPpGwbmNh2/CsHCGrvNop+9k1h3g
/jtVnWLfnXTcST8R/hAQL6sl8PRcQLnSDFAfnuwFv245Zp79H9wAyaUSLSZQ4moXsnFlVdzKrFg2
Y/32sSX7dmsLheztEX0fC2PRw6qZsbaxXv9I7/x3WFqcj44blkEx43N0LBG1eSOUPXXP1LILNqoQ
HReK+TTG50bMqSQO2Vhb1/N5yAmVszCjksqV7hsQ0IfdbkNzOfG3ro8mw1gNytLhaQ/Gp8Rodme4
ifUnDoSyQXJKJ7DH+GENM9dhZjGY/J/ehT1TDWWOndjjWCo1PSUKvqn3Vou1y+ytq+NuswGei76U
9Yn8GwrgHDBnTc4+pCd6O+AITzwjzCsR/Uyw6bFCycNiyg3+oZIEO4IYN5qimjxuPGS9kc2+q9Ta
l5fBwchVUxya06OJ836bgMKlC0JVt4cqJJB+oz/VTZZyUb9FakU6yrrYr2Wi3kkm4qNQWZ836m48
QZS7JO3R+fNz1WHaWhOk/ynszVCZooyB3q+zQh/sFVM4vnmeHPmddYKTNd6ri3HySTbJxjYl5Bc/
ROqgl79ZMoKrrbrc3Z6NZBCRsR4dJGOcrwQ0wk0stRRtyu0zhpmsrTRYGMOnwywv1v69fPkVSDBG
hAuh5acjAtJbBSzhNPPkWjnDImUvakg8rqqWyAmurCqcrk++E/L57jk1UrIwZuphwwqfeLgB7PR9
3Yn8/CSkN5epPRoMNcSyDWMAyQSdBeByCMKpKFya0PyvRtxXYGsd9QqG6/oG4n9bg2eyB7wYf/Gu
v//cWyBi/mEDL5W6U58ppOG16BVjututbiPnI25Qou4mPDoSldrkQwr9KD/puKNaoBLZLlU5YQ8B
xpz+Eiyf3V/E3rtfusuoIAlLZ/Vl3kULwIKVmBeVJLLh5y/bxS/gI8iUpekpSFB2XF/ZhVXh9AFn
W0JPKtD8QKWrpQykV+3u+CJcnZnQwh7/RdDLEN0mhv/W6V4EiOBMTt5eHDN4uAtb+PvJ5qFgYhkj
oUnR4kcNbkOZ+gk7lik0EzjH3SrzNgO8W56chZJ/kPBq7ixGXrrN3Be2XL6oe5vNGcnpL188SBT7
/E3KX1hsKNLvE+rWjJJ2ewYDBmA9BNarPHNZtD9YNaEF8VrCJbvVFuEZUu20ks89cBWdTynfqqSI
/Dw+74dQbXhuYN3DmpfRJnoUweFZmbQujt6LJ/bLSTTWOaYwWP7FNdIko0a5C+f7bPASb06ZGjwv
7/WHGzYri41x9pMh0+1wBBysqoZcA8vRJdzXmGCfO+v12EogLc2IFlSlT2Dy8Yz3lnbyPM/mE6nV
G4mpeIjfL79lflBSul3S2s7x1tbHsjwH6vMNViTOK5ev0gTHO5eUgSJijCU1cHe0Pa2QNCcCH4Ra
lsq6nJ3YF3z2Z71+yZBSwuDmy0slWwzmC3ZFVX+Vw4QQAGs4FyR2rcknxrzukqo2xT/kXFuRiTuD
CBtH+YIKgHoj9/8RNeIKcD6vuHFr6RuGO2U+nJ39UpHq6zL3Z1vIKGg2TLyYWOmW2vqrap5UgcSg
I1hNFAAJdiIt8gNsTW2rx8J1C18lsCCT7wpi4+2vp9SsqYFYJCz4gNomfHBPYBZO6mM0Bo4vUZC6
Po3R2nLUhNzFaOhEOORuKGDtD4V+q/8hXstck83D9h4AII9irjVjNWd+bBclgGBkgCbsdnak5D4n
riySGGh0wD2F/1wPZEMlo7BPk/97h5V2QoF/Gq97nWqmZ0zLFlMlKHyrojRrFftsne3H74RqSzUM
MYYUfIJexAA1wyND8q003zH9Q3406FWtBQTEzQaES1SOGdcXjlalJER7DklNCj/5/X+UvSRxvyg1
zoUAxT5aWuxd6zqRBZukSff6RoqSaPwH0raCx5OtxL72EihNtrzSb0m4svEmNFThzeRgebycz1nB
KG3G1SeSwNFYs8DqAJEJd1snjHUAAmH75rbXcZiHUuBsI5PDjbg9JZmvjTSVRBeEAw1dxOKD8OtM
Nm3yvTFli57GdTlbCYzhOnj3xvzokvFf7lPr8RZlBklItO4/UnRm6xOO39YxJxdpZo9t7q23LbU3
pdtr+L1CB1AT2WnYlaEm7k/R/uES3elV+qPU9RpHbivXYcbK0ZrBYRBHQqILlsydHfxIBavU7hbU
BspoQdRew3YJXikXA3TshS+x6dHjeo1F4R40itst1rYPU88twdOEYTWduzn1nFSNYEf89FGMnTyW
9YyZkFebRR8qIIXmk/qZbXhUU4gC06q+DvT2jPbVEqmTZviMt1Z2YiHoztMUTTEB9YIwBlN6YBDS
KMSJmXlxiubeMhh2slrm4fXNchZKCIA51C94JVhfCBpuRc53CT5M0dBvqw23dhsgHyevNikLo+Jh
dsDfirm/Je1PSrJEaYwQLQb2Y6qlGM84A37W3yZlas61UnblvONi6sfd5LVDDpwWaP6QMHuoqmVI
738XCAFZwlbxAB1Or/2TUPSg0d1EvkQjNrszMCCGK6KamsRdoeHwRF3reaeratqYffHFPcG7i6lp
8fGGmjDUbjXq2u9/M2d/Ny892jexhbu48E+4UP9ZE+Dmv9UQfQgiQDI7JolL6rEPh+fWAQNNaq+G
kEZLs/34r6PTE7/qQupfJqpaEpLGbAoBVG+G48axeAU6GrMUyopjXjW3YE8jaQ8Pi52JdIZGtuoX
qwy5V9p2EqoIFbcJ7wIaXi6LDXn2Nkvj3L9FR9FZEYfIDMdcqXEpmB7h2C6KkVBc+dlrsGaBeiCA
jGbTbBXE/hnksd1AWD2hVBFLw6A5F5Hdaeoh6xGpUzeBKf5XmXzSgs3Dv1OYAf619ngCzR0lMeGI
8kbNrSdWGV+2iXKHMMISopaN9zsFCQhx0cj3Bf3f0cEs7pgfkevPGcZv0WIU/QqKSWcVj6Wps+wC
WDZWYTVH9SCe7UqtefL2LPE6wswYpF3aLAr5+SgBstyHMZDLFk9Pdq10Z8TFgi5A72kybNEXtPcR
WWF/71FDz+bkxVu6OGMWr3QzqvDQebtbvyk/6AE0U/2B/h1m18btzBXq3WdlVeoPskdO92mGNDb5
ByainzIPnprRr1xQ3Bd4NgvtUOqLXRm513/3SKLoo6Ob+yTznh3sy5B2iGDJ7rQMMwVdCKzi8Brs
Gdttdd8UKlEEJwv3KBjCYcMvE9cMGTh+n1ZN6tFucDd7VvRycdA4HOUHAYDK71molfm/uHgvD1pt
4xYb9X3N0DbQpdO0UknT+A6uWutuPF0fOb8ZVI5k7N8ws+hmDYGm70VoNYjJ5ADUX0b7K5zsZOCe
ProrD6iW5G2hAcAjWJEUAMr/7yPvxGjAu53/3pC4Q6OX34IMU7U+Klg1QR7u5qjTG7fmxte/teJi
4yXJLJUXA0LaniwEEz+P6XJBTW+GXsYIXHtict8wP3NAWSMYiJWdMY2vgwVyi/NDQceTQm8Z60tk
M43MJslDBJeT30M0tbKflzLqh1PE9ZGCoOSgyt8y8Dzh8/AjTxLZhfkA93ZXGmg5P3yKmhSE9PPF
t7eHxPytVc3Xq1iNnnXOdJm13ksWrUP8tofQz7tydpsN7DrNlbDUTaWCYymoSkPTu90A1/D4hpxo
AObF9l9FAw0VVev5KshMoe9kpFgrUxth+rwkEaf0Ognp5QEynQSV+GEzJbv4IiM/50G68jqn3pNt
x/bu87mlfQqHsSX7f7n8q0aQq8Bj30ytvOQo+Ani9tnZQ8oa9Y4YX7rtszeJALe0Bm6i3Gwic4qE
WCy8lpj7hKdYiE7VIzs50YdmCHLnQWZCcDwu/0IYgfq59l9t/FJwjcU18FcmRYyPwhKjQailem9+
V8zKL11uBJeqCBBJ9ifzsWfhCEFgAdh1MKtJ2u+UXqp+WWTvNoN6rDmpfdA2DTCHE9K37zQFOq6p
0ws4HKt0aFfAEWYo7viJs0SaMSqzEldXQTjyVI/QPuGMZX4DTtbQz9Zud0T92iAXP514FaIO5OfE
j35+n7n6LcZHVRshJthE4+2ex1ehfvFD+/qpR/71gvemWpUF+SDdGwOLb/M2Hi8QxbTYKbJnybuG
tynnlPuQAzsn2scDBbJadeYbwqG4QolAz0E5aEIXMnCrx0CyMIRR4vlWYGPtYEOOGrXgkRSbr1Hm
u1aCJyYs5P+mooayWICFe1rn50L4B4VfR5rF0iT8MOBKgAU9Jun4RlSEfqGd7Z1OLT7xvAROjYCc
CzDZWyYFQHc3UMvOdkiLAeIQxA9HfUu3s1ojdBVxDn2MranjKCn3mjqJUyd6SCFEQeLGA2Nd3zQK
chKrvV7jszzLYdfTsfxXYmiBaxXp8szyIiaP+UR16AmB3Xd/yaI29IB8/4hPDU1aEpCnYpunz7QC
ZHa9jicAWek24O/3YF+xjWVfAewcodM+3KdnmLdfP9rmNo2rX39wKZj96id4neR/1Iqx5xOByric
cVODW9fcFW5mAwWYa1mPURJZVrBp13MaM7jvWCAEtUGIoDiKpKONTFetrhG2lSlGHCM64PASBIRW
csMWHARrLbRnkKFZvmrwWWyaJUnFoTsxpD510cT4oLqDSszTRG+H2H9pDP0gkUThpXqo5Mgxy6wP
mGKXVmn6nv03Hr0zYVauYKdsM0oLArrnyU80Qpk8SvuSlBX5LKas+WHviTy+drfypH+NjfQR6GNe
4bP7OO7w+t3ysQyTB4AjAYRI57Kk4Qwa7qgxNXYgjl5sDt0YFflpka8m64n6NNy5iWjmqQ33deSB
/j7TK7mb/JH1xHlFxMqxzI730Mx4cZuTc9CuH+T9xBswpRF5aW+/dM8CHfd0tHvGFCRSCFSpppTv
AvWyuvSO3SVVa9bA31dIV/5oKSeRWcANaD63yiaHKG4nnWXtS9D/Tb/o6PXZQZGjeFgJWK3LqicN
xlqBLHG34jgoj+/kqLWY/cxSdtcv6ER1S1eMH87o4fdvNW8HZ0bJjErG2xSgF1An0PzvXRW5b3gC
IFa3IpRHWhixjLKya4X/0/wnkI4bthlIk+V0c0aAqWPT/fReKBwW0Ft/Lwa5UkJ99lO1gD/sHjWb
YJ6h75YuphriMdbYhZNG6MTeDXdy8tbqh+daoyRds5dI8cE9G1581F5obQ/1cq9nN6J6yokyp4Xk
c3IL3RMlXowZMwOsQjmzyCdGwEw4qvHXFdYwNX4Tahs98euR3Pb/CIL9OGO653pkB1jKxfYgqH+Z
KIkSoyzzxn69xJl3CJqVmGqL1w8Bci9uv87j9zOA6v759GS22XKJ5f7UqV9MVBa4NtM9QutCd31H
hzV/c4Kc21uzwHOKyjLQK9hvs7KXnzt1hVYJNT4+eJCvxlQAFrpDXbT68ohD2EJnqcqtKlMGYaTp
nnxjvx7J/qWAZdd+qJAYDXGLJfcdQGcpPxQvsQ4u4nK47LawQkvuc4Md0bAh2FHadGyGJ+Lxviq0
fTJ5eIoFK9kQH85pDG6u5IszTYONoCt5MFi9/lRCdd9F9XXU9ps9CExuVansEMNiqmil8LVqNEqf
NAyzDwHdiCZYTfQSFP+Z1nI6bos528ODiqlT16o125As1kmFWGAf0X9lbdnwxiBOVqYZ6jq8Hct+
p1krxAGUovMeM6++HGTIkzb9rxk8Mctm+Pmhqm4IPAD6PiQ/DhtNZtQ36PIevRHXN9BYJoj7e73v
5uq22DxoOkngEZDAWb/l/riJboOV5olrjD7M8YYi6/cwrARFOn/zdcMwsP1AU3sFhZWJAUhNTTKH
mBbel73XOM9YtR2EYpEseZ5S35jxsaGNDFra2u27ckBC1iAoWqvdVvzQDgSIYBSxhmVoHNCgJxVe
sZHvBe07EOqnfOohFpWGX+iIqqTtmGoyBZqUVyMn2I0AuNexFTdYTd3kOr7arHbL1GpDedaww8Yy
7DX+i+NEezbxWWPio+BzFGANqi+08HK5bD5jaLHAk78Jkd0OctKKyqQ33gFeAcaknkcidgppX48V
BOnVe+n2FxKPxLy2ZcckbGAAFpWNyFG31Hrq35iv1yMwYii2SYVj+1p6o0DwdkkdYy9UwraoF1rv
SsvafWCCjy3OozPjKJyC0Hc0gYDYd3qURXUX+xD1Xn5xcTP0GIWSBndgQmkQN+/HcYU/urFaGw4i
/LhThpSJN/zeim2UK/cQ4b5cwT35ZTbRfytaMSJjgSPCposPHu7G3E6AJAUWoh8A+VWoac1eoUqv
Vek0U53Cg55SexWPrW6s+2nDjBHa4FlWKN3jV0MOJw4GzKMerPiZDcRvJDDJytK8d7oN/2C5s0uv
cQ8T/Wj/RW2F4jZtXkrUJgjNOVK3i1urHW+x9+WCXKkbf65NOvaIVCRPX8FEBwql0cbiavQOhLGq
W5llusJcmG9QuDqNCIpEnsgz28ZEMTfilEwzcSA3NGwm/Q0iyiI0eK9pNJhCfXAEVEEVj3lb699l
G4mi11d74nAUc1sCMOidYVlVo3hRKHbHecsza8+GzyCnd6YgL9hhct0bEE+IV6AA6FEyeVqzItV3
0GVqd17KkaamOzJ9RhVAmQidx8oZoh4vujbY1rqSFdxhKKfFqyyxRBryOFX0OyvFTIQs4h2A6+b0
Y1gU4HnHi+/dCXM61RmkJ3BPyFM0v8UL/GhWnxxehVHPt40EUEupyXsTsnoDHIM7GLFPex9BNIWl
BpMT/XfmftVosKKLACiLRwJTWNdYkBikuzXtNq5o5ALH4vkw8g3Ome4B+PY0t9+KYkwbEpgllt0O
+8cFLu6fQ0i1KKUx0C9byIxb5Ppa9HSii+vophvuXQWzjTqvpGkBnAx64Jstt7y4k3KleHooPmUe
QzxqSGd4QPctF8aOqkuK/cw7ZFYsWjWkwhACv/E6FTmeECAqBW+8FX7XlJ/xYcggZLpqOJKlWxkD
HrlBNL+xOARGqPeIa/iM8KV/kebrn3XMBHT3HyjXk8BVbelYLbQqXZ6ZLkPwyoUWK3igF62A2ovy
wlR41mM23bGShMvfknjOi1+b24LcEYHD+IgW1C2Tzb/aOaZefJqnzJLu1o93+Rr4JA+J3OqQbobD
lEAFoqL+P9nv/Qa/5oclMjClfr1SIsYi+kZpurikBRoGSaxskj9wcRa4tl/7KXRMHv6VZtRseCg8
FfTNE6v3Uw2jX2UWMq0FZGlE5pt8V3QmnyCFQK5g3OgpTwgvZcXpQFLRT5Ygpb2gQyzzHtow0hEK
tJPgsHtIBCSNoOeQYPLZ5y8+QmZiZQZdqOOuhkmPX3TQmZ5aBrOt2BiaF6Zi+eKoOJWB7oauLS3S
aTmsVV/g/Cnzk3ZY6ZsgshSoYBE0b/TjAUMjBkofMORqqbrzaEyuImcdmHlCmCWTopx1WkRx2/Rv
aWYprGf2mg1CnlHE7cRqA8zPIMrOsxR7VACLVHdsRa5kJTCeNbS9/bXhCHAsEcqId3+X15KFmFz4
j4DxovE5eJ/dl5v9y3PWRD3c4qSYHopfjZsAmag3E9TerKB3OcxrZ3N8ApI6vwp0dkwaS7c6RiG/
Z6l9RcshcTE8YDPbv9zEMuktz7nKnns8HoCVQy9afHbNWjmH3e5x9OOf+USgycqQ2hWqYL5ESJSd
r3xu+n1c0Er1+xRbkj8g2xpROsB+QYd4USLNdQMvfKeVDW32RiowUfOVQfX5Oe04OL4NFPsRawG8
03HVd3rKkyR9n+hpAkji3aeMakKaxN2uSuP0hwugh1YfuCQMJvmwptnx5I5NbK5og47fLrYcwIpZ
kgD1z5KvTldU1XheCfn8tufOvUa2apVFeOZDHbPJRV/TWgO7wqXixhH4ClzkYZdGsrNaIEciv9X4
8bXqwgpo/ww3V8KbQMbBaAy090CvLkm11j7iPD+uHANvJC1eMW1sZQjC3R3T29QNJakOyqgRHNfu
r453Q8JM7HkT5NVz0z58Py0rlMuOqNkpSzI+X0ts3OwAJ7TplgDEfs3XmvdypMRFJWjNkvbMX4b2
4IfV1nnwSY647acmcySuzB0Jjl8KQEaMYzaRzemm+iQLiWKAabqtk5SYbvFsNZxvP5ulNNiWpuH+
SYpdj7Y/Xoc78L7EKl6thEmuz+beuQ9GoJAx9q+j9FLpibYAYbhoP8vYiHA/aYJ848ThSn9qrL5R
pFJY9MWTGSzSq6Xj6O43xBIMlYznRCEieaTwTWiOdJX4MfcEuLYOHdkU+BKR1hRq5gQ0vhP4V5a5
QrsomVVl3fH6Kjl9xzSR/LIa0AeXUQDkqjC8fUJZCBQUVRs5EG+mrqtoyInpEh7sdtA5Ddwno5rl
oUeLpM6MqamVVR2vMvBAJHnF4B2DkALA5xF2gZkBLbHA0vNMKD+07ymLv5KgFVvofMbTo2DoewmF
KQ7Jx7gZF1rld0yb3/vOodoF2yx4Bw2rAfshZAWGXl6XMs86adewjIAhxK5HaL6oRciG2jJ/+ldh
U4uxrAWX53ogFeKreFvU8NnF+zW4SXQZsUXc9BIA0L/B3ospvhrZKYtAmWRpMvUb5DXh8EZwpOsI
mEop+yWAaxXHX4KKcaF5oK+LL77sWLH3Lg4OJOA3FKVDo5HBRf60r5Agpl1I/2qW0NTGjexiHYtA
qV7JxMdQBBFUAboappmDeFYeFMX1enrMkWstdUznCmsD1nXBcn/EjtLCgkaT43XhBG9J5XhO7HjR
7nwjbdH4/Jk9smfZUa1tGhge7wdOdcQv9v6aqgIIJiaFPxfMOfzqVwVPxF/zrtob31Ky35URyxZh
FxvWw06zV3zgJNTBASQ9IkvTX9v6dYZ1BplYvWnZQNqQa+txQuvRtpiN0l5Oxvt8k1dVzrvL/fDm
D+Glah0SB26BsexJh9nR4atioJ585kuKO2mVGUdK/hs3orTeXVgEzUG+xU/RB35h2OOeXg51l8j1
zQoVbBnFXeljlQ++WO6kqt2pioCR8Lqiees4LcUh/fI29ZFVBtXESdW4x/VobqOIZY6qBSeCl/cT
XUMv9T38U124mM/syQPAWh/uaDmhiwFYmrrtXl4kn0GcRwi2dq7fLEC1pFgw8eka2ZLSSPDL+ZIT
1uFdIm6Q0shmkBoVrPhX57MHLFu+bdGz65ocF/AYWu29s2MPPuQxbE2ZeOv5Tml9AdVWRjzvfw+c
Ae2C2TnJel/BvIix4p1Z9Z+R4ZFv3q4HRbHtOl1/HIttjQSUPQzNlAhRlUgVQvh4WH1ipucE2ikd
EMd7bBgswmvdkBCaRx1k192cCUowipqQrx504SkN1FdYDB5Ccyi8druURND7Z4dPtbjiCAEdwD0t
zE8haDxtu2NXvFGk6J3bciAK8UwNXGFas/QEx4jiEZRLMQEcR5Pryc2H9WfgSGSJT9IfTmoY8F4R
7LkGBlDdE9tMlg44PLTXrhaJBhKqz9PvaRQqtPNGxlAtn3YpP2O/tyuZJWfTH8zWeLojYEdvCw3J
97iPYyqLjwn+gWOahIkpux/wDeVejS1Cm+xwCUosKcdqFEH1T9xEJLVH03WEEJxNVLPpS5lxyCwe
ym1WjmHZbLJMia6YtZpo74hA1sjCtO65VQ+etWunOgnE8mJ6SVTJKdfYbXlSrdRWLUoEAbpsKrdU
U+Ey1szqUyahf5DmwLsgAqDQdum4LIOyWuuqL72cRaGFtAjSIHoBLvRTRZExpZIFe67G9MELVPVJ
Nin4/gpC4FvFg9dH8cVQyAT70Q2M486ugrjSRtvHANmYAxUufCtXp/99aaTcNl+2YPzdyN2TmfQe
67s7iaoq7p9P7cLF9zfMGzPG51ydHIYXux9ha9uoZJsY0sBIiGcJepqCDjra3ViESUhkSIUAxJsR
xcoI9pPELPRrAKpBlECwnD+zOT+w4gyhvP+1gbFjYicHlpAyxzrWTO+sxNz/JfBBjov0hVqBN6K4
81+qyv3j3s68opHaC1TYjhhVb2yBJgtd9icmhsXkD3y+WVSzkxnentcujrOyAjo/ioiMKqNESo3m
PVfBveM4WDIabeQW0odV4KbR1Gu6zArWVCT2orfbNauf6JYm7TCGxPEC407YOKix9QHSRu2v/EBT
UTVcXXZBT3OV9oibUYU9gRgqd3kI8ilhfskzGoKOYZehjKbZY/UzLgGpZqzVizDqFEUcePe/oCXG
IxwAp2PizUvKI5UgIRPFN0HFfyDnqpYGc/mqBkRSrQJwJWda+nDKsOON6luxZf1C3IMquioH66Di
r5EeuKPb86eZbOoe0fW4m0w53B3T1pFjCcsBWQboIP+vT9bAJmEfdKujLwxWOcx+8seodWGUcDMB
HNvJ50Im8CY/10EvGu7ykLgz+XwwK6SlXVb6ep7M9NZh1XjcdCppmDDDWCo7UmUeaMQd/bxUTO+a
6DWftrkD9SgzQkBO1p0TJMU943JuW484+Lgseb+A6LCLv1cdh/tQPWsy+mfMHgEGmDuFiFeFskY5
EtXlGzQ8YHIOzcGeDiWk2qj5ra17deMkSRkK+zTfb7BHs3MHIdBRNHRL5AyBD5mwPmdU/OA0jjXP
DsFd0nKcMXpDZqENxzZpuQMX5lmHrpF2jqYBf06ZCeAOykjyeats0BIBd77QzhgtbGwRd4N9MUQK
tfofWSywGmQpydo25pZPcES89MwRLXyLV8nOp4q0yaoICAcZtxCWWIni5UI39c2EnpUo75R2o1WR
ZiyXG7wXzJ7kxkh36mKGW3OHZcmzrIwPDs71Y5VgbYxfaZ0WzQXURg9Gc94FtaSTJpsnPOooSvRU
wgXWwApJ/y5ibGcPFhxNVopEUxXEtTgCDIL/TqMrtz81MlQR0ASahEGCBgcP+iy/JgF8EhSZ6mTK
h9s8n1jM8anCX8fonfxmCku0qhqiSjK4nH8HwLXZVLImtoaQV8n8r+CdYbACzUe5S+0ADdUYKuO8
zEeGK8MyMH2xa0AUNvPv5FUhELnkHglK/6cOAdt787SUM1LjuRbk0ybb4nmJ7fY69reNwK5GacDm
NvOleuAGLY16BbvQopaWjjeb7TsGS3znxLSm4ybehl1LXP5tN0y9lVun5cX9qkqS+zY8r9moVCeS
Y7VncEFsR9zSktF/UD/6mfmhyvZHc+cdVvZ0TqQ2QEaaJFhyi2gkZCRuX27PCRZpeMIGiMy5e4w5
fDnInKn4d/EdmkjO6W6X0i+ekLlfg+2zqEWd2D6UCX0+7Ck07Gf34dYCVPOtZCHXpyUD2fOOYNhX
G4clocBQY3c+I2J8YwKVr73IPXXueGTTusF8pzq1ieaF/uhGVED/RPZ9Z49wv9A0Pcg1kamvEBQ2
+re+KuAxVxF343q2oWUTjbHP6Dmnu3AbMpuQXVExAJl+YYUumWYguubZ093jgbeKExs1M9jP0PxI
SGD/MkHr1it6CsGN0vJj6dg6NOyHuMceatbcTwPDbTAVHTW9OhHSTptwDCvRQv2Zks8fmsoXH02d
/Lv9IpCiJIuDOEGX4EgtrLz3SQ0ACGpqktkbfgRU6UZ6XiVV8dYI34vLhIwlBNgXAniDmRkfqrv6
qoNp8D8WdRI3MrmUUy0Lrfzc0RvcXiX3t48MJn4YwATnPlpV7NHqCHjqzlt+KJSQQAwVrL5f5hJ4
n5QQ6RX3/oa9whv1AJ/BcovJnBKi7ADDsftUHwDslVo5cnq1j42W70CUin8tey78pBHczrqDEQGL
ZKYds+CRLtruWqXTcZ86Az+x03j89s2OJPD71FAOlRjRsLJO0L/P1L8gBC1Sr6NRdInt8o+af4/t
g7QucbfEi0EiXDtGlY0CaxW/PNrkJ4jhUzZXueZJ9k36JQsbRpLApgGr4GEJofw4rX55j7gDHICZ
WrfHkwfoBzzwCdmmMmhbzrZTILb7r/Sw6xzQYpCCRAyFsCfd2a0rDIzUfv7tBE5pwIazTQUyGjIp
ykooTwuvq7BXlNL4DTWSn5IDKTPocCHBZjIgW7xjSzXLWKOCjPdGGJZtO56Bl5Hp2cN+jCJD5Rjj
9Uyq2uUBJxLySwf2j4+dzHfBoKL5LmDHW/FkPx2NF3Iz8ympwLG4k+vDHnd8F89hn/VP8NpQgebV
toQXmMFNoQL4CJh28GCAtxPygLCx/uf+NAeEcGAx7Zm1aNEDG2c10x/jP9p8w96IW4+5fjRMDIWD
7YouHZblfaXJJa8wS74aqUmqosMuzFujspRC+Mh7wsjU5QUiHi6Pcu2J+lHkOKZtZ++ITaUzG7YV
1HtaFnIjfgmjQlFGeCMWfGK4X8hYFjpGB0la4x5XBzO7GaHHEumnO12kxmAmlJMCEmCl+vV5SEv1
9CXwNPL7B8RWp+1YrUPrhDIGMMf3cJyBF8ajaaHee27MnKq578DNZUfM0uR/hVx7KESgAk0KDTQW
wsYWt29JoeNu2r4/OFzLZCdyOHH+VxujCt+l4ZuMMqxZ3wTFomm1DV/w11lMZQ/uwrf83clQNN5Q
JuQ5xgUk+73vTzojf5f/x8k92EZk1go2WId7nFYUi/NkCtbgTV2rLIHBKiJaUKYh/JZ4CjJ4Di3M
KcofHDJ9KBeKH7Ef4/S5+vFVl3U/6t8OWner6nb1VTcjikdB9OLG4OyT4LAKUSvr71alEw9cq1vA
eM5Z3rkH1SQ75ccl/3KogiUFwsn1rRcNqsO+AJ40o+uMfFjfj9JzBJh/4hotoom3cVIlP7rwG5Ud
oIfpjLJi9knNGwwjYOC+mNIKnvYGm0pTxx/uucK4Oel+G+Avjdih7W8882y9W0CSDrzSW25ZEdww
MZWsUaRNX4Y47ixBWoTRyG6Im1olJIUgcQKVmQykSc0exCQQH0Nr78OzhaYZSp76Dg2WI0rUWX7E
2cpaJ3Dq0qoNVZiFdYCPduMZF2LW/xJehT+dbc+UnWdt8dJk6W9V4FwYmwzhoQnpJl3VWFTZtKOW
aWuzcBbHjM84bbcCTrOFFysorc7gqOw7Z5mYeHeRQPT9xVc/Hl4Eonx39imRGnY7mYPXo+/09iOO
Zhl4xSI7FvcO6FJjGmlciPEH0KYWKORCcbOcgaSTeFjYiAYZbPrTy/bU57z46zK4TGuwcd+aijQd
1nzDD9uDzpVEk+gOKzUW0X2p41PksDZj7hRLNM5t32/3rCoO819B89aYylh0I2GvMsfYtfB1qhEH
C3g9psg1n4qVq2TfJzL8X0NFpMhxzNlNg5vBVJVjh3TiVhQNos55de8aT1usczdfCBT+HjfObPOc
n3HeUaLYYO6qIC4SxLh9BO5NvzfuOBlrTy2WRGO4TWNHSPYEd7Tme8V2U+3hAHzDEeZgmT5YEsx1
1uQBQfEDM2dXdVgVCZT5l4zERWntQHKC/AzKFnhXkYwDmsSg6evo+ZOzZgjlwWqMPa6YTZI3TaUP
bvk3Qh6c3re2lqZDVkaN4jya0b5OIqOPxa8nUI1aBoFqLFEXZ3tWQMV62nhrz257IVrkq0NM9bTV
G4XhYsSmo9V+V3jovwXBr04QDHWZ2sXM6ozoE7VnPZ1jDEIPFPPAiSBeA8K16PNZqfSSFDtDBEZD
rsySMpIYB3z8F4fP4U5zpRKdfd58wUAmaJWEvsJ5NESeYl0oWVrT3ylFqbdBAUUGUXqZ5Z60swNJ
mdad++f1gpoLyZJWGrunPSOWjdo9uwAA3rhtbyD1YbvrxN7j3BYSkRhvgK8YIlojzAVy/TsqpiMM
YMMoTR5GKBRPjbp3IIzLrorimvv6bR8bhahghd2WhX7aYNF4lpYKEOl3XO9woTJUy0wjT1UaIdMB
h/NsQBvKc7URBNfsVZYzJWljx6dEL5i9SJWrQFGtzqj7JcSnlmbkJ+ZEc2wt2qJcH8w87e5vH5gE
uFHpjEIA4IrHgeiz1f6pDvqo+Rjpdce97IN5854EOMqmndsN/2e/yfp+u2PAMsnPl6hqYsXVK4GO
0JOwtV8In0QC0YoDRGuBRFoIg3PM3/aBN1MpJ8ps0RPHsXbFbebnEE5uLi5nN2/cK14ZAJV85Avm
tpwL1nqmngCFYdQ9SOTNmtnskIWTf3CjrleFSuuXbIcbQfh9ARSBPcpeoWESiXAe4ioQE7DttP6L
wNMnMZTZIdyBZduK/LptTDl1mWZdDwvQNcLusCdhjsY8mnW/+jsAfamiYJQmwUP6PYUrktfKWXEd
vdiqVY5yoqpNgEOGcMBdrw6Z4rShdl69L52sRoe6hCc8uB1xFgKDVvixHQ0/ajq3Nfd6RgHg9qW7
X2oV5hnD/lJTuRjEYTruyFpd/2J+FK/QBvq99FefAG7MZyD6euAXmGZOR/UoYUtEMKR748PrSjb5
P2jVhPCOe3G6rlmQjH0q6MtZY3XkKXHO7yjwntq2uoJOOHw+tV8MojsgF3lCjD9N2oNfygqL35Sw
pXYZj9nHS8kso4ilayobg51+mxta36cnmPhH284GYwjUQvK/tobJjrr7oL4zS1BeDKK/EA7HX1yN
KdVw9QNJH/pksIRpgvRTE72H2/XkPkrrJ+EA9UTASMhaG1K3avJzyiQGksy1VjyQVW+0Sar0MmxJ
A6sPPUnEHP5BXrMEhTr3jOqEXghwOXurwYnbbk3HtdlfzvUEXFMT/Fi42vYF3HRduxFYYktvBpj5
ymNPmH4IF8pm+xsrDR5TJ/yDd3ffmnsP+ukB7qwzC9hFMdV2tTzIZYSiNEsq8qr/6PjBt1tYBhmk
NRHqN1ylMTDed96F1pWdfyeuxdNY/tkQJSyFzJ3NEKKv5YxgMSyXT7EKJzjdyZkNSXiGPGW+F/Du
iKyFekO6s6/8h0ct+++tMWgByfLQCbyMkIRMLU4It21VkcxFQJzOJkN0Bxi4BTVnh308yPhXZP6y
rW595FQh3RchfGVh7GifVbz/ZHM94+dSCcPwV7Z6HBKTZeDCmd55EAYdr4/rlm5A1WTCsSoxzJFk
mf5z9V9ryiFjx61DM18yWkxiwBN5vIP47M+/u6DxtUM8COicIuz+63ZerDYQ+/dTkxV2bL0XSEHj
JB9XwhLw1IXXD179HjH1TxnFJzrkzVEnhz9GmA9/dhsdPMXwFCOgMZTh8sqlPzEuHTHsVoQF6tHa
QBTTBIbrlixPL6M/Q1/WFZY20h9NxEZ7IbvLgErTrOcln6Bz+EmwJIR4OxWrQu4visk1mOhefTH/
tRd72TbwaekeZ0wCqK5hhlhBXF+EaPxBTQW/5EzHboGT4AAAIshOq77qkStmB6ikmqRsFqzlkk9D
x+CsUQsQ9YRVyyesCk4edNQ7KP7TdDLcIF6KamES3A7uV3ZwScbZgHDSSNrs6whjBRHSzO22Fj/x
asT5vnnGn7nOSFKT7PyIfzmxtzAxK54S+Ugqom3NVQcq4k5lbzs0/hmuOs4cKC9O2kWW00RxTslv
f2DhfEOKQ71AeixdrrzvGnj5pInSEy00J4hiLozT3biJuw3KIv9lueU0RGdu/g/nAIjjRXy1Zw7s
OywnfovXvD0ggOZPR1NhKOjC4Gkt7QWIlq58RKadXudqGovLxzMOTs5nGndxyPxxiPqGU9UwoCXE
7JuJ0cg4EOQtDvbkholGiPHzp6kz/KwnLJAaM8ksDr3rVKk+ZlusjwmYEaPKZGNEN95O2eW3SE4/
VjALO45sWHCbuTlyfkaBEYtpUC1jknGUfIel8qVpV756o1fmMquL4vCdVioG3U7xL9rInlZmRVN/
RzJzIFx51i0vZVvKXF4HN65PfQidvErJbT2xviefMSCa1RvtzX67wTUcA2zCoszgQ2oIEik/mo3Y
NIAMKRiYUm/WswK8BGfX5cuXhgGNJx6IXCnz/NGmiZZf2fbbhJ27Y+MV8s7RLrDmoV8Z/Seq9JFB
BApZzZwk77FSOxs9gbqTTTvyJZn5WMslwsFIxZokYlcpQtCpL4YLU3nJVD+e2SrvOOs4UI+jm5f3
BnP0UVZoqv5i5gBuIf/D6eA6Fv1rGTGX6aTd5V0j/l20mJ9/UxYWKKOROzsRoOebUnBYcshpwsIb
/mWm15+ug+RvVQG5Mka9d12L9PTc6I4d0lWz0dP1hUvZ3UjbG1pwVta2aHz9NpRZGRBuE0hCW2yB
1IeqcRP1+Iupu1Xl5iPHSPNUJPYpHa8hkwG2pq/BPZyEiSlm2/7+YP6zCU9I8FdRMhSkgN6v87CG
BWOcNGJk4pDg0nIUt0ts83FzcJQgQg1Vs6GcIu8ngNH+ZIiWr+toRUx8fHl3n31aHmoO7nZydhMm
CO68T3bh+CP65T8wsAj4lvSWfXntJoVTY8CZmubypr4bCx7b+azZzSDmp2d2OSyPy6ojyikv7Y5g
vLtYVII4OsO17hGm50XeAJGquY7FPlVwHTyMPm9vtRW2Zi4uShgDsLiR07USz/E6K0Tlv7nq5wyn
cZjcFil1HOQYq+eQoktB7k5xLjhV14JWEBNAjC1kpQbb25PfvIHsMLIcY8puaKkWOab4GXdfB/iK
Myi2Z43R8Xo+ZwK5BV8ljz0Izz7V0EOLvklb401wBuXsHKUjkcrIFKJ1nDEUJPcMUdp4XFntBdBp
bpSDd5fz75ocv7YoQ71L1JdhFMZOvNvwvf9m0NZzN865W/c9Z/6cNO3CdoKSHCYEeJoXASkWqA4f
noQSPxRLjskQa6c5lL1UdZ2XpIQ/v64m4cpv8BO1Tl8Dg9DMAt3wcmNAeLu2PDUIqlOpGlOz9SBR
3jtNtMcq0nyGEmNHOhDZ9DmsxsfYu5/I8/RN/pekMLkgZZ3w68rSa/X7hZxurdJsS+7/AGiNXOJR
opGPhSEEcFpMdHi/Ijq0dd/bAdE+OHinmi+WSKTLUIbX78JT4UBUDUoM6hTUeE/T0FiwFX6ycV1D
bOhC05t0kGoLgZM4QSWnmy1Nli9zTYu0nARIPV6cXQ12HvmfZfHNnd6aR3KLaLwAFRXRA9Ssw7d4
ITH/x91TMBuwuyrW7MiL8X9DKj6OagG25diZsEDxFtLaAY8faj4zv4SUgimSodh0kqPgwY65nBAh
j8uiT2894/a4+qnblUCztbWx6duO3+UVK8F0ZLz32tW7p3IAmZjHv9DiswI5B8HFkZrc643ldw8Y
wthv4g0XqGojQDBJZ1Zxyu8Epl6+HbW8Ce2Lw9ftPKKrhP05/LZKHfSlHR7l6APiI1c31fiXnJh2
HcKg+7uMYhWk0tXgUrgC1hDxqmPYDlaEzo5eOOTyJ89HKXTsEwOGZp1EckiiWqJzxqS5SOnqHQOr
+EqeD28h/ouyj53gBohrvoiQNC3rtqilM3s8mGW+lTm49oc1ixxJxbbpIJYrTgryWMnJU4DmuPof
mUzsgdJviEx1VXHl7pY7QLnwo9DtNwT9ZsmHcUD4uLXEFEF4VQXiUl1nlD1wFOQp2oBK4qRYI7Iv
E1RxePZ83wyNghAcjdQKRGWCNFV+IUODe8wYztqdAAi3mGDIn0MvPf8p+xU9fzWQr1I5A9F4AmLG
undl6UvgMRxr06PHz00/Z/gKQm2/I66I6VOoEMdFf9sGmEgQZ+XnFJSW2imQqTbOzAtmbc2qaNO1
bKGtDBxxKiOAyrqCGf4fx980l07boWv+JebYwouD2bVIknWyrXP7nlFqmEcyb67JBMsqlUeRM2fT
SkKfuVn0hGQbCKnxbGsICG5i7W3ujA40kIk+egS2md4i6BmTr/SB/xrVReWualGlVOqdA0YoQZTh
DN6zpEOphThXi04wt6mmattSWsE7kQOvoBDlnWXdxmAPcKQ/1n59I0fzFce0yoHCRx8ZH6Tp36TP
9YdpnXfe5Lae/R5GRhzEMCkmmqWZh6HFcM+oN66IDMzrw0sHzYcBAmXY3zKCfJSOaoScfgzP3GbV
MG2vwcFcHfM35Mpr138nzfr7erugDPqUnAxBFRgk3IezbAewH5cA0+8APA+v9SgSzZL0L8zuDoi/
R4NmkAf1ikEseWpNKXkXLRm7Y7CSemgxbxh1xggqjHwjn3XfVem7S0kwly8rwqT0a2Ov+2amxJmE
LJ6FBxRqjkdLx5Nr+xbi/vo+WKIlMo9A3NmHCmkAOPhoCStyK2zJ73/KU3JWvJUYPGAffdE5Njit
3P0wo1JnOIKkvcHy+NJ+UM6iic9Tv89JxZcSChVO3JbMy+QqFGrEKYAcbUh//K+bViGDKFcQpJVh
4KxczzDQfJ2gjMGi6Ky3h7IgTnKJfzpAW50oPrqtDdS3Qwus38PT63ssNvJP/5OFDluHc5m5tz/l
8Y+Z0dlnfKN/J2Bl/cnguS0ln8gOU69xvgglQwx4WJtGhlRz4505gyBXL5IBpxpiRPPwIwI8D7C6
CLpyqCxUYAR2GSk5CkBBrJT7oqPYbqNT9MInlteTpwEvbxJKZ/IkMoEb1/1Wo9Cxyk0YX+8nd8Ci
zeESaUrUhJXNKERsO7NsRPAk79zzL3V4Hcc93sx/8Vxdy0/tHCJa1DYpz/fElam/0lwgw1JKgF1y
77Hh7GgAuxIpj5vxHuHzplmIzOzRs3IDs1qSQ2mXgyU/pE6/QQPWv7z5ayiBI/IhNGM7PVIEdVdL
dI+PJ30npGMsPBck152mbWctJ/t0Xq0ftTisw8xvJdUtWNLshtYUtJ/dv5pjbJD+bizko9rgYxGL
afYy+pnCkMUIZl/bmKFrcBGbiHnmQUaUQ9u2f1WMwdZYxgu27FCPT7ryq5N/rCpJ7dtuSfgazrEZ
LfjAQc3K2xC1f5VdBh4+PQvo5xBwNYYr9d15cKX+sggygkuDQ8TQH97525iy8IdH8ROv7F7ihWn3
Y71dYciIrmajib+tao0tTkRjK7j5BqUUH2BTo+nIPs9JtBRmY465m6umuyU5xDLMZqzYQkbdukch
tJUDoadB1jQLzqv2gcp3UnutLrKx++cvKz+vKHAi8YeAgA/R3Q7HJ6q+UwY0u4LXLyKBi44tvH55
xbyoTc/DRhvY8+cgqKYRh09ej/E8YdA20SBsN2RrG7ou2W1L89rKARsvCD3Yyc9ACM8FnfPOiyFA
rg0o9FYPpC6WKghnAYo1+c8f1tM2UP+Y/3r4psI0UDR2fuH7fxcTAplzsOLeAAYH/nJxrOsp+nPO
xkxM+PKjtvV5lEIOTuDwsXztq4JylYMVWRbFRyrmQBSuPqGKg7G9mkZpJd+uoRmY71HYgmPFo5tB
b4MJXm1QKqVI1A2s/eyLK9oONhVEDBmLVGZ+BvVm2hoohd+qlMBuLYVmf52aNWKPMYka7Pqd5dGn
e3gYFce/5pzEhwZTgXDafrqSfPwbmF10oE9Hfdk4HsDgtIX0QSbYFQ13XL/TNOVKteCR3gDI0Wu/
jaxw6LPk50T3LdgDBC7WQTqP1pWRXbwx2c5U5dI9UPtcldK6ohiGkKuoVipTS+Kl2YR6Y3iKv5XE
v+l7BwwEwwRdjW8zXjkSMxCFfmrBGm2URxP2z5WJmbTETFCfGfprLqhhlqUEiS3xqsE7oiKLzuXR
SK+dgM+ErcIh62hZJc0rnOYq3HIXsyNskdi+ebclYctiytBdqJ4y7FPaLnuPBWMdn3KvWqDFE/oD
Jj3UH08mUfb1t8HG4MDomeoAo+aIsdwJGR91j2dcipGw+OttMU3aX9yPVEu/rDVAODOMwrUprtOe
hiYmem4mGuGo5qbPwUsJhAXfVXaDNKfQ378cQZHcgib56rzgeOqklWoc3eRa4vc6pBtcMCWMSMU2
LswNMq9Nvc5cQyUUZHrc7kp06E79fk1hiWPLEgrDsD8zWKVWLFQTuP53hT0/+lAUTPif/rlSpF/6
aGbnsz3tTknxa7JUABkcmY3WiiQG7DP+vcVSw8kmR/Jt8TRS7tO4ixDhwIBFmYYMKDlK0YqVB07Z
AbqONsfAVtL+/AZziMnu3pnxfkxsNJrSBqnGqHbjDiiORX/SffiwSvCzHjVEO5PJINX3nyCoqKXg
xdHfH4gVGEFJ4H5fXeetq/ZUQrYdTDQBzLt/ggeW7mbnnBvaCmergUM7BM/6CLLe0Q08Y1vp+j6k
IUD1ks2bGrtknRDCQgZppBGRRLqAlupifBCPYWsSMPKolTgB/lZnkLvCY+DCwlio2SeoDxxJNMud
0g+TpaUyuuuDFBwf1ueMUEWoJW/Z5661/Ng+0d9778Xd+gzoq2Ks2Z17oQwjuUSxc1Rk3XVjWHMM
rv2+uOYc1+70GexcIwo+NAaeXbyDcoJp3rBplYkAoPfoXFKddXAVUPLWYPKOBnv/ezPZG453l+cS
Olrq77S+SFUgv+q2gBpL1Zzp27qmzy2v75Oy6/TWvzhFfEAm/jiDa5GEdWBqOdhzhgctwv6GqP73
oaWrVMzLsn3nhQpv4OXVUbj1pfNcxpm7bGsqT//Hl74lkO+Gav5UQ2bUDEh5QbojWmqVrWy7l2Hd
o2pllcpoT00S5UUA8/XYz6Rib9NYsyI6fb87BhiAxsdlbKPpz7/oYhfF10SkdK/sR1OfdsL3bWGd
fgEcpay+7ZnjoJkm7YwAt8D5qwG98mVwod0Zropd5moG5gR6WNJdtneZ98rGH23sbW7fsLp17Dld
nt8IPtcYFTabU2t3QlYw/Ep2o7yq5nFw7U6zpbObXqMpovK9bMIzlvFuK+N3oQm82RIn3xATmt9k
qeu4giq3IOP1nhaV/g1Kzq/Zg4qUMAqL+Stk4CXvvTceG3yV0s2jnT2AphT9RcYvTA+l0XoPbkPV
8IX8ISpVmMCbO5swH1dG/Nfc+gk5WOw1FZDpd0Q4UgRX6gNAaVz6232dtiSGb6/vLr6rsN+DjVU+
eNw3Ht/5BGMcIVffQRVjlJpb5074hKjDrOBOiAipHU+zIGEbI9LteE0fVPXMjj1J1awO4efb9JyT
g1fuhzbzuF3Nwu4IhvfJOi7Mqzp/OhwhMHs5iJYtEHMew4HFmseDr2jgGIekoerbUy9UZWMdHKCx
q5Pfy5EylqSC1jY+n1LZOW6VxdmhDx5toM71xqQPVaL4XaTEx2Jb22jFHICOY9QcohZ7JFCT78UY
IwLme6crsH7uyRiAofs4uWG4FgEacTsldEhVQoioXoEW0Os2ik7OFi7V/vqucyPt9EZ4oaDaWgw1
CdpAi3sI77Smx+Zpoc33Zk2XYx2q+GgFMksAmwbNs4mdaidplqxexza73rOgQ3fD1rI7o4ftXjE2
yoN64e/S0lQqiNRRTc70QQIEH2lMsdKByhz9N52BCUNt9v/dDuq9pnpe6bL4jGr0uKG1b10/1Rh1
PmOh9BJW3N7Un5t426uovHMUscSOQThIC8YgY29PguQmKQwCxeNkx6p3psS/Rqbs0I2+yaQB2UkP
YukPt2i2jo667cStzh1LtR5e6OgZ+la6wg/Ffn02dMVEltnVOk7r/FxHehhMmOlV+9lz+F8T+Nom
KmzxsiuZFRhssd2KGLJyyX1EP1BYDT8FgadOzISEMC2zqRXUEdgvYoICvyGX94g11t7AyuK8vWgs
/yu4E6APOFG4/J8bfj66QHZKXHozwnD4yMj45YkqR1n8dyDB1ICp+x+//TsF8wX2Qw2ayXZ+Zzec
ltVkEAMz2NEnwIz3Q7+be/NkUHobesigCwkpBmNYEboEYgR29JeQ3BEvZX8cLgNjVVJrw1REQ2L/
EJ8Qo8bVQs17EmF1gLtA9e6S19DqSif+f6L0iJNd7mh8eLWTY9RlAPkFhD8RguVb1ssCIcfdKBoV
pOSUHBdcUAjdcUhMoBU0IBP6jpsLw1cmVsPQqCYF5rRXUSZdy2a7JGxGXg3QqPxS93vtmUGxY0Ku
TtrsXWHqNaZL/NDMOhLM43w7ecMievOKNazYq0StT82DaUJgLQ0BwBMA2M7t9SNp9igylHLBtzQy
sAqK6H6PSlRBfZZaqBTiY4qoW3qGEHtufN5R+f7ShPGFy36ZLHw+SJtvCT9WXoXVEyMPeDJX/bLa
StUaTIlM7Mww9Dtk5LDbfZk5nVhiOK2ZybzJjm7j2SM2WQJR3Z+CB0y5k4PmcuAxZD3bLAnRXYGW
fUsAgndFo9RfzQCKIduMjYzWPHE2jOV0T6DkmCootbq8lP2hZ7/ECc9TDwVYxvYpZn975X3sFMU9
Fjpuvy5RJ/Rcw4QKr2caynwgEYLQqTjW/r2kse6xoMiOVutIwi2OvaG5O9O6XxXDikTIK+la/zNT
nHNqv7tbPHphZkNtgOIj2eGvuihE//jnar9n+LPZeoZCZjZFa/Qw6ri1ekw+sXEcJUXjuEBklAjo
79LoBGmDjZ5hnxGMVPPXHdonA5PfixxqpO50M2K1IuqCETtDuTeBby7oSb3nKuPeRLU6w+YQK6UM
rznlkoPqqBfwvSjQsXWfzeu/a3EUOaSdy1/ADmSYePzHpdcadp+x77n8+dFzsUoMUh9Xw4uOW0vd
6iR/0IRw3DqIUalF+pdL/55mdLzd28TYtS/qWD7znjT2RADj/ikxjZymmLememlvlHLupZiTTrxg
q+YarWu+yuA5oIn0slMtNQmC45xq0Rkl5bm7gJ7FUOQPRAaq8LI2b22XRD1IKnypEy66jZrY1u5o
1RFOjqlfTXi+r2z+NEzrovO07kaficnB+4/d7hfLOV6s6rgaWboDGQ7FY4dHR2WVV8RTEID3YnO2
zRzbNku23OJH1fqPsJrXmoP8aRavz9qv+fe4C7rlIBm39bzpqIqGON+rANoaRJDPfkuWOxm5BgR9
hEdamUKpc1XcAyDJL7afd6ZkKSf9euZbli9bcN7BHw5xCtsJ5jAlzjzDVvSdouVBINwnXi0k0BdM
NwmE4GpSmx98MmDm4T9lVnwClqUcR9hdNLUuB2p8wbyLsB8nx0vQ2mlU8f76Zgo3KpsfZ/XbOnG0
v92WJsuNtSuIZzz+tO6efEe0QZ869vFBJiX+8FoB3iViObtwGELgElSXxaCgFTAwDv0p0xvYQWAM
hiuX2g2s8QHsF4FmgSNMWa1g38DD4xQmtSYwyHBqgMRC/ZLVyP0BY2MvHcb0fJrpsnkyJgZXrRXR
bGmH6HICa9TX7UkqQPi3S2BfUUbSB3PPTl9zy45o/1xGx7pAkMFGqoWLcqpjCdpUQUveu1OJATaR
6jKWc6dEaa/9k/cdajB56vK+udRNaNZw/AuzFwhVaU0uFLAsJ6C6dDtvAyQ0vn2zVerbD1A1Pf9f
Hsvqc3JHdBi1s3sd0N6PwtGHyvqlI25ISSuz8yYnwnxTkWAJN1Fxkt7SOD5NBuXuJrqY4HmgnJiL
SIpkihQrgBOJxOLdkdYiZ0j/o484QjLHSuJHBaIgLdn9mcJrAqth7FmeGMX/rrzetSWkPTPVH6gd
qgNtmcTw6lY3uvaNe+PSfEsAML068SKFM+q2q0c+4D+UF/0iVCjavhuQaMsQrPsFGk057Yvyhq+6
lJxs+XF+H4L88hniFL5WG/BSpL737yEKm3iEtQkKBhBS9eS2A6oGKzzNwPyr+Jko21EAJ8kXEeQZ
S4d0J00qQbc0K7yRmW++5/Rm87eH7Cs1qhy9yIFgvjZgnYOGzylcfwPN+vFgKklPMgYU6NEx0VxK
DRqEv5pONkgadyJqdmxnQRox/+REQHAVfophGXhkTtHetxJIaenOGg2BflNdYZPPOsVyw3XeCyLC
8t9SxduUah6X0ZBeHXUsknOTW/QIUiEbk0Lnh00ae1ik3arxyGypC5gD9dlZxzkMW8alfmXMdyBe
ZPCVEs0tXCl4MvQeu7c1+jqJj7QhlTuZd5BLd2dsI7RdeiJIbxhdYFiy4/FxE3hP5p7kqr11LSNf
lww3AyXkj+qG+nL7P7xuO5RLVt1kn9HYlmo4DR7h3i6gd0SmKrfp3SiljTvBZpSY4d4s+RO5SnYT
gPnw95ktIQdUMLBan9yVpH5jEqnLggBsNzrBv5zRh5+0ZAClW6S6taDJse4FoNd9MomP+FA3HP4t
DxQWWxsAmmG0vorJNwu3Hs/BHKA131tE6JF71N2zZ9OmrrnhN/oWci8YVgiRGVLij1J6tnb3TP//
8lJb2+j0GFizCS73N2DKHCmkKtBKrmLlbATnywc2dw5rmGNOe3TYofG+/eMSJ1smtWw3LQGSlppg
LfofaAEW6kFoXeFxtIc8AKKCK5gT7nOf0X3HVT51HfQJ40+xA/5kq7Xb9HVVGioieamA2Our/pNv
5C8zG/m6igvPyuhD3Y/+ISlYxN9ct+nzeSIPArozuDu95wMB+ESQaofnPWKeb8pOoS9/Vehp+LcI
9mYBXcwgI1ET7ifo0LI5z/fmZHJXrfrORtM8+cC2+hjUFVSpZLCa14sJua39vJcnWl1YZ6ZYS+fK
jwVY6XqkzNoCHfW/VNa5cxFJN4SRGdmAhIvcsYhSeyAgoooCH0ESucI5dPCJwCQsRbQERIS6judw
q3ILi4XCJCOjf+ScgkXzCC8x+b4l7/AQewNfL3KF6pqZlkCrqtO4INB7HR0swT4xkPXutkpmrR4n
vsKpUAj6KpvnNK8OCf1CRNb1MIxZHXxUi/WxU6AnmvdVO3yB3KW6F6UzYDWJ9n1fI1eQgWRgmE2m
RAHRT/FWMrxco/X1OaPkpaHml5SZlctKVstBTv2AyBP7xDdf41JLt7UtB2fdWjikoB9sW1i1VlQL
Xz1P2+hWXMybH6UVuRgClf7nCxVa6yw53WhBM3L1+uCJgKonpa/dKoE2NK7/KEe7SVbYd+p1VvvZ
d0ZTx/kiJ/HD2pP8HExHMWR40MUy+hVUiRwbcxaHj2wFrZwzQVk8n4yIQscPvtm3l+avBrpALHkB
p7tprlVKFFNQQQP1hnjE2Q8HpeSlybopXANjsxJ7sExUuU3rumjOeoXuA5Ew73x2s/T9oGXWnHo6
gXeCwttbOsT7WnGdcGsmLi1Oz0GZlt3bkhsnrfv18J4wLz7gaAjodLnJvVcLtmVxaWhkqLcVZN/W
3FBJMt51VZ5yl24qAKzn0r3n4PnEM/OTdjqIZxlQbVkErSvKiMWdhhDdz5TwcRYmD0pfOXagH0oA
BjAMBPjRIjFbnDj5t5M/CE91GJgyo/4tv8m2sLWHEzwbS6YfgyLw00oG/UZeyM35gbArIysJz8YS
pgmjsFjv+hk0z8lMh2JfazycnGb+dzee7on7QZscOHXiySCuArPS+djvu5Ijv7wpEjCnctKimTrk
aLy2jhyZKqaYHzLGdHeptWHqqMKIn7gPb19iT/S6EbP8WHbTJCGTcXSGTufl2f+AJPtrARaYllBy
lmK3Vpr5ZWoktdv+RNJRIY1cNkxSu54B7mxGoKiH1epGnP7ZqiovPkB/jkd9gXaXobiq4V+v0ycw
YPiPZOjkAoYArsKMhC1Ld200Vj63q7jVXdp2CJWCMQbUXi+UQ6xFkEDekLCd5vDEuq5ElVHTtBSK
kJryduCDCFZc69fQilODEOw9i2ySLJuPnWPtCcElg2donsi3KFxVwcM9lS5K4C/94FB/P6s8VbZm
m8PMeMLaHFsy9HbiIkQYYlLOPgIz4ZfC3w2Os1PX+lf/ELuA1WTbo6OB4WbdU6r9Th4UcMtln0k8
BY4vTJf84JKqct7GgthEGbPqoTpdaIv6dCLOqtbReaKlT9q6DcY/RhwtwzSWqvVdKR7zoIiKKMLX
6OZobmhyNT2j9D2F7JyUhYlpNLIAsoLjBqk+LNPCMMfmfeJ9NEUB3K7oZV0UFfcA+C4CWXwtEMmn
VCYGZ4+Qdsq5aJMvDmEf8eiIcmydpwpsBo3qMgyxXKG5wnDYKWPgKZkKiiuok7s+qMvbdR3iXn+l
oJHYBDPfNUKYFZKEf5FPOL3fwqJjR4KACLBV6ARPhw9yBDQbaW3nyICYMEDQS0RvDT6j+bFaOWkk
ic6WhmfMXQJy7e+ozfgsDk8kpXkwJ9ld5EP+CpXVLsAcnXwavdpnLKvpozEOZ3mrSons+SxE3rjR
WpFSldURQQ+zcfdsXgz/tNdAmHhu0MHUJHVvI5SOqpGqpULg6/kUhGkCzU+STnPNR/qEBpY+B3Q3
0dp1eXIYAiz+fXc8HufuXhwidSRpZcH6rAlaySS2cVBWFiORVaVbXYihlNRz1ZD1oe1jPk1/MJ/W
8LGnRM633sYyvyCJS/v9QMcuOysA2mTiO3X9O+Pkg/vZVEseISOq9REZGjaLEdWn8dxpwmblKDQ0
nRDwd0A7gy8rVauG7SQ89F9qV/xL5rJOO5akQt02Obkpoq40tyRk4guf/E7mcahFjF+oRF3xF3+w
kGW6DIPXJ7THQi5UmMFtA6OqukKgUpZvpEn5L++Xvq/3gCdy6vmawbmBa7fyzRjEioZDlD8sKN2x
0RxDuRTetdcb3CQuBOKL9ePUW6cCbLuN9pnJkRhzLEJz6eSi3CgNp21uRenUabkcV1o6rieWBqdO
wsEvNrJOjJQMwVjDkn8IRDMCbySRod/8mu/PHgt7RRjc0DX+RYQdXLI74aETleZw8IcSwqPnFgBF
A9j/N2rCoQ/+oQtlG8Z7EWqzu079on4R8tmLKQhh25CMffV9+oDXET6cNIqVWBCYWkn3niXlfaQq
m4DQ8tHVpZUceXErf97yAstXVKSGtK8eQfqorIvlilxghA3AJ4MoskSUgmnvcrMw1aI+i1WVT/Cx
Q+gUYdFtVcDUkcwvKxbu4M1Tg0axi4pnFXjO422ge+zc6BWj2h6pBvnScMHMLgA8SH+kzeLbuPNO
r6aik9MMVWlxDXxCHjaPYxjZ924bpJJfcPijkwkNfBCnwmmAARlBEb1CJxJDTQDcW2KVne46/195
bgiqfTaLtr0no2t7pky87Gr7pWfDNEfzaE6aTw+kxKNMsQ1HZdHE8iellu22/N/4v4bmBQmz6ZFS
eXW4xN7pu/AboMRwQSG1Fvy+bxZI4651BcZcOPCVv74x1+fIh7NhldZ3SHooDPNzYGH0X0PfdAXO
iK333YWtJDlIbv+vbiqhiVYb92DKymozkEEGwXDydvNLjl56W0eew2dVpmiQuDvbTtZaC/h3vkIK
f5tSH4SAjYg9EUkCaB5njD0/ALsKcO7x3dmgG4JSsDZe7G8CiSzJRkQXfp1RTNPAY5jinRaWibGe
Y6yLNkbohxzjmKCU9MjpaJLteglYZGOiXWsbSH/7Gr4THWuGdljEWXIB72puKwXcxrGEBEOEqXXz
43IA/GBwPcpeKZ+toJ2UxqXivYykcnSpz7eVFXLPh4p/pd/1rmfsvfgtGtr98tgp9YlShh2I24Fv
YHlzuEN+P7v6XJSbMTDcf2Z9kUCbINUlcRxuupKNH650Kks1GQsfdtJH/yNoAUfpjxIE9sHBJ28W
uKLohM8zZpOeUkCohziBJy8wuVvCG2ri5FKIcMOfCueTc7Ziq9OzX79W4W+WatUUWCb4BL0+rek7
seLFsurz4/WlmX/LZZ56fsm+l6dVUhzPguxNLyaDrgW2E7eFLnsfiTs4998rNdgE2UdDymJJwCLQ
XeP70PfOsiT8gCQ3e4PqlxcEa4lVuPfi8Jt0RZhRnPE/gM7B9cXGPVshXB8otWFYRN1Bi4gqjJtP
xUT3zwUDq81EnIi1ncd6Df+by6TRLD84X4xHQV9mOw+FWfhfkcG+z81UAjw/vKXB0oBy0tNpZUfI
8KgLOHlQxIscSb8iABz7fiHarxLTFWfD3g7yHLuiftt7t0HWKciK3SXmclumOWqN5BPbS3tV7nbM
1HopWEVNSpZt53pp+qjUWHCzouvDzK+ZCK6YTYtjAAuxC0kpDYsQSqaTdR1ih9E15Q8Wu2gS0Evt
/wyDYKn7L4n9xewpKPh+Pm5mKjcz/qO5cEi0dIghfbqM89tD5dQWxNcizOfVKdBWVaDnFsuhbku6
dOLtXQDu+iFQTxAkg7q+PlGuusECNSLlns0AnEs65kVlWmuAg1w0CUK795DASi2eS+1V0oUDUaMD
hva6BevPTgU4emp6bf5fLkdZeZSRt936Viqwb7RkbxpnhAuZqW4xQPguZdjMi/plgfFIX/8gZLX4
Qor6iy2uHUPwAH3IzFSbNnYAzvpLypVd0dMVULh5i6vWW2BvWRZ/BnRE0/vpOfyCN/9ymWeN17b4
yUNwX7HexjIkOyXmv/f9xpyquEm28ChBde2GHIQV9IIDlrvDF1VoJFiMhFkHq+jkw6SlDY/sDhSs
q6yH/b8sFRSYAp8+yD7AXQB7hpW9//qgDVX0EN+0fYxCK3ul8wXwYCBFSQDZZgtKrmKrpCL8cnO1
iFLsOhEgfNYTCQsEkx7ECOwCJVFmGqnnL1SjIj895nNdJRdoyl5GT9RvSmwC+uhwTZVZfnWu+qVV
clJeSq6JplQelHLKLvN6YVuXSclwaCK4kNNvvy7Q3UTICAaZOQcjNoTFXqnZ5fyLq6TMUrhRHl4r
30dTNX7HDGQLx/Nu0D0Lnbtv6vnpBLKL3Iuruc22ki7Skw3P/gxVE8DYgaVIvBu23a6tW3moxQe/
+BYfZWFu/ugPi3FGfz0RgxQXaZtqH/2vu7kqIBB0Ay6/1oAUQ06rrBDnYe4cbaTRt9UFoXhZKtqo
Qscj7OmB0UFA8eauLwITBr7FcKNg2P7nm4shqd0cUNXHOgzcrw6FRpcGldnJWOHK6dpJZb2V6Tw0
IhLEUzIofDHIs2JOv0KzbCSyuyv3AaRuVeliam5wbFSyu5CPdPs+wzFLZD2Vv/3d1hRUgtaGZc3t
dYCCRFCfWAC9wHX5VSzvGscTrwx2lTYDwn8veCdlv/d4H3zIsh7PMTrccopksAsFSEA5k5MvIWM2
E7ii77pIAlr0Mg6m8jAsztgPQ+BjHZamniAZjv8HRXJoztjiaR05y0zlSbMdOH+q+3xggWFfX7cv
A9oSyj/jfdIRZss7po5vBtvBCoGP3m3tRpJ0vCOl8WYbqS1C9WkTsMoWC/4AOKvkjcm7WAhYnBnI
hQgeVsm/g4Qb3i+RrTVYmgzMrTWAULX+eTVkwHJuiFN2MjC7q/maQLfWkp1+KeybtYNfvGEVvxH4
EkHTNnxJYxHkPjIh+QdH7XsflCwCIdgDAlT0PFh/qk2R0rgKXyeLR2y0ihCc2yZWr37kncHO01vI
RxDeFLgdl7iUqNnVTkbbkhPwgwbNOEMZUHzR8Sph2lLgXgQo9oPTnstP4EG5Cy4H95PkqtruHVM3
CaHJ1Xr3ollai0K9kiViL0nyB4eqPeJjT0SLh/j2NuolUYCmxbIKnGRAdNYKmYBTqlg+WvTq1s/j
bPrDee6OZD/S5fFjDzMaWgTe3eQcEycHZJ3Z8I3qvQZjzJSZWr90MxKDAPMj959irMOw8vSnRR3F
ix3jF9+nhYv2QN1lyw6qrZDKNDKJfBCiORoH5lkeLZ0IvGuu16WhlFbY/DSdIA8dYf+B7Z0n3xeU
E5V84oRpCutg0jX046JXAwxQxyoZ9n8posTjNxHmSX07iZNx7V3E6b0hCbNSMlW5U82KOC2udadC
HSdVLFUAsV4N0tkPJbANqTDDwjZvthLIYnprym8Yl0h35TrZlSVbFdAUUKY40wlLEHt5Giuy4hcy
7RzRHAykXGyhBy+ZjAFQu22DdCX56FLHbpUIdvc1fEAfkdHyhqhKpPGEs2YdfcR+hG5YwOto03Qr
XK5OSzcHIlLXdp6mLhqjoqlvCrDgmZNAYwIDt14fmHo67OVEGdBxdi70LLJt8VZPiaVuUsd3PHHB
2YgNaEH/zVnOE8Hn36atQKi7i55f4IWkHzEZtoGBzFGjzwlxnKBbn1ky8rsa/nSUkBg2tMRsDN3r
M32p4/Wx4XVTXMIEMPr0n0r9nqaL/j8s+fQw0Z+9NgZAyUUAsYLZJ9Um7+JXjgsKXfq75z0ydelj
773S9EMMwnOkWIgudB0X2rVObMnkyLbqth3N+nOr8hsdfdnyeUbq2QItCwzTkXB66Dpp4i/lAawJ
rSE1e60yPlSmambACFKyT45SQNd/OoV9c9CdI1/ALCxu1/NMPM0sK7lWAv33S4njXIuwx2o7YDD0
cSnQghGK01xQropsQIpxu/US5QS6v4gMGWvptcDQH2Z+A392NoS3R86fDtqYjjB69GHteS3kc4aY
BEpGl6LInnTnDEK5/9KJex96iKaAmZdv7orXrtS4dh1eJICD0OKJYIpAPGLy6OVK2SLeh3Ikim4v
txg5dLKqoK/BjuJo7Utn7jANYAmpP2QoTu5ligj1ZrvaoxOYbRwflAsg97wPCCH9xF2PKu/KxM72
F5zyCLyeAd7OyY3EB+3T1ELduZ0vDTS5s56yFGF5IlQeFKGaeDikMOVXY9Q981VjH7uerTh+CGqV
1YXDm0132fbfG8wPb8UOCMftkc0wNaCup3EuH5sfvZara8Or/aATFf5+OY54MbhdfagvknUz1eGk
ULrCsYrgFgl0WQjY3xGmUWozcgChaWiYRhBgw83ScEOm+w0yGfqn6XWeHF5xicfNi4x/yaP9Kxs/
MJv7pLI0f/XXn6xHP5YBgEFKFBDcbW5l5008CO2hBthw0rANe4STp4cIbsDgTBgRa9U3NAzMzGwS
y2WCtPwUS/ApfKDHgMJ8PmK38DKEzzT89F9+IGfkXQ4q0S+HXLsJMBhqZXUAtNtvj+eAG/TOSne+
PrLn4x/wbayS0M9GF0YfevyZdTijo9VXCjYp2NXZbbX7W4rISFSg0VYifoNeyH40c1xMCQiNfVT+
OTFNr9w5RRPR4eLdJyYPY/gdGnOruhG2M19slK21l4DtUXCsvNXYL3W2SCAJWzIA6AemNnEy16SG
2EPpriFqCoBpB7dmzNvfrpGr9MtzzW0j5fMb65TbrAnFLyLDdTwOvUFtGyGXTN6PjPc1r6q1GKDY
3qRLtnnqx2dBQd/lBx/ZIAg6qkY611WDUTP/YHpiidXlqTAUI4Sch4KasAQ6ZhuR4VKPD01o7E2m
L2uVhQD3u6Q4gLJUEBM+lfOQVAqcUEURBhujE3/YOvmW3eHI+FuBmU33DpSwsrL3ZPycTrp1zWr6
yWYjOfQLFHgh4ynGhwyFYrv/Z+ouL9ShjgHfCryd3aIwdt+avtVhBAJl/3Cfwu01BYyaVpv5XAB4
fyoAhENwk0uExLMhIqWLG6DGPu9P5zR/cL5/IcvqMxCxtp/nS4RqTbH34SHv43yoFCWAKmer+Fv7
+QjsmUXSKNu8tt31MgptglvFHYIxISNO14ORCZ5VkuZmK1lJkPBoa7Ft1fUgnzKtpAFwElDVM9rC
IK9BngnX0l63SvkphBmrkQlGh7g/0tStoB9rd0MIf1iLjo/59BPV52soRwLnIQX6WMVr8gf17po1
AZy1N0OClY3WzhPdaahs4EjIjITQ4nKd2Y6p2mUmvluvMVrLyFUzmVbqKHrnxOivlvyiAGgul/oi
U8cjUdLIZn/Rlu29ZP0cyd0KLaxsmV8C7nBVLaa04ALlGu3CzGAPCcUnNp1V+y1ntpkboCZHIb3w
jy1/hMKEemZFI7/Y6pIDd3EpITZy1MlNURGvtl24+0SIZdEv+jYrO/kjWaJmGIjx7MTx6li1C3h4
9i5a2cJ1MoJ3iyJq1mvKkgcME3/netpwxxOU+mzBrhJOdFCJN77uPA0JeZapMr1wIFDMrX0/HJls
75UVf46RBxZbnTHESdEbs0aSk8H5k27e50XpVqmx5nUNXHmi0Wc03grd11outN75XT3OH8agijXX
ECgrt47rc1rMXFq4z6OeGv08yXp2RGywkWUGl15s9+2j8t7dAz4v6y5T1dlszT7sFhhsATA3uUUf
pm8vXDtfqs9zLwF8QxAwB9Pnh+qK2cAepnUo9VOaPcH7S4zg8eXwP2cMhTFu60qz/Lmoe5h0y+GW
p1OXeD8Y0z4bklGFwJl/iNOEZ/CNhLe40BeqAKhJEUiQylIendS3Zus/HFu0sKzX/3DvV6xYBu8N
7x9R2rXGHgJRjHqsjikwjjfi4IM37H0Ylz4HxETT9KkrGtQuAq6WYU2M7xeL4JtqgkKc/WbQjw0j
hO3pnFelwC9dsGtazvLHfkVarOmfUQtFZ0G14588ZL3sH4JTBzSm9QNcjc/3Vtkfq/FQDEvirNxz
q98q+EiRMCNmwOrHdMNyiI3OdiG/eIaBVEEKhGthsGrZhzHQP1oKSWWeuKWyZEkibWVV2w/NM7s1
FGxvYXPCLY5FbaRSPnZYz6Irpaqhv4qkIm7S5e6AH+MriIEj+rsNUuDShSTNb+EERro0iQS3YIOq
B3sngGlChzR7A52H3M56bidC8oajeQuFokRriepSMZ8ofXNSRpF/ztKHYGpAa3WU84B7aB6kV3MP
ZaMEBckggKWAYHmhUeE9cKSZIJ4P99vRZknXDJWHaip07v4tAp+dbnjI29HiXlaWSXyea58Jqs36
OgRg3Ib11lM5O1teyYlHyFQ9rcG8vE8Bd1EoaAcFLibDTQPYRmWDhn/Wr35hj/tKYgt7bSzl53Pl
DIeoBJJbIDEP8HiFAGOpKJ3Ev3hv2sV9eaEV2tvZ0K7aJ8sBiCAN4aJfW4sGH+/WOUl1gqAKdqIs
WPhdWAetbtMFMeleFHKwqesxEvLWwnbyi7qfQ/VmxqMsNMFTnd/cS+ZnqS50Mxlw+F8nPh89KdEI
957Kjlix9A4GZMf3dyYpUCjVOJj/KHQbxAbF5gb3BSZLgfCZktTNVSrL82O1ZtQ24EW0qqDNqkhU
w54HCz7rjP0kKVP8mohskM/0Uprn1ZS3TO41EqeaLCuDmSr26do2Na8zqTvIqMxYZM4MpDRkuHco
WFXG5j1Szk+wakXqMuWJLB3Rp4MDfTXK6uHd6dMb4SV8I/m4ibxt1hRVTbIaj8BbA3w9zqJDhLj7
H/WNKR9cAkyb5kbh5SodBN/lHq+RD+RvWUUHYRa4V6CyNeYD7aX2vtM5PdoOjODDGZOZqns6sizz
HlZqQ8D0qNiCttwjuZDw+kuVlUimh6g1+1D1z4tEGDv4Q12ZCjmKiavj4/7U0VJ1o9O8FiI+Y6hJ
l9wxMqMMMPBASzO9Jo1RfH4bByQUTpxy2DYCR04efuU8/ZpZFkVk2oVpr6f9jxUcCjaVIF4cbvWQ
W81xaqri3gLvxq+5PCuYF3wpgJ/EIL6+H6Ru1cld8a/c/s42JwpneBHhVbfEAj8KM3RiuFSMlp9E
rMuplxKJIV4+wlmqcwM7xiKaKKMy2/FRSS1suvjMOeBwC6amiU3tlPk18A0tLVj0ejbBPZKpxHXI
a77m/xyPBInMFlMRzdcRre/gM9nGWZ0IQRH5mDpBagBNbJBTnXHfEbQHRHzyJVjhXfFvh9yJwtuu
jFSV2zYKrlj2ixYGlYOFJozqqx3t/bVW2G5n+xCv0k/mo5K330fAOK1T315voUiZreWPCoLVZ+Zn
5V5fuD1Nxx3uAdSsOOrHSXIQLy1K0qbJJ5dHn4b7DjtPtGC9/NicBLsBeBdpAYDSCmXtc5I9Lzcf
zhzy6oqmlUJnclG/HPlKzyfsDvKuuLUjwpvnYp9VqTqH8VkKJxAQpwDYaxI0rwDydgcvPwZ4xpQt
MopBsIqy0+VM1mEj3iEUuJ3ic29PR3Q8D7A5FWNWCgp6f3UxFtmecIEmo9uO8vk6uCcVSBs9nQv3
1FAYDCo4nYx9A9uf2Cn3tz5veWc5SDs0CJFRsvOqOsZD5epp6ZiUpyJ8jN7tfCMKh2G+nMwL059U
jI2KcdsLGoXlQbbzUs5+ee/GCbgBobL0PiQXx9AivKFLsZKhBAzn9jJGxi4CNlwSTOhmDNdF2vM3
yddieTn20GkoHOfrmGEbc2zOFA4bsdkNFBXbKeC7nG1/etFn7c0S1j8daDwd6mA1t4pJe8m+RRd5
lUNunPTUlFPdp5T+4HjBoYG0mTJDb03JoJq4isShIINqirFgT3svfzPb0QxOpJjz6dWQ291I7svx
4mcctA2h0/s7nhA+DPn7ctYHaVNtXMVziIVJOqp2CJltzd+kokdQDqHnOAINBUF5ypkRsvBB+DL7
pYHFKwZicfdSTaEiVHQU/f6e64gju2L7V6+tmYQUXH59mV9EXZeHpkTOC0R3pKZZ7V22Lw0ulZzp
dW4OmtH86Vu9jHMkSwM5FwUvOlUvl3aEUSE6d88pJAnqn8BEoNKkPXDYQKEmXUpVXKk60xH33CWP
hyRRJQIA5B0I0lgbLS83cJfcgKtM1bOgZe/qEQDIvnpTs5JOskoFtGXQhMlibHPttwrEkJJlbd48
gWnOnr6+uw/Ed0MJg6L8yAoF0LaGE13Eg5MJYDQW1kOnEGzNSnkIKRRVmvK5axamaTtVpyApkctD
Ln0wjMaKmEqKt7TnT4qw9wuGXliqyngU98jvPkCyx9UGP9pgL252FeT3mBC6ZcNAXUwMGrFsc6gB
xD8q1hPR6OXtz+cJzjW4pzSi6RzLLfZXRt/ViXgGjoNi5l1xvV2zrYbEGb3eOmkfkHLZnvjth4CZ
mFSolfMxvBqv/mw5SKNbJybz7jlJDJB38revTaMxrxE8CNwlhQqTD2KZdALUHrc82zmie4qFH3nh
5thwwsvAwG2+9s0+4YyJoySokMBOj9mgu6V94xu8liq8X+wXZk9cTa+cfz4WcFNxU6JCsBwhyHfs
7wOXVx+pKvl+e5BvrwPBElBdK/NadThZGiD1ewL1F7nBPh8OT0pvI2WtHihlNlxbdsJwE/KO6/oL
2B1bbYkmmwz46b+sggDs9QWogNpZ5CSbQA9tw4Nz7Rm6ExeNgfk940KE73PtzBjWM/hgXscS5Z7v
w/s9IOi0lQXA7NFrRShCk250RmypG7loBNQboYsZvHe1402tOlItyHfFWg+TakB8TouGp3a1g/4l
e96yNKXoiUWeM98pYsHzneLD5lPog4Tp9GVAM8FR8RVVwFq9++YBApavQgXtbMjvxJfkyS9eBBcT
qLGisuhN7IrlnzqOlr6iq1Au5p7ZaRUe2HBlhS2rCZrb5ELQqvCJFQe5PXz1lEyR6u1nta64kzJG
Y6wrQw9bkbxydjYksHAuHLImkz/vQ8ZcuLAsxEMZTr2rn1VvnSwVs7lvd3atxBYow1z3etvfVAr6
xbR4dfoxs80fsWd3bMT75OEuQ0kxujeSvlV9tk4+G6wvrUBYOmdoPHkhg6tAQm6C3XUhe+jTQXEX
aKfP3Cy+nDbAXUdw8S3zwyugiT385qeGrFQFNe2FDiFWxdvG48XbFRRzOjdA8b+ANLiG+ZP6f+7F
+69scVRiFKxloOqcnTDBmUbBSCApdzSHf1Lfn9C0kRMlr2bwHVhcoerHmty1yuhIqcxNGw78WHIB
+xmNPIG5NR3OKhCbO3boTNmbwNS2STL+T+v8Vm98DMbJICHHFkZIKoUdqXvQEBBi4lzCZq6+KTNA
59w+bOSzKX/MUDut1fa9a+xrLSQ6fY8cA6fD/BBahETqKE4ceUTcwx2QO0p/NoucWDDkOeEgmeSh
T71VoTOTwvrPJB25k82tbHyhwEYYN2JIDkmgcy8pttMRIgEGTrENXqkO8MyZPLef6aswdBp95D6M
VNgo9jOYOQ4Ae81Q7hoK5BKxnetJi/rzrpSuuJ8uzDaGbLoC0Msunc8LhdCHSVSkmt4HcEx7YjeT
Q7hUegb+//tvBVA1HaSO9G+btPMY5NT8LZNN207f9F/mXpJuLrkKjHvAAY/UM7Zwpb5Fo2VbZdYq
jgakqNkTEfs0gI5QZhxpyUO/1JxU+ex1LoEuY5QPoE8To8hUxMhEAXTK0/G84agtZkBouaNCF5Uh
0kucrxEdlELGU8Ca8HsDfP6CpmorRrUATzv0KJzDFo8LrmFopuPUYF+aSgiWbVewfYKWg9zTjtgL
QzVsdTHrwitH5IiZq3g59WAUN3z7WI50PXgtFsECyChKhOtaVt7OLkBMWYNW5zBaSlSIKaem1TRM
tDiMZLCLMafB1InKAO13d4VyDufBicr2zydSIjFkcmXTcP3h01Bq2SIEseYQts1QFxtdtsjPqOWK
0O4azmdfqIZuEziGavScstuSTjU9cud/9HqEPDc+SlE4rrSuiXudgil2QBVdyaoqFSpxUZOByp+6
cpoC33g3eJ8fl9P4Kwm0HawCjP49Av2CV0Fdo7OK1DcgOkyxNGFzIl24+WvK1w5jcBxtN6G5g8yx
Hh7HUpZYjYGgSozaGEPLBFUgZDpaYvfZUj3BKsFX2wG7sTM1WHceh+1SGuouGKQ+XHRWImBR3/fd
E0whkYTYCzqQfJUjInzG+mrMGsc8HxHrVmb56PMPym/MYJ1N9frGyjjgF7S+eezGRkdYCeuC93N+
531JrpbEUHWoJYrrks4ZFGVbq8fRRxQvPvk4IY1gGCtDtrzXmqOjugRYOzYgP/UuGLnnGlaDtgFx
a5QdL3L/XDyfb8vKWVcxjnPqNH0AzSbl3FcofpNTB3y94GjR04moPkqs71W3gphgsCu3zWw2ZRG2
VSUZpY0UrXKOqvpse4qtQHUd0spoPXvNz37cp/N2x9FLmj+zkFzSYCwoF/tzEMoalW/g5YeDUxmn
dUeLzrIXK5UT7iZT4iNRviuFvc94Uj2HN27/VdsHaBtvKP0eBGn0D/aBaKtq8Xrt7c/Ti/C93Wx9
e98z9ypwnYKHtQkay+5nauR71Bs5Snyf/mDh0lnTuBjZGczwWV46n9PkEDKuv+NWmKeu8qHGowcw
GBJ/r+IOKhjrQfsNJj3pTQ4KkDYUnm8365K4C4Y9FTsEbp8ormyBf7wDez+JK5dp+cFmyMvG/ZSq
WDhpSjTFc7LXqHo6lhWUZO3WZjAETiuS6qFuBOtGMuHgUkptZO1QJtY362AwglU7VMJfE3MosKpa
TCmbpGekeT03eIAnbMbECMZ2kc2F79lVPqfwipzZ4naHV6icVPo/JqYhP38cSSy8WYdskyRPY1LM
EpS4zH+2aUE/3fpF1INUynsnH+jPRDP2fec31Yce12HbA5YLyKE1Ab/ZqG2qp5po+FOa1a+Lgb21
Q913Lj93RoRSw/40aaJBQAddIqKrvHVs1DYP6aTo7KQj8hbV6os44ereJJQKl+svLc93cHjchML9
MclxDee8QFgScBB2o6Hswjdk4WwZS6xeotmX/wmn+AKUC3ObHp6eLzLShO98kbeF7JJYIhdysVe1
G+5+few75sbdhwhJI6PjI/HEMWB7tW0onKyBeItHUlNfiqS0FGqFAWP+CkmeQMx/Eab67KJNxoXW
B9/uA2k6pZvoceTvsgsgrLte/i6DIiC+nd+QYAjU5oQIBlRtmzzU42s7Sl1t8rEs1zfxARIa/buE
CxSf0Vgc/L8UQ+TGdWvppTg6QRbciBfDciPGq71PDgDkFuAK7sCVhJDESeMAHaSTB1WWD7083LqE
KyGe+ECrNvXyErRFGUdd7yeu+qQDqQKJJG02+VVDYEyocHJP6wrirUTmD6oRbS3wR2dKsb9Q5n/a
Bi+36W6Miaxkdrv40r8N6MWcMDpg33iL4k0v4MuYHXmpx1ZoOa6jcEmzzz8wvyHaX3W3aLsbjlOy
9roRuUGnf+48S+FGcRIffZb5SLSOEOZubPICx00OtvvFhkxp8DyKwfe1WTm8e+AY+3azjyB5lP3o
2xcgZzhGR3QaUDyvUw9m1jWCjytqpo125GdU3xACliNEApG6HWkv3nB8ChuFhG3VxvnHN8K7FP9s
Nkdo+7Ao8gPPNi6uF6q898yiYKXh/hzfWeaPDyUY77cUhlGUUE/7jSYNsIRN7slWqI79aDCHkSf5
Goeb+rMaFlfhdMJM64sCZqe6UfghHXvYKqTCGW5rg4MEb+VwM56I/eNwD5ATAqWWmyWNyLbLNtib
pikrpQsB7wxqHgehB6IClf+dwGL4+s6B+ZUP3gwl1ttL6dUC/p97/KTHMM9/4Wy7OKEJdtsJOGR+
/j0lZBylhWCjZ4SFsqKqDJSU7kH0AYuG1s7qdemiIjFwHzsG3T+9mDsYdU8jl1GoarObBuYVjvuX
SXNkg3m4F/l98+91AOvKHDs2f0WM8dW+Tsq5pGTOQ8lUJPtd7wodQOPm/34Aumpuga/iVhmn2U9E
yWqIf3SnkfAbOkNuj0/vX402KC9wywvCiXIKVVbCYi4Eji5FDKSpfwXYrg2DvBNzTznN/T0Cdnw4
OrWqAgsMnuuEpxBpLNalvbClvc/zye1E/rRPp83s8Q+eu3eMsE7ORTCUVC6zGO2nvqlnvl9n6Pv7
9xPigBOSjktrAjl7aELxZA5NzS9PhQ/9CFa8/118cuga07aX2g8ffp/7QtioEizJKwZMeIu7KLG5
9TwUilYxNaRpHF2qmAbWo6TsONsS7Ubeh6M/KVz41KE4o1GZMrbdPVWbn6hmp9fvui6XchhXqpxF
8HZvGZRdDYlveYxIV1a0rYIvsPppKkHlu9tJa9qUhKjnAPYOixCgz92mms0Fa/pb/cp3FJ0o/6JT
Il0FtUAJvzkxnw4tJuu7vR6MEjdL2w6tcrkXk4Ja1wMqkERtt28s7whzmTF9SfCUKVEa+k48r1UH
FKrzi04/e0Bx14cNlh9ddHxN/17BAQRYY0CAsSmz81Bs7AMX7nkFlA8IawoQaq3Chx/8QWc0a2Cb
EOhQgutbEbpY54+xi/Z+1ImHQMPZvA81rn6oE/046jlv/VfAfbIzvse70zG+C3c/PCrsU3H0mzM0
ge7bg+KeUcI99Hlbls6QByOBjqRZoxiHjp2QF5jS7ret9/sgN74JOviKhgxgnMnRyQ3nhUDrWoWC
BaUocaHEIDoyD5FPkad0U9rEM574QPIJf9Bp5RL0SiDj+6BHAJZPAChGOXN8O3o5TYVOvNsUPz/e
zBuXqtOi4dCvpppoff0uR/FsAXLe76TmwEv6dSocRCFZfP+IuO9IIjHDiT2CE3BjmubugVew3ECc
j5bIi5ULpgoLioksUMkI7X/LH7+zz28c6LRPqyh0Rb++gEt2fnC31A8Ru1bS1mv1vNlmBy1bASbC
YdmutJ1/l6PRFG36JcM1oyXAzXmHCFxwSAloZmMj2oY67HDJQrAfO2HwXbu2T07gE6fRohLwsvqS
FBKzcwqsGJH1M/M0fONakUiIvyMXDmY4Uq+QNeAKVTu+ZYzlrWF4kf9JHhSf4vVm3mARNCDvNpp2
FpaJToaxTHoEuhW+MKpkhociHA5jfIvTn0LbStie/vrxHJS45eT18vHlWXDH0W5s3wtzZFTZxnpD
2KgWiduYzlg2yp0r5H6hnB9tT6UdJk9lKD4Pwj87DfFFFEbrIlIHtbMRflizwYY0AftyvibBhv73
Ic829EhPvoaZLKikqr+od3sNhF1kGANjS1Vzg6eIJ1YIApJVOV91nNoHizI2fmYSygSGu2Qchv82
shUwgIKkIyvN1pCEyxRj9pnw7NVxwvc6Gtmd1ldCH0VeS0elsn/dPoPBOvBewlzraTn8czHE4wTr
3ndrwUElWGKvmBbImsxW7WcQjsk8/5YVGqTu6fqtYI005GUDRk9cvWtmjCuKkHnUFlys16+XEJW+
SnACZC+84wY4GJEvAm42HOOBkZBkbxIOl0e0Z1l80lc9xyYsaV0gpTNQpj0lsR1C7aJGsxQrgE1R
gKwCZqnMnqLACMf9/PU+14gdVha2bAmCP1qkdNfJkkeFvwY2eYUqhSYRkJDhvWdRlW4diGEIuMYU
05N/WoWrgk7fqwqtUFY7d+YYo/uqifMzEqFCEfYaQDdOTAZKAZBWtV4DqBAH6HNt9UMTNKxjN3WU
doebucPlAkHBcLNHsc6M4L835ecbDrBbyN+1zfPIO4Lmlh1/Y/6ieF5LYtjGytnzYTzI8oUGyxqu
OTlMuO6PIn987zelb61n4zgmldgOEqZA61G3A2pX4Z25Zf231yj5Cj72/Twi/Tom1MV9XwlsmiXp
Qc2ZKyAseXf3oKA/5UcjjEelgTqSU1U1Y/myFcfsrr50gTjSc2F6ZR6X7+3VJzhCFdUhCsNSu3Jb
VMc9LNsAvhk1KYjhdxzK2Gt/ZPuI6nkViUuHq3Y5qu3qMCmU3bDA97ju4IDPNKWkHNS6+vfwSa/4
0HD9xcsDxgGdZi2FTpHuBAGigCLikRRqZYw5wCTa9jnhK57JD8ASc5Xux1ZRtTR+QbtrjKGNb0Ct
bNkvATq6j7KpsyGLrPIPCjyTzxC4n4yQn1FGEvhsZVTijq9lt8OR0SkIrLXezwZiEWV+lZgCOGUg
CHnLOAdGetoOtICxzjJVwjgdYfZxaxWfTpPDNfKBCLP8bBd8ejtb1/ViKYFew00kk5ezKbrW1+48
IDbFSWQBp8f3AbiKoeEwBSDfykbZUZB9Yd31cyzdcQ1ROHRGgZo7l0YB/GoYzds0hMYSiCE/igAe
Giz3g3UziiCKnSj01/GwXlzcbQBkigz1YrO3NyCe8RGbkG1Y3xfgham71giuX86IlLOQ9rXOz1B4
m6ggAkhAmXhQdFpiwd0LdZj/qsqlM36Z2GCCj8/qddvob7TKbQAd/KGwuHW7cCIc8FzK7YRAt6Q1
U135cbcepQ4wUf5DQo7oz7SYn47GQXANpL1E2LqJ25sNIxKu8sVAMsoIQfWzL69XEvnlrg8e6+YZ
ypk7ulY7K2orFcR7Iq0UA+XS20Er0ZM0kwXezF6kH4uzLo3fKTQdooRWKFWowYAQT21QflrKCJRl
Q5XCCftVkJ6EohvmY8wdAbb8sRunpnQhdpXZQTefFbEjqePeVB1kGs9Dh6vzsCMN6AX1twtefJj7
O0qHn34QeaUk1342nJBt3a/zva5HIm4YDtUBoG3+bOJDjylbEWs3cbOSQATPoqAwx8BYDjIaSN+t
eLeYT8u94Rm3ZB8nyGOai62rJXXtAn1i8tUX5IFjhyTUph8jtCOm8meKtAb3+P4mNsRJGirhhWeM
l3Ljr+Q5pR9QmXru2QSWmqDMeFdJXpPAaX0Hfw2BRrsahtPge+zSVWuviY7Z4NXPvN2ohzjBcIYd
2+YbVsrKlTsv1I10huafDvGlw0tB7dYatGdu1zWs3kxarbx+IsxREbcDZIZB5dvIAwlncBEaO0nB
oQ+ZGMxkmhJlLgdwtRyPzjssLlsPOO0UMCmVgvpKEcUucMyEh1zyJ94k+/OJBKukAOCwk8BbjrVX
bidSH+OaXBWkxNgcGSIPvTis/siw9TtiAKNr6HxUjXeFmTgpImxfgq+02nZf5fQaBNv1zNUk7m1I
z6XQ7u4eVdFPJBe07ctqCh2TqrrSkYxqxntrEL32FoOo3sV3j6A9rbLOQ6A3wpS79BcxA3+miqzB
PdZS6srba2tkQn0u9BHhx5W4ySlQt5yJI8ELrq0Ljixj8xgpbIQbIRJxId+fAf0UrFsJ44rs5JLm
4I6gUKRnoFpmRo8SLJEoFntHhSEOHMmMQ9ENeDINdlskigH5I3w383zMlEN2PPDhs3aCLuMOiQQr
9JmSenoeg9P8/pA37lc0LDulUs06/o1KRz76equDtd7JdAXYkAoVCaXUinOuMi/70RzHD4+mtkZ0
dHEF6UUNrEdhIgd/Gml/lZaO2+S5qxlkWR1EJ63btoOKrIEfxGNi7kQpa0OaQ+Vb22KUMx9JOofg
TiJix+vnR3yaxV8k6+nDzMs+xM4BI0uTNH/cotgxTNNalCgOsiwHwRZ1URujsOiYbYWTyASVoFTm
rFnVzUHDOUo+CIaPYkOsWnxyACAIOzH6qrHaSv3hikTtFVs8CiypAlYStUXpyAD81w7QwAIJZ7iL
vFSKuWyfj1l31jbJoQONE732ZWwsSXA4IrjG+BFWBuw4XXUO6+qk+5ztP52FRdh1f22Vw2whoM9n
b2o8Z3iQ3yPWrJSFHKjhUGMWkOnWlCRdTgAjCaODj6T+vlplQB4KKuVfBOsSPupq/9cmVQx0Uzve
aK5n5rBJEKkYV74xR3Gbaec5X+SWW2V7FjfvhrhXmvMy97YxPLFiM/+fu4ViJcC3hcRpHqcfEA2R
XJZHkR9BCF0DBthWB9vUBzHSsoBYQ/b0jA2eWKjge0V5swEUx1VJ7XCxqNXe3W9oYcvpeRdPDWH8
065dBWjcywPHIRRtmBHiZjkPSWyxxXy+8RyltXTCmfpAXcT7vQ9uPFuUGndG9m8yDbF37OFsjC6S
E19+iNRl340kZ1o9GSiVxCWo02KS1E8PJ3rHmuNy9UzkM97h+9Si5f4DOx8/dzv8u3Df+RVluR1C
nNH4Lg5ZBiSmIkQqpnn7SF5kgQmPwoz+/FtPOuNXgxpVYYdNwLVfljXuZ0gR0Q/X+BZL1/ruQpJ0
qgDUgdLfd5CB2O9vAbAWw0DMpbc+xEy/83u3+v29T3p4+gfJ/FzUEIrbtIsPDfF2RI3ej0ejHdA4
N6Me/Dx64AxGwGE1tV1iEsYuDXPps38kSnCwTe8p+sq1yvaFPd2UjUgoUiZAIL5l7dFEDzhf6AAN
3qKctNI2V67/KIk7EkG9FF+9eoOUIuMMvZYa+Zwoyh7MiPoAklkSidLNV8GQQiFD99V/9OulizBm
gnMvIZUYJy07YCTh9idxYM1MLAJnjMhykKC7TMC015FSIz9bo65Ah+IuUwbrMJL4unoeHqNXKqEK
X+9y5c8G8zHHA8iB1MvntLx0ZpRVVfwXdXTz+BltOmYhLXrEDt6sN5GQHwq5jJqK8h6lcx+ZUQ8/
4kYFisZvIg63bpR+U/p3VICYr9MagBp03azHyNP2/HuE38es7t3O0dHl1awb2n+jGAOuFOv0hd5B
yHoLamhbujbjK2Xo/gJiYJCSznvIKdnY4azbwgz390TxWE8F4N2OugZbbTYkPPo3EzkOORTO00oJ
+bnxMl2hIyoQnq/XdSuNEZMXpA2KiQSi9yO+4YxUNNRWK0ys/gRxuvSpgD1UXGHQXO4gyGio9Dpn
fZAvPYZDqK7+pHR10F0EugBhjDyzdqV01dxcX77r/HMLiuGaXj0oQmWnuTp2+71iqr9Tv1D3TXRw
TLkDnfH/ZWZYnrftflh3z8YSRPKWDMJLY/+nAf1IYt3Wz8V8xlEBeb2T6cJH6xRXH15x3yRq9E33
88rFpyfaewI7gN9E5mTi3qcgEYLu201qLekYATKpcXUu841OkQpm+MehP9e1N6TKRStGDrPkc6ZZ
Silp0l3u4TdZ6GGisMq4lllX3kgSDWS/vMdiBuFB4T+WtKgTviK0JKbAXgRxwrXbXuMDfJs7Yhy4
y5Y0VoXlDhbYf0FN/JgJiKHc1Un/9KxcNEloY0FZIKQJsq7bMuvc8ZhEmgaEdZI8mYOSF8QbwjSw
K7VdlMDyyFPGbK/unmrmOQgGjGvRJEdRrZb5L1pskDDw6Amo/n4mX/04BRQqCjLkMa+S6vNbE/Wt
fsliYXV143PNRArjom6J2BfYuiCrpzeDGC5YJjHWAzPgsizHqglBdgUb1cyHj+5lLajK299jivKx
MRVSAVqucut41K6wDJchK35+5eE4pWJllt1d+ZK3mYQ5fsa5YLEFTSUpLaJH94DHKdlXTWxuWNmS
lcQ5OyvsHpQ5ti0HswwsI5DAhoiRkM89VQh0g7l+DQLbaKxTUyKbmQPd71gZ1fgz/0K5buyV5S2+
hOIDY511lD/OH1OUXZyTQjF2R+sb2e/unozvjM4aDC2p4A0ba5kxhKvLNtzffDpOCFCUTzD01tDQ
n4PMAI/12mKE3VR39OPLqQk1fyXTafETL49bc5cV0enY99CqbfOvy1hmT++PL+xYNHFL5negkE0Y
Iz8a8rVo00r7uWZKc/brs2iAZ1pbNdvdALDWKWtGeZcwJHiXLOfvqrN3N3oBH60uXqzS2icZrrZ7
d0zOfqozSqtJ6GuTaQDemBwcm3+UXQoltwXCTdqvj/Jso9bAgRvb/ta9Iss9zc1Qf+QoE+HcXW/r
hOpG0r3VQJI4rra2iOgV5fRYSWHb9p1zKXx0qLdVL25HqFA4ICVlH0JVG3pT+dlKKsoVR266OKQD
lgeXRRbftWgKi2MuZaAYII1OiTlph07v0zr7PQ8sr+lqZrhX1GuQLdeVxBRbaPNdSn8sF651JHvG
jGjPAMis6CZzfDSHIOaNRIFrBQs2NAWpX3f4D0usy2c2uqaDiCt9XO+p73fZnb/tZWtVrps26SCA
6oYM+PaUy3K2tUJZIwA+IXCAdzlDgf/YNqY/fL3BD9S1xIlJa6f+PXvR4BKnUgRnuWJWNu4tk1zf
J9giPqmZCIVrodQKxPuLGvrqmhaR6S9xX/Qfph3R4thOZZtIqpASuILc5HUOJOb+ay4k/k6kV8V/
xF+13o58QIzCoeoZC2JIEnLJhXr4tKhILzaUYu1pqttelGkFqTfnznJSBAJp7lU00oDVGrWKoPLF
u0WwV78aIu0EJZMb9ljnImjznAy2tRlLxdo/w0PAEqI3NiGPnORWGg8dyh26I7BQlxKmrw+vWsjo
LiygJpy8Nk4LGwvPxWJfk4Glcrok1EQ0kElb/mSbTSmkrMwX383IPzp8nEagxVJQmzzpneiLef8n
5IqNmnibgViS57EWHABWwUb832qJ3OY5ZgveJHf41Cx2IG2Ta/67+KhDqK+Cf8IA6xPwbYYu7nrh
YU/uvn1jGhp0GCU4tEsq8I8kcbB+vFK20hgleX4GfqEhIpiABHheYSed8Jk40KMEs9Ckwd/eMzgP
rlPOn0mY+NqO1XKlHDQUQITOlGUMYAPJSUgwlT1Fd0xkmbL1dRghMcyn9y4bw1rNEOpJ528fWUrM
CyuNikfubQpTSbL2dunnskQFFzzRrCJXkJB9CPg8tNCHKsBOHZGUhgwea3/H8wMV8U0aVhpZAxEX
AW/IrJiriv/3457n9PLazicNq/wZ1zQFYXOJIsMzsFK+iDCp+a5c7uOtXD12sCJ7iHskTOy1CUMh
2Fx+59VgLqWdbRsM92S6uhb3WSCgqbrVl6R6KxUjivbXMzzMH0nIPq16kSO+uMoYXBwT2WeWFk8m
rGiWxY2ZPkNZIOIKJ2iYgI/RUBJv5MIWbPNj5kRk7gxN+D/fKQnwEbuoZah4LmEUmSsg2L5J2yHr
v3zO4P4t9nAAe2O/8usmUMx561p5zuB86oOXBTEUwEXpInfxJXWswemFp/xKc73q8t6Nixlbiuh0
pK6+qYEtcERmiTmjr+ByJ0iEMY/XlN30Y8SeleuyVYmsxwaDQgoxgEGZ8yDMtrgkY6Ijz9Vt08mM
VIcZ/F1CH/P7nrmvrVVrZPMWQVGxDIK9Wjb1lZzkC3ZO9wchV1W8H5VQZWTF3GkkdBQpWgIIpoY3
9yqSnMfkzjO7NFH7HpS+l72Xx56dI0/dvfHPej7MSWfeX0swL9sXZ2pmFAJNWQuQHQsPdtCpQBNS
CGqMKMETKg0ZfG1OzZNOLgVR0pL1bSUYTILfIrBnNY8UZlFAb9Rd8EEHfrzPkmLX2AiOV/kvXFmO
xwDUCwXtmITfeCow76A2sZVaI7X40i9BlvnFsyxPYM6o20WvyAV2A++Q7tc3yzXitbrlMO3VSfyv
2EiHk+8B8yFHFTYosblTmYf6K+PVLtJbuErbADlls7I10XmWuGHTHo78fDWRK81RAbrjPYU8oQAT
31+f5FKx0SUzs5cTk3f0cx/PAw0cBbMMPq9zcliq4i+mbDO+3LxlqZZZaGjvjgeuyDSZkDXHWy7Z
/AGH8tBx8nh7DsgjWWZzvKvq+OKZMftt90sYwqam+oW+NcB0AiyOWn5OV3DRB5rT0BcFomU/akIt
gusnNlHRal9fY36RxqcNDwmH9eUhR2RpzuH1/K35f7pRRQxib4qc4nTJbvP/lKpb4epJTmBdJWpZ
JctRtbGjlX3mrq0yfTWUkoe/ML50hSNcEsRH3MfI4KL7UlJRGAW+IJim+xo7XdmEggFRvAS5yYDK
y3p5SpYQywZGm2bKC5NM7m9ZClS6To09emG8lkhRS2SMc4d3D0cb3BfL8mXxqRwVMO74crHDN/g5
b9hFN58xp4EKoXWho/mrNX8sIT2Rr7hD2h5BqT00T4uTfgr1P7qgUZKLxtldo9zdraJLyBKe5BEM
mAzC0wO2cyvb/NFHwHYsVJIpThgQtVi7Qynyzff4LGV8PVK62Y3dNF5ZSV4kL7/R1RtH7yjEFdIK
sgDHCDg7TGgYFqn50Qfl/63piHZm/PIbIW4aGCx72UDctjKe4K8xFZVIZKrI+bx+6WsahEf/Ji2a
Wv172osr7h+0J6CBj0m+bMi/QsSoUf6XB5TLunzbpDWgV+YrgcMUc/dR7llUi/5uokRjTKf/BjDf
CmzeE9GCulUsohphAlxEr7K/xvpMSgXSlWZyOkgAB+6Z3AJNUkdXrE8VsgusHS12JRhV2bJpaatN
PkD7aWzj6Pa/U/YgCbyTXX4MsLszj1A1UyJJAV0IxwSgvhIhX24jaFwx8U9i4t3ujgXFoxEz5qU1
CyXM1uw7aVjH60Q8jgZag/toJtfymzQX+T4stUPR/wb+vn6dr8FH7kxMJTPlwLlHTRN4c2D07xnr
UaxWf1iasgOJkmm06VDIc6mRKKFC2NCwpfJCVnLKiuUgV2zQNXfIF8Y7pD+oP15Ss0qZ6Lnp+Bq/
BsITSFKH/vAlPMoWu+/03wc6KF/6ylA5Pf/Bi9vCWqJArad36fv/A5pBrvMV9q2gsv/7lo94Aogj
EXyAPDu4cZOzcFqe9TJ48HTERP1sfp8UW+rZCUkFXYxudoRSSSCgpDk77fvwnIt8STnY9cs4963s
6szYowP140bt+qnAyk1yrUxUwYbdeBRcZ7V884TMXArQR0EOVxkVfJ/V7pxA1soi2Q/dCQo/P8xq
BDSfls3yMGRYpHc8V6Eh9fp0P+WFk/RWwMoxaik+ndMNsGmPGXwumS9iq0xs5DXaSZ7Y37mtrPlG
bf/eAmAwaejKa19YOUIzUp12tdihC07y+nejXUCImATML2P3T43meQZerNJMPktB0HSK7l9EZeaY
Wbxwao36Gv/xgZmG/GcbNg/7Tp3HWO6U00XZ1o3rhctuJXneBxI7dkAsYhdx/2QmXXDNl01F5eT+
eksXBfXzxo0kOoCJFTe4DAjOTayToWQTADCaL7cMWNsJLVGwhP6CTzzoIF0jZZ6bX0MXkIy3TNSP
LxhzDxXUnrSztqTDWE/pxoHPPdKwSIBPHcvBO67l1sMM3te3tzDb647rneImyPohZIsQOSTgjHDo
s9QrvJi7jLak3shhQIT6/nh+pxLdCZN9ZNyPHz6z5WZrlxv89I9bryALSW/JI875ICVpiSehBIGE
vJLxsG0WDIp0+BSGe4wM9jnT0yKhGfA4XlqSOFPB2jZvndvdvUZURjuV8onwYOJIG0zE3G0R4jlS
Y3SqCiSWlKqjLUnJ5W8nY6a48b1Hs5jdHX/S05zlUQWaRRut8cTCQb3TiYY/EcRteJ5IoxbIU3Rs
daksjc9KXEgiQmqVZQU+Mj76MRpZWydDpTQCxQswSqGFbdwas9Op0+39YFcgrCOd2K3s7P+0onAM
nD0BtJwF1VBH0QK2lfB5CG8+lW0AZZoLYSaQFcsxMTZrpTSrD4rOEAlH2zmJPtLd3x1E0fl8U+Ip
+xD5iotMNE9u6xM3BXOvygjOGBHJo/lSIBxd4d4OXlivxYKM4qTfsjyFyTRsrOD0OCyzW/Ncp03C
fSItSz/RR5UJ8l7lYLQGhzQAkSvpk+pi4TNoLSKLZH2Dmu3AVGSjF/wEJe927n340ngCpbtQ8GO0
I04ftzbctPvw5bK4QHhN51Fo9SCp+k77bJI3UAD7GRJildLvU9quBmuadhYvvmO7hSBVgDhiktOC
f/7DyqQey5H1owfFHd7vDZ4SD7Z/fdZ2qUepB62d4UED7U4U8e0ahbN6BBPfMlbZm6BUurMfDSgQ
Q83MIN4BNjBiO+xUjXFclF/maxiGT7ydnLh9lb6skMJIxkn/ps+8WYiYbqZHW24xzaS7pf+UBnLH
MuHMym38u67T3myW8lSKYSiow3JiUxZFnlQ61Mov9CdbJodGNHpfhpvNiQtOqYK4Z6c+Zoh3OZ0j
BP6mKBnGBzuKWVur6G+eV0s07Edz8ycyhqkO67DfKKqo1emK2BeIz2sPM5aLvN3pmgXJlQ1Ff+Dn
IHToZUDMPdMKov0SAqnQRRh9eaPs36F72+UWRyg+R1bdj5cgHJfZGWKKHAhAzDB9R9FQOyL55Rd/
TdlT0G7MgI8kpAYlW/IN3vn7TTdjSPCzS761ZYxJerbxrf8XIoo4yRBq+i+hXUIUL1Gm8GgqJAk+
ux8G6FiDAp5jRq8dOfqk/sbrmyPfP5IkNeh9Ai1nH5kzvRpVMt9tm1dUQgfoELV81SJLItxCF0QS
edBlprfGg1auubPP3lrJg1dBpPrUf0lKER6ZnW4+ARK4/tmjyqeFh+4P3kwm11/JReDsXNX2yX+Z
rRbxeDrrSlH1ZNHbLzbhcC4MNrKBQyClrIDjHuSGjPKONLMhwJEmrD812vh/uCpKn6vVYRKkJoNg
QWe4IVaggC+GtrIeylvNtqWRz5iDpHcpUMyhTkNj9CNUYSe7qv3uAnFocEiIFbZrMPERLxqNv8zz
pJhsDHs0NFGnjYj1+poi1XJJT8zm1vnXtvuHpFkij0Rp8vZad7QsrPpj3tgjYF1YtwWitNckbk+D
vHt/gv6geJxkX5QccPZAPbMDFlzxMFDMfE2Rir9wXvM7y0G/cL1Q87CuM6iKP5og2dBXIR6DS67b
yd/B5nQaOZMyTZf5skNgIMfMSpA3cGAjtZppcKHh7d9k9ANzZBQ4crJjqGFfpBrlI58EqOxNIxan
XfspYXItF1P2yYvSOcr8idWR649CFylGudl++tvUUfyKXpRO8Wx0WfKiSxvyDXjoolT1la++NEBW
bCp/cTOLc+YmoRwHw2dI0ec4UX5JVksTzQrqbaXoINi0fpxm/GDUb9xuVxHmE5ixZgw6smvY8up0
UuC/r9Fan1/YcU0XwpsqLvhCe3IiNL+3v4L6DCgbcgaGh46vXuEvg6nnrHVgRlNj6ei6/4sRAvLo
KayUuUkeC+fcuv9bBa+dA8nKcZg2qCsA2lVbMPXnrkRaM7rbOQfWPcY9EiVpYnxAY+bPpxeMWhfb
82qJfDGI6ljkEgz/+SjbR2SC57DmWzNhlW7TVQdFPAZbCfuqV6Ep27ju6wwofoBrp4IDiIFWwUX2
Ut4U+pp92OopdUSMrcT1GgFYg8N8DxnEpvOlFTFb+/fIVWFQ418e6fgOH/hFEKO89TU22XSlBKLy
pdzNqF9znLD6Y6yrRSFWPu/TpfIFp6VdvuKYcbG1FhaX0NlLj8sGHbmrIpcCq/okGCxpDcHSlg9I
j0VSvGE66OFRRInVegRFm8j5aVlzfcDIQW7mD5N8A0tASXLAsP0qQfnHoYFoPYsv84PZVZYLtu/Z
ghy7W0aVrcv4lZxcVoCR0Jlu4+TRxVOKjWz1wsVTwX4uHKCSayFvvXgtuz58ckwxnIDLD+4wfm+W
+ftjzbRLkvN3u+RCyxJdbHJL9VIkgHjH5NliM2rwANeGDtcRIW3mLFAyauOPkFNLeA14W5HiDGKQ
cmZr8Kdh1aRKCVhnb34VxDPIiUpMsUYFC5Iz5nktZh/IKa5RND7L0cvnTGb6ddmHr25JwApKyELg
nzF4GRVNAIcmYZhbK+FQCUXzZqBmnHpwOHvA6/CdENtlHrDgpYf24y9KAowOba3Qqad+hTrfA3iw
IYOvKaE66TRBHP+g3pXyFyF9dFp0HyMTwu4c0mM4FUGKMnVDU602eGxL0Y35l6tTug/M3xBi2daS
sQMPtp+qc8kq8We9Xw3IzCVPCs3uO1ZqJDlJ7z93+PXHx+q1o418FSw6XRKn2/L8FRYHUuZ1GLRI
RMvgl99LpSXZSeWyQTAWr/a6+xcjO2K/bwxDBLPo6MEjMCxigM/udQRj6VoIMNZLz+7X19BEY+e1
2do7YGhed2Eq2n+nkfz20jKiLPUKRdOtaD365zSGuv5E5dSV8s8byI0GGIjCJ65Yu9N6j5sQM8q5
bvyljLNdvzKJcfl1lJ9lq7iim/MXHcE5M9SWmP66X8DU7z8FOzTt5JJYNzgwdC78K2yAl5KWBf9l
mTdsDEh32WyEIqQeIRXkyFd9BmwOuNdQ7/Wc6TzvQpXx9vs9Bx27hoNZu+JosEVvt+EsYReN2KFK
U6AlGQPtHCCkc7h+Hw5+I9T3qykXSkA3FAYSh+ehntw8Zwn6y3VLOH9VG3aF71O8ytX5KtFDHygG
/ZQ126aOXPvgp0DbwXVTpsjIJoQIiiewKC3ZBh7E7bpoqIp+qZ29jQnxnip8UirlKcwhk4Zgw3qq
nk7UNEFwrdJhW4j3dO/9o2ZVfRwSFjtDAhYSxsTYf9+shnDLEK1MRi/z5XI3hypybgGr0dM9xroj
5F3LJHC2jO8rqfHcT4ChzvYkUxNvjysHTMmuy47+MAiYZPYqgyQh+S9UUiY9ipM3HfuHQpNeT6f+
PTeqh2lmVYqcEt7rf9gh68pL2/sziB9PDg5p1AVJ98qRB3zRaxAQEBKD8tJDmHkqb2S9gTSuns5d
jotIgSXn6Zn1rpV9qUWkNzxM3FJhlUgALQ6Q9obR/T3d2FxhEra6J+wafeUP0i6tnrenI5s2i0JL
KJV5GNSFasBKbmp1SKXsuMLHV5RniGjm8csVXhchup/OIleW980xN7Jbxg7OETzsN2ZgsEFjYsVa
tY+xKk9t4KIHL0TsNaxKMbpPFIS4bYK/Qc0pOkTd7V3C4bz2ic3zOBdx8mrdbz/t8QRJFFlx6mlm
7Rr1gybUgQEjmORpC554v7mbFWqG330xwkHaaYUCzTax362wq0Sr9v0DW2uKHT+PV5dcxyvTdZdi
UcdXNbWxFJu65glf19aB8ruIXXM7jT2BxfcxDyeHQhdX5MrkziCxWVHew0iiQj4W59GsoPys4tYN
jAUCIwRjYxi8OSa/UtabmzxHQ0LDCZQZNSxcteVHWxBjfhWiBYpJs5UeJ5GMXUF2LYk6n1knd1S6
XAm0SEywQT/Y9VbA2xx6yZOZj0QXLXb10bx46NyUuRhrN2GyXXXIV6coioe3rgZQbA+yd391PyGL
Tzv8Ww+1tToWBtvErTKeEzfRlgqJwoZfalzoP8pM1RkoOyfWnRkYhmgfJErXErIbUSpqy9RvV55x
VRHm9r/AAIdUFlEnljUlCEAiXdbAhh+AUzLrLjCV6VVnLOUw8HhL0iC+AoYEMpDVD0yjDfA3gr3+
wvMsiMqm7IxS4M1F5OsFpSPqNhSKqLgVXRjazkk1OgWkvnkUX5s3kzpAbIHgNLWHBjGLIuQODTWu
BgjdYDTEny6/C2na1f6RV0Ja1057cNctOtgV5AybWCv05wAQ4rUCLcQDox5KMKK7txKjwasN/94e
fuZWn1DGHrKJs72EAdhhoh0PPIzz8DIcNXuaRYGuPJiHE4rkyeP+wc5MM3OzYDnf02Nw3tnY5acL
uOrCjsAWM1gYmEm4kv0dZ4JxloR8DewdNw33PbyGQCJNilmVaZp4eKaZ4FrVpHDvVVOcvFe+8IL7
cNo6rT/4AXbOjrkcPeKgDCe47+UMVqaBYS2PmwD37kwqR6IIkcS/WqexZbw5MHmXa8Flb09GMQLs
5og244gdetqx54+gfjKRZ+gMwUzn3B94WA6KUzmrIG2v0AfgWi10kRwSatNVIfSuAj5AT+sIoPSo
trx5j5I3umb1gAxjy9CCS3VeYwQWd4xte+asXVcMgVl8rzFTp7VWxjztdN+TLTSAUuP3fLCJWqEk
KQ8jqZHMpbezpbPvq9Bpy2iNcUKivqgrTaEZEZO/RwMYkBW2GC0QwS9aPgfVgifd5iWF9O0qgsxH
nIUtQKtTVNf7lHVY3OmmtMg2QkZT2/DYHnNnaFebblmzL03GBQQ0S1bNB/1U9tukTlg2FSHrxrBl
t1K+RqaYAOsZhl1eavqCzMYgqLmWy8nT1HCMZCp7OygeZAOH03Wcbv85J7pvu+Y1QtNC1ji+JvEj
vREorSXQpozn498uONfb6nuoiq1LnrZ6VmNXbkBU6jTldUUfcIoq2K0oxu7HQjlF26az+uj+lUlz
OakkE41nEXiebhgPSV9WtPhySGStswUNSBzvCzAewhr4CkQwY1oSNj1BuB9pNk6vssoQQBTJrOsO
GciICteBpYwql5PP6Oiuqu6lLfjMm0XWy+lznqVUYNWfwjs3dRfVv1ClxkPd05UiO29e3axMPko1
AN3zi0KPKq6plyzMi02XwGKJfulmly63fB4RQCqBThqQx3k+kbdeLl7EeyEMGT1U/NAIfOAnjBEy
htC4UT8R6IHKMX9TLwEkFpSgJ1XdVS1s48wqPRb0AU5MOD5+aN8CWpE0eWhmWsWdcADSZpsKOcWr
LBWu8yKrM9lhBpwkf+LC1nbmoZhIT67R+jFR0bSu4qtFMnZoF3wE4QW/Ev5ANpwkJUvs1bISAwsA
A8BUpHD5HP2W76ewgf8VppeMIsQiZIbJ+4/ilh83vJ1QrPopAb6QKBZ0nl0J94uZYZK0emWMY9AP
px6lqXqD7/7ZIMv4+malgDoYFqFmAFPbuaClo81T7CwLhPGCcFiMjEhMa4CIGL93xAg+WG1LaUrQ
mAZMtyfJuukKFLo5hEOjNv1VmfL6ElHVeLVFCmR2aStQdhAj63yEGlxYvjh1+fY0cUZXby3ni6Rx
TSN2eby0UsY8HzjAI7/83Dy/xEZDtMiQiVyurz8KmpBGSMXYKVDAKfgnHjMn4l6PKE1berc0auKu
gakF2pPD03wZ0DSQCkaJJ33JTBYbPA66hb/PQYdZFIHHsKz6iCXjZ/XhLYqtBwlfSIK4uV8vvWDV
UxpkY9ZSB4ZrI0A8pOPd/XiEuOUk+n/p61orFo4Lwi5SojC3aSje/CSxI3297RoLo1N04jVjGvlN
ILIhrY2Jn3XcQ7l9GIGJUd3/OhO96Xxd1mxuQWtcNV2BQcoEhoQUbLQSqwa4J9IlQWtMT/HEep/N
/XaNxKKnUvVMb0XLuZ8VbRZZO9dVztRfvXnde2DdnLlKRkzdvyxGuBuHETcob72x8gnSWurjELtg
k1y+T31hQXoWAri/mgu67Wdm8K+GHwzVPnrcJi2LMtl+y7u9Z84jdzIEHetCR0buWbZOm4YfrQ7z
C9/HdJi68xFrAwbvohTyjqebSbUjFxzcQdoYDYge857tOt6SKMzYh6n03kKGsDsueFXeKUyfMSD4
mnLjnDZpEzJXk0nVllWUlNtixBZ5hv5ya7R3kAakT5y3N0KuL0fUQCKCzasIBdUU8IPSvYqJEI5h
9AFAz0+nzV07zvzyPY7EAy19BHL1s1cTyHHPWP5HUzFNAa9/U+SmnxStg13IhNk4N1A2CXnPICDS
pYP01U91S1hwBuQhmbaDlODypg9FZLkS57UoYlYnhOfCrLiS+1IxP1nEAK9IFD/3kYiQ1cuwanr1
ItFIzMoY4Hz9y/bAiFpb/srY3LunUf15l/jS7HZfAyMRRQF1ALzNx14d/6e8oT26ow7bhspbJ/6W
asP6k5NkRK6C8xwswyG+ivkb2pf4Nh54MQ63gSMUD+fW81W0H/KCGTgrt+ZD/CdrGTH16JjxsL6a
wvay8+TqevHUmpfZF2ji8Y2159ZS2Y/0oAbcLS35tU02gt7qnxRa7C0iY5imfaW9Cd0iVNTD6qZn
MngLhfVq8ehALRhKgmJn3l1s5hhTB41d2UKnB9kUNzQS7PgQBFvcNganw7y4xSWJQjO7sU/Lc9kp
2TuWBmSISzpBcVOH59l3VSkNVRe9G7WlS9pIDe6PV1aFi0ffmGS7nAK1PZXMPxj5uo/eO1dmGjgB
y4QuQqV17NvnSv/oBm+xadyLyNCZO9A14N/3HS+hpMvjhMdVbnUMaHt6jlqI+tRPm11STT3QiR8H
Jac/k8F+QWlBQDlA+RE+jPiapC3h2ZAkM8F47zBeh05RrTA8K2XNW+BAieJGQKSdEi60bpxFrEmg
C94Boq4tmY6VkPHf12n1DW5NVaSF2QUz496Kj8Ax6qLW8Lo4m4U5gkezsS0K5qj4I0iZ0JwY/eB9
yNMGIdyB7HlGkF22zlfr8LqFVXhfb26BemJVeWPWxZUMvjAW9NPoQN5BXmIUBQ7HpfKNSYDLyO4W
14ruQcSLFyhLxFCKqdiveNhDKYeQO5XFt22QWvoAgdNN/TP68219uJN6PApr4Uel5e0w21WANDyK
+f5Tx/jSj7hvLw4qS0N2fF6OdOU4HAKuiR+Lk3y4ppDQjY7svriG66rgGlbU9NNVpKRShhJmmC8j
96CcIllEuNjuoOhYJ2jigJAUbMRb2+o1y4dM4md6JrfVG2ozSzufigRMSnujBEzd4x1wFJbby/KL
sigKb0DFOXwdbPEsngefFDPLBZW0aYB7/vjhD/64/A9SOzZIHil03UVkkZtZgpb6B6i3rkP0h3t2
xf9GhbpM6hrxNIJ2mdtqIB61H22Ba8ArOkiMN7SvVcYyxrKYRKVy3MkZR5JGpI1Hih01CIxYahrA
6wpo3jsmSXzA7AuS99Knnh/bawsQxsE8eRoDCeXR3kwfi4Ik/EPCcXSTWaQYkyfFClQFcDs6oL5S
9rctDSo7ZZGN7v15UUBqNCN1hL6HhDUDyRgzL2RGSDkHlmEu1UaV4LLCo9XLWnfma1Pvpx7BmCYB
qalV/8MrgMRNPsfoEhwUQ+pcHWEI2sIBpCWaQDEq46CUaN0Y1M5j2d2BBM2+l6/xc3u1PfjBhvjP
Jl3EshcDJS/Np60uq+OuSjsnyI0Yki1cTX8AJFsOZqTnwvyDupkmQ07Kkj3UNtowRbq2YI3kXhOo
tTOOYiDIZLuylfViUHYSRx2fIawCpV7HlnuQaIcRdsoaPi+kpZ5gOiA8wmE8xWBjWQTc8PIWibm0
r2ELiVgI8NQymJIp+0oPol1G//TXNd6DDecIs0Ihy8bkDHA0doDwi8im0pJU5fqcS8sx5xhx7RJH
T4I2UVVXNftMdkrt6tgiH+wwTHbyfhyxoTgn6hpPx31AX+m3545GnxjMPMLi6zQWmHhF98KB0lmf
q+E3Bwt6rY59eKbofZH7J02UXZltIz//Y7ejd1omo2MSKvXpuWkhX9qvJ82V2S4FfxASCdbf1IWZ
2JwMbpCq1iqWjaxQBaUOJYZFZAxuE2oKMxmxFRvi7Yp0fwtDFOHiaSONhJJAxtVNZh0ZrU5omi6e
TvuwLJBGYNFNSCF1uT+xKIZeYWxyDkNosktHCFK5jzzF126/PrV3xH5hQ0V1UU4esY2MM1f+/JaF
mVo3JRccLtp1ppwCLB2qZMB5912tR6Va15xKZ54h8ZfgJ4ip8GkU6Xosn//w4eN2XetYbx/ufB1O
5GTi+qS8+OYemwgS1jqaQN/oKuoPjNSyPnK4RVfTEG9DhZdlCVoqT0OXGPlqfExtqio0dqZATbtV
BdtI9+lh3fj17Br449VAvRlRljbqD0eGyEleiwboGIqJ2m2iHZtdW+BKQ58n1UX9A/dpqXfvaGbT
aSSKfwWoQQZ9geTXrC5WUSy/a9OfF9sCn+lgBryKJZok/vCM+xmD5YjZA+iEEuZDlJzpUPg9ugGO
WFUIEpkxC6tD9u6mPP4xBU3m578ceOxwoia4dQ8zCqTeqKRMmEUOZJchrEOiCDexWMIHwlTrQ6H2
5cCaIAxhJOVfiKOEMXWBD6/DPuMOlUhmuVXNIIYmzhN6q6CjxOu3Iwi6MglN0lHstj/Ew7nX3wMn
rJ7FGKRTjjLbwUJn9tFsgaT2nL5FXSAX1+WDIJUOX1XNIesKN9o0IMYfYFyJSe7F7xgHpfXwnLOK
EUSmGR1hfnpB6naeewvsg7V3lz6x/y8ulZLL1TZHV3eTb168edTdohi6UlmXBOj8IWqFNgaKJKMA
ly56nlvmJVMUlNR/RLll1S5khNTvL/b1phHaUaW1QUa6xobGO417jcEVYipoAv5ymM00tdBqLoMD
p0UeWVi0jAQPs5slxyFnZDUr/GCxJ66Pg6+9vtVMASL3doPNf2HAp3QnAljz8R61MWM7BEDfJlIe
CGicgUvQaqrtTwchNrqvH1jZvlGR752kAHQ9LxyuVbxxCuRX3wdBTVgeNXFw7KcNAcXLaX0h+Fv5
QVOvmrF5bPAqzcvZII8/k+QE73tcTxAneh25q/mMXOKJoI9bqQhcpvaEQF1Y1jL2kZw/lIgIxqyk
KdDV7eKm+KvrnAu1F+FS6QYLsAmj3rzzHvVbN1rPwMsTORUeNfGqYCAAaGscR8ZZJPFNp6KBtmVv
Zy6aPRIRd8G3U3CruqiQ5h4PTux50J0mVKSKKeLbq81zPQh+EVdB/hiEl2fJ/zsEiDgs12SpgwRN
briN0p667V/qs222M7o3TJ9pJIV0hDd+fuu/20FLFOrA1DRcMGtmgpd0yqo8xnZJd7BR2XaYJlIh
hhDyvurH6HdlNNTa6R6/CsK6r/paOcC2RTIWZbRD+BNVZHxpgnbGClPXfRh/gcoBHwCHnfK9ars8
Q14199lbAv16xoKmE+reZxn7h72Hodb8RW1iGYY1o++Qg33M2XEoFJpG6DPtfKkP3GHG2gWXEU9J
uEQOTcXq/wYGP5ZD3U1GXQxy8ttdMcHC5PKXyQ1QcpFvflCNpN9wmxnLC95Xun1FExhrUKnJN8gE
D1KCEP+fRr0rmwJRsC+Nej5yED9gY4qtHPMk4JaxcUUO/wMtqlt/Z4oky3iLkEWZ7p1yQtusH/4h
KR4pSJR1HvrJ94+LMBYGYBUWLNvHnz3YA/O/rX60IEDU4sbUl/SPpm3s6iIp+0W+S+G4E2dH+jtP
Bj214Hu7jVLVqzu6ovcsbG4p6Whe2wJscWIL76SXg3iRawHAnYCW6x54iCIvyEaKc6zdbzSl1Y8f
/2KiCwVNVRA+NgBzJlx+UqaSy/y6mRXP8t2pt0RlCV3kjDBoR4FWlqvdNVDUEyk83RlwPGwuQTSs
9uQLuMVdftkRrQ+vlLDXlvBwQ9mhzwV/TTGoqcWXNLn/FAzJjMmhpPWFiJrQHblcN4/8F8o8ZBQH
x1M9VGT4cSJvx8TNqNnwiv+wKc0r9ZkUf1ouVcq0t1lSKX2nj5Z4t/MF7zumYGNrYGVyHuTm1yWi
EaXHL5bV2dnZC+wUmW+KlkJW0PHpFL6C950R68zSBknmy5gWkwwMo7fxPcazJV8nVVSKCBvDn9sN
0q65PFXZbwr52Hhi53/MNuik8lHZs1IUdLywVO6egQSYRkWbfL+5tBtLaRUBN/NYqvNA5q90xOAW
JeecktmGq9raQ4lnk7ZQ8NqzsaKBpvX6WfjvksfqQVgL/z+E/U9N7MzmCeeR+3qiVd8IG1jGIpHu
2Bh0j6PoNcqCcmTbryG9S2V7spaFXvC7QIsTF9jYG9ZgzH+85KYfiroqnpHHApEvYQRRzuIOTGct
2IgJww29XS4fZ2LOALjatJn26PsMJDQkHCbQQezJenXdBqFSSOdRodmMVhn2gWPzzd7lP8kKiEZE
pBonjUbrbF2BT3mlWMyZFOaKGGS4E1wk3vL0ga8vODb+ZkgXjXdI/0puf6xcIsw9KeVLs9A/leqw
488oKmQiPdEuNrH25ll/HN63tjbHG5CDmqI7N3GHUAmUE/ZcEQSlYa/injRUMQIDC4OqYhpde8gP
aoW7/nGoY54935GE/RSGJhvdyEuIO849hg7ryi7mW2Tq+bcp3ugfEgIPgvVMqW+jlppkFqDpSct7
vnahY6Yzt5nGkPUlMqS7pNRuh1jVFzPrqyeyOM4V48SQ0wD3LY/BU5IzNdb3f/X5NfyP+MT7IuqY
s8hcKgD2ZjMVcVVrqXBCTzTju+r+JbzW2W/4V+Fgyx61GR/5wB8ZfUbJFCikBRVZlUisEH+ZY98X
8BwFRPHPNxZfN2Q9qxnADFsAv7jEwR4OPFKcVYHQ8O26TFwKTSJBhe0uCa7WVs6ANdS0vgXkXZHo
AxmT26uj9j+JYVEsKwIn3kuD/GuPQWkVsXaKJ/nY/qhCCMO6trrIGVwF8fN2x7siqBWwIlci1tlJ
iGBJdigXwUPCk1W8BxelkF5kYFLPnfRi3fyeqd6EMDBcU+243m3hCHA2vSHlcrghL5jOowVE7hXO
cijtXMITDIu1EyK25TI2FW3nzSlsIRiF2uBz/gqnLEftqZ2YEPNtKGut4C51E7Rlre7ch89cPuUx
dxH5C42DUbs1gnhvMs+R0xY0iwlRxJn3AnrLSH/bCi6HHsWqh2GJQWRHJp/49Tpne0t5qhjfmd1E
ChANj/JyCkmnfp0q6kyPXGe3872ReNpVWFk+tlaheVLvyIiLddWu2FE6j14UpWgLQC2qYiRdxxXj
0FSAl/EYY1P/AtYuOauUNiIZBZCGACXZGl3XbKuK+Cjbva6YoQLKWDnA0SvGpI/tavnMBJoy4z1l
2hsA7n5ig6KIyeeaAwztU5zf35fVLovfMYK5BwMqqlESHrWsf0GEThqLoFzhQNytAruvPnxRM14P
0JFc4thJ8096seKXkJkQDocbtmzJCBuoO4Mm9eI00Tv/YAS0eidX66JvYrHHLhRmQLNMkPpD7fP0
M0y2jrvE5BKXU8DCN0bFhbE6BiLROglomcFAnujIwjuk4ebufGn0SczYTCMOTf4Tec01C60G8kWQ
E9CAZfOOOZEGNbMwqTkQvCGMbxvZ77oFDKiQVooUckZI4raNoFkVownFNXhTGA2BCTzSFpuMlZ4i
SMPhQJbdllEJ0m6FS86xlPrENE54gT3o8LwHRix4SEk7dUq0NN04BXxW9X2WwJX0YMTmOkkV8M1S
ZNqg0a8zxjprQsLgS2zGXUQFbK+8vfEceH5Gm3TgtevTHNUmswwq3XlUaA62grKOUxR7HqvXOtu4
kZ0iEpOIVjdg1Wt19lJQa0PbwGVsgkK/JMuBinLrBDn/6GcN2/ffYFz77CUVzmSGppW3kl8joT9o
53yL2yQphPMAE3kGJHxHpiNtqI/VUG/fbzfxfzBHOHcOaqNOnTdLIejhriDiSegvn4dFNJTkjg+5
QHE5VvlUerx4cyvzzVjTNT0VjQU7Nyq/EDoCPmFkndv4G528KZs/2/9ANHznK1r2sPzH9VApwBeJ
f3wmVsJKGVcTtpaiz0KSsl7VWkwkkS8imQo8YUfbEmWHsSRmZGnhQbV2LJdVYGciLETRT15d0MqL
j7e1+ri9qTbm2WzBewYnvD6fAfE6nwiK13a7RGMZnD4UwhCRKXVO7otQExPgaNMBt6UCGQF1kss+
BQi9N4D1Wu7sgMzZLQ24GJClqz0+yLZN4h80oY0WiQS1E+n2/PG/k9z2TX6zuzDC6wEPVdvS/tbf
uzl5BYykohMbeNXAF19tnqkrtFTyDy+eYXf/JxxtN/6qAJVyjSm/bMK9I49EhHe9uVwO4am9cfYw
UNDNDNXCRoc0dJwqEzst0+fvOsNXRXNfsMKARS9T7WK8Z4+Ia336ALrjWGKDmB1TqwG/A5nLlkbb
12alpKGsC7DiT8hGlJ7o2i8O9HEetY+klAus/rXFtnex97wR1gm38bQPhUy4zIb/7ZgBi6RsFNII
LBulQGGiBqzqnmb+1ogk1vddCvx2nAfsoh7Pq1EYhZHpTrdFxFX6tlgFnCJXCau0yaYYUMvnBL1Y
oreVZH2LvupOm2M/zyQRlHInN0wXFc7mOUw1ePKqXf6XPsZDp94P6y99wYZim/t2tE0K1wxmHCgF
8829bvO8epFrRlriVAkyMYdDznkSd8aQI0imbrpc6hrav27vPJgWcUclFVHo8xQYW+4QAV0Z8Kf9
Ci+18vS6SVKu4YgWmF7JvLJXRHlo+vEJo/5quSKI5h7pU9FSokHb/+zlRn5PKU2azhWH8swhlek6
DdJLJQwvQ7rAROaE+tVuQhEvwAQB1Gm3b8WJiS0uRJ/tUVuoZ1Nwl7DcOzq5ZY1eEzfgubPie9Nd
nwe6ESADjl7KoFvbt7JzLi6uQbz1xDqrI9x2g2ACGpGzcvAST3Z3us1fLGFO8Yaiyt0EzpBbKTco
fCHFGgEuGkR2SmcURfPLKmBl6Lwd6EPpS4TzLlNrksgDtwk6nwv8iwUCIBMmVjX9eM6c/JqmRR4c
R7BIbyUqIbDHL/mjIJhKp8SLOg9gv9x5fAJaftSrodAFAUyQzH9+eeqYTQhSBJfEHglk4Xvv/POa
K2AtgCDx2v53YCQTzyN/AM/mD4KaeT6zgnG8RK5jTnbwshotmeOeFhdzvlDhXpCFpGy0041GRlKD
Qiz3hEZbGTdT7e+dcm5wdXQ3y8/KjL+0gW2WfH3JgNDzLs8rd2OMxlOHj3FsIiyI2IiWM4GDz1qy
pACbyd1jNC1REO0x87DZbZcMfr3U2trCq3zWvnvjiIEDHLJ1hudeQFhU1XNXp2UtCWmfLaiLY7Fg
/ec4TG4KwX7H/eTnm8TVdrWn8KAikagX6ig0Tp9ukvrJGdD7zUzydQ+k+I1Eiuz6uXHKDJje3y0E
NFZJyJD9HBN6fIkZapd17UkzRpLXpAbJH1bznk6bZ+wxV25B/lbXFIfMjnP9YcUj2N6ghvp53HgB
pYaibJW86/GLS492sgGhn+R9OU1OIgqJlkdjuyN3vm8rITUeDRTx91XZC77fG4NxgZy+WA9VIlYf
iX4X+TOFRCCqWcC2Dcc2eSh3FKtZ4xCW0fdNEGxYt6GaaxSKpo6SUcuZd10iQ/xL0AfRg6kF5bAv
IaEK//V8oC59fC1wZ+jdcKTj6+3jauUlsrTCfGk+VRhvYKOz2KaXeyrMfiNXtnAz1xriYUJ/3NOu
pwvTN5Lq+Qx6v/s6EuWMLBVdSPfCqp58yKxEjJum9S6itT2wBlyFEqtOhKRwQp5bFz6NRjgE541b
5E9MnssUNDy/Gfy/Z8Dzwv17mBX6jFKFcrqWhrOqgPyZPn4YESo33kDY3XBx0AlctZAU9wwd8V9R
YB+k65qw3fnyIT7zA7d4VEEeJDEgqvZ3pi7zKKDYJY2paJ+OvYfbqJKwCeMpOtc2bIPnimFfZ4Pb
sMHwIyj7Ie2DQ3cVy5DM076lkChgzSZmoBALvwTVU5qgJ7ltJhIA0t/OcA2gEbxRvTNdpRPpbzgV
akJ7MsVDFzUbiiRoQQMDKEd9lRT0BL6Y1aEcXseXcqY/RJT0MoHakHWjFzEtVKOJo34gBWCAuF+r
wg/clI2dLyr3KeDrpct2YyZ6924I2EafIu2x8H/MBIrB9aZsuw0Rl0X2UkQFCL4PG64uIvRAEhUF
k0ttnJsYtCkCYx1QSI56WXvf3/W2ap3T9FSh8iECxnaxpdT3ejL7hX7Wzew/6KYHy5m7gZPlpu9Q
jWenAkR6cRAd3KkZdp1gp5sqFnOEveyMFAMttGpHlRGn19lIQ0+E7J9Inv95eqB6zQnCNesLWc32
GGGdmPt3VMhX0wAOaIZP2tEzelxEOsaqK1CXPQCDfOw2bufir/t6reX3qwKUiDnaxrGfbWPLDD66
1Y5j+RlX2HZ2WwciJ7sOfeNcw9C8WsqKzw5fny2AHacYfDucP1y2T/sxJu6fdFMDOHu5BigUJUkx
lMIU2pYRSz5HQskgWitk0/taT/ACiNfRhP15RpfKtomGa//4L6FlSubponzJG6SxujuJuYgHPPz9
9lRfgeDWk5nwK6HS4zmJaxRfz/cmzWtFh+p803QMgMMeg1QllDyg80NiYfdzhRzmOtuuRHEZSTO/
tuq/ccqT/5lSph2OTo+MbYaXvTMWkAuETIITjFTva8uvzLCEYoxHLktoR8z12BsWqKdWzllVmZzw
SLeVWpSXQNzoJUvYsmLtMWaFvyMc7xjz/GirkxaPDssddlHazKTP4YHJn4LFesi89MKDadGpD7xv
bsFFS1nzJpO1uxQuRtgIe83qYOGlZ3C8klJInZ+VTPGBd8FTLfJFwkMoCplCeSEwM6MdJ/s/oRHG
Srmeugf2wGfi10a4uk1hN/8clB036Tc2S6cMtoZvtE2kIKF7rqafaiQZceXfq6QrY4r3huNsB8PT
wxcv/ST954yVPU23YuxLA35FlJREjwrvCeKHy5vqE3SpnOfPCizxIdV9b3FSHoBRJmyJU/OvAtEt
JdR7G3jDUmlGhXMekIYT9eBbQ6UGO+7x8qNgNTOo5YuHYF/WqYvnoCZu5/lPo2TEZzzLY5bqbuG2
SDZpUz4T/Q3OFkKoHG1E8jEyhSCR9fNRsojTYe1ElIN5A6bvoT8sqezYzkQ5+GQh65Pya+jho+h8
LfkfIoYI0gp1l5c3xr6cd1jxTmBMw6n0owHeEXol+K90/KFISkdAeKKBURmHIaFzSo64FgXfH2bF
5SV9Ksmr8hDi7DR/xCL2PVU0jT6d4HKUu9Pu7k8YokPG7t4UHGNdo0QhRg4F32EBWtTmCzEGemmN
JBme9M7mEYNNEL0ToyqavXRxt/46rsoM1YioLTY2jCBin6p8NDO6hKfM4ITjSNv6AZUVoO+Wo31O
mTTE9bSGavCdugDonXqnCOBX7EMl5jQ1g4oN/Q9bOzznybecALUgUdP0flYA9BKVjHUSta242CPU
MG5PjIkxdA/I/AKIHIeKul3hdN+kK8YVPFTZ9hjrXWLrzneJdx41peAavN9XMfKYWlnuu/Apf9+q
yvYDPtE5cu+ejn8Ntd9kLxK0XGvikmsm4NP68YQQFysWXG04fPE2tbXQnFDgeV2c2fMD7sg5Ex0W
I4DA+/A01ZRF2h+uWdpiqYdDvdaSpOWhuBYFKCa/K782QhjAEICWWe3xkuzJLEP/fOHFpMCXYJd2
b7Nrtb+KkC15SW3mUvaGTFIEmVLOsJJuuGPih0lhLd27Pyi9AAx+kmZSlwTXuDSrlLgpWpci9sKz
XUi7WYHW7HzH7BNtc3mSaVjua6M9hYuMGG7ZuTSNtEcdDAIzdg+75GtbVN3cGc6FOva4yZmXoqH4
blaQZx3b0u2fmSE4MM5Hk5O+hICDYiYg0Bc/FsX/2JkTxAY9LmUK2G1/VC6bO0nasFOG4m7i7nOf
CNGwxZWAH0TCDTF8e+Hv2C8pVdEhoTImZ0YrJZps1dMJjxn0FMpILxdP8gS0j6KnIdqE74/L7iBB
KBR+6B/6RMY0uUD37uykrWuGSIwoZbkRnY5SIt9BctMhOTYJ3muEmrzPY9IOf/nHFSwXNSBQKdpL
upIwNq1FYyeJZkY8oe4/U7gMSVcmGKqGgdvHlXKU9hdt0AFkFquw1H8iru6IuangbLV4YlslbtPb
VPum4MFfGKOT2qwTe0LnHUkFQxnR3CdbBC6NVwdZg1jyWsreB9l1Hqyd2Jd46dC3ng3hNJ9ViSoq
fVEaafjIHwmKH+juI18ICiCXhKkmnV83oRkEijxFiXcy2rx5aoN5bRq1AQ8cUzC5J0AmS+GjugL6
8Ptito0BPUvbU3/rIzDdaNComo8SslSXJuH+8p0GUwkMVvKv0wqg+FWiCS1KHlvSAkDfg3sJOZpJ
xK/1NZqVzf5izN0b6BSUM5bVMUIkICpPUCTgeY5qz8oM9ozRXo+V57QQJSAouOVAVhTc2Z7HFREH
8MW8OLW9XVb12nvY+3kipDN3VgbSXhL4DYgBU6nE11sKVQH8xaMp8yCMR/SnLVjyJVbaq+SMkzpO
19mAcviwWtYjDYFaQHZXA0WWJ1ULy9d1DKmPQEQVZQXLF2grrM/nId3RtmovVcdAPG9NuUKFGcfH
AbvnIpGKpXx2IEIMaDqFhYQFeBoOyUa2HsYP4mgHl8xylH7nSbaLzuihB3BLNrTuH0ZD3/uD32P+
GCt/T3He/t/FRRHrC4bqDtXJjpQEuQOJNHF19186I41/Hm7SsCJbqG9NNY1borx4hRYGP3IUVYvE
sM9O5b3S2740iOkXki7rBUBNj9Nvg03EGyW0i7sh4sRnid4WtCJfO9ZdPKbDru+C5kwDBjx+domA
DLewcaDX9XnVPuN2aW65mawWDel6AIAf/54pnaSCInk2Ca+7SLyRs5l7ybT99C/W+CBhyDZ1cmvb
nYsBXT+5cHReL0kOnLdsi7zGlYIZWDjtkmiUeMryeys0YJJPC/eVUwa7rSgNdEOQ7zBocT8dVYjX
Vv0VpNAG6xLY8VaqK9Rizfv5122KfASjgFVOLRXA/ddAOUVeg0QzVxTVnHp6eKsfsBvFe7+wnfvz
VMGJ1Pdgo1cTyvupC8mBl5dpnlFduoDONr4i/pWDc2swQL/p31akcLq59u75BhH5RLyWrFjUWMKc
LoTdUhrxdK1ND14m+zI3XdaTm6yY4I67pYsmHeBzP8dRP/FUK4TiyT/oBk4kjrmq41MfjDtdA/i8
X3KBaintPHYujhgRAi2+ydKV/FjNprulDCp5vIOeEnQ4aB9I44YqR7u++PsGjH2N2m+MW55Pb14s
WpV1tM9dvosDwJszph4fy6qqRAqAkEFawAhoUzButxfmcfSrO2yV0NK/lXsgLk+BOdw4Vpf4BS2C
hmB3OiKUyP7qLWMJcw1I41wh4JzCJ9qd6DInfnySzqR2v22mJE+hKkIugsLnNxf56WigKzPwo0+K
FYsy+riIsOIEco6a/T5OlhfGRcYwTtqyqXQjQ3qrZQb2OQwpgPorUtGUTj1Sppb08m3SW4zF6jSH
p3sTRJ5OOa3iwp1RQd2eSodYaT51rTY8WPog7jdklZ0ahLqjem6QKIQM40fG0yLgu7c1RpbHWPzY
/wNNWGCN4T7u1GNZ1rzu6hiFimvcIiAffeAtXr4ZaIhwavWP+vXKyiGL8NV1kmUjhAEgZvTuUgx0
jDAh2vFRsbqoIx5o53fnezTv2ZbSOs1U8nC3LXHaCr8Ff8K4Ww7TOyFz3/613l/k0c0MlxiM4p/k
EsTn79uXv7mRPbW4cyDVusYOt4iT2Sv0eMB3W74qk7/nGLhYtpHRw87qKyL887Tl0XjlKUIbr5xY
0qQLcjK/AiYfxl0OCUShi9c93AEZUx9fxkKEaoD6PNtJXWVTOwvAB/bADeI9nh+2mqtyNXgLQlfd
4F7GFl1ANo/l8wRpsiGLiUYtZSBwQJDtsdSOUZOlFOjGNcbIv9UyU5z7+qUKSzc8JWHNsCXzG0DP
o8JjhyKoZ4O8GqEHeIIW/UKMOMw+puutXVhzya3BarpO5nVWfEZUtFtYLba4D35V3I8y1xLQTEe0
/OqxYIreCRQMrQd1KCgvit6CZUTRpAPPohPh6OIiOwNUyHqy72imyixiJsTKE7UApQj4y2l/2zWs
QpvuBn4niXgsR3ZPuVHUxHvFN4HQ0DqvV+WJ6ny1C4rChbBCAG2DmTzgSn0Rh9KP+rpFHK/232Df
rK836NYWV75BS7Lj+ejJAmYyYY7kkPzAklT8hKf5O/9iGRiPjwXp3EoVYq9UZAgYkt6wL2Nr+CsH
1tpgcjX0gHYum+whpGK3IHYEsvftfh2ui1L7cQm5tPUrxrnEJMdBAv/3OQG67Bm34NeMiuFBdpAw
2uw2jO/+4JVOOc5WxEnd2FLN7x+Oj9DhqOKzs63EsA9lfgDkOHfInBguC59p7xi9OzU8vbiIxuYR
l2EOGJbUN+rOsw+RSl9C+hpBIwXXXCz2FwJhvNMhB0ioNS59RIh1eIHz6PqKZNUzDrJZV1BMQiiQ
SjlA2+AcDw9RdHPUDhkErG8OGzftcueVWsVYQyf7/ze7+HKtIMOXRXxUzMj3UkNIEkDNHDtjKF7q
2TTSuMRuBSTSz7uCH3OiL2pmKi5PBn1ujf4B5mkRprLYFVpYlPHPb3KELVjvpStXsJOno9zUyykr
lc3hqZ1u+C4it5eJ+u4Qs5mKwmlw1qlo/RWb0m9rvZx3gVWGAoqmMgY4exgyxZ0HtGFo2zqS0zBM
haZ9ACVSYskDzDBb41dI2OgqZljqyosjgHUSrDqWhywILuhUHUdC1OYNkOLtwJ4pRU8PGKcRccdZ
rEqu0c5nn8eKrZgiwKGXMyExZYBfi7w+PzoVOJaiG1cHnrZoX3nJYiVkkdUsEmgNT0Kc5KdlQ3sJ
rEXA1Ny9juTbY+k3jSQzpTYJDax2mVGU6qFNh4thuiFAI0Qq0UMkfVDlyj7wIjw0gRIf9r3VPvNN
wgBRujUAcs61ja/B8ChcUDJf5jq9Idu7CEEUirHHu5nmDJ4TXK4bUazzXuCVWxCi8HWvcyVXurtv
5H2MiCN3GbrD9WWFDnxcZqe204UDWcWp/t5F+QZTy1w7JPDU6buyBqbfsR7OGGP8g3uCyc/rxKW8
j55EwhLOa7Tkhplq9brK0EuDUd3VO33QBI9OJ8Cr/uVwwvU6NZgnW1UUz1GQ2zrkCSS64CQHoA/3
N5bkFarnVRycsEPsp2VEKV/QH1dqpCSdGHHnkM9H/Dt3JFk8nwLiwjpB0qYU9NU5UT3Vbc9gbDlc
Xr6ifQZlu92xaVfHiUwSM98PqYoCiYjFoyvBETN7rq6HW3bYuWAg6VR3HjN9um/GL5bN3A87MoS3
UJkUTQAfDgY56ykXTLM0Z79s00K6Z4OqjiRz6oa2tLFEU37e580RaL/JUG35sWsH6aUVJSt49uLW
PTEfzPMb7WvesAREDWJordpmDOGiWE+FABObhd4V6vt4skcyky8AkiY7ss3KWiSZnzuC8CaCFTY+
XEoBunEWShWLeG8SnFOR3V+72la9O/prOLJy96kw0qREzParfCA8oQwmw9+MU3WcfqoDwLvBXQcQ
GiRqOCvHRhI2UflsjZxHH0Buh6iOF/qXRsDCHXUAsR090jbSqDCDsZboVp/mgDuKDk5sYMpx1LuE
9l5bc6sdX9UvLwOCtqP7DURvRpeLVzlVQA/uqj4n802R2Qy3ybqppBzkXmDfLEMnBgRPYcEixNiQ
/dX0aarSf3LOdNU5WfRDfJHO+2h29MiZ6gWxcrWYZKGzImi7fdQ2+SWtMLcuI/cYDgZrVZi7X8ZF
3Lk1UpqimpXeY/la3YvgMrGykw1BerrJndlD6iDFiqbZ+1AXKMY+rh1SaloypVBDN1Avt0GTEHBd
LsrzYxCnOHc5kHcdLONM3GjQ4Nmj8xudDGOuNUas17SZLSNnGwLu+jktrmhbCnfgATGvXWI8JIFx
3H7F/PjVLwbYTL+cJi0LcSY9KrOgGV+dTTgxn3Io5kaKo9pDOGqsztcMjL2YaGIQPB+pXkOtGb4I
AbuXWin75VLrQV2WGFjPUmPOU83/rhLWPSOhHlzcGyS7Jo8WWuinGdTA5i78PwRrSZuMYcNbPMBa
Bnpw8kd8uaTJW4+vubTBEusnuQRwjivp/QsU9MqhtK44c7TR84+ZOiy9Ucnb9S01dmiE4G5Uis8S
jNS1+0d05RU9P3TNPTmxLumkZp/5n8qOwI6kSST30VsBhcrgbCET4lLVFsCVm+OQfe/HFe6kYv/s
bS2jVjCzGAEGj1zbKJAK84v1okWI/B7FIbJmUA6YifkTXstpziZDF8e41s8nhoFSPTIdBwJQlesu
H6aojZjNUOxkxkuaxvwMlng6djMwh2mN+b56fXF+hlCelgPGrV4cL9gmgjt/hpdCTT3uZx20a67q
UzPGF5CDjnUudS5KdbvvUXS7clgGAeeiYK2ccPd6oADqvrrTmAYe8R/fOJ7RAk/hu2e7jGuJuYVQ
wo8Vru969+0GcuWP8hNHMJLK4nQCcDOD2tiFOMymQdXsv2RGe+mwTz7Cjs5jut44Un4eeoQg3i2Z
RaSjPc6GAs6zNIFLPMcpD+17SIcNMPcF3D0QUSojHsjeUyApep5HWQyQLvUv+ID0w3ztMfexyTH+
bop29vihiUEfnhwtgAoB2g6qTB/dGlUN1rxReBJMAOryVgp99H2MZ/CHzT3G4mpQ2ee7DiI2R2aM
PUICZeFaPO2BN8qtUfDVIQZpJDqfkfO/lVpuM/zgpMEUDcYDTAl6TigIx5ZYltvKvJJjp0/x1tlS
iF82KykavX6MXhqaXwYFuKT2mrHJfg38gWX/ctJt3Z7YfMYRiORawlklLMu3TIEEzUXCgYMCNUFJ
P23+9scLVdiZhgu7EGrEB79I95YfSA0wPwXR5AfFCR9Ct240mLnv/DVBXVOufuyT7EiGQ/OlEGhX
XFfUvUKzEOXr+55r4CIb++crQ0eY4cqR3C6QbE71HSHE2Qd/VnQfnEFbAKrbylgOMUqLnSjda7D9
lhVdcbVfVhdU+ZDXm+EVArgo9A/2eVy2xFOuK6jtkKb4d79Ue//5Ml+63+9zqa+L+wejOzWTW5+q
r3FR293ODNsfWJJwGCeZgzN34TGwe7tJS65Ly+bnAy2D2g5QhQIZyAcH+bsTtRX6tGxpvzwB9Rqj
Vor+I6r2qBktdkIp1DkfuBdCkJLib6KXO0sSHzUXJG0KSKpxJsQjswDOP1OFJ86ywze5P0xbJ3qR
EQ11K1rAFEs3SUnasSbrqRNDillTlfwe6MDfabKltQu+hFj4zKC/2WVei6JxjHRJqs2cs2qNfjWK
gFyUlDG7fwQph5PrdsytEZmBYP3Ymcgpj3qYK0SbFtrQt6/7EoBA0BnT02WWMJuxFQ1Fndgc4Bfv
/4OO1AQjIF1WMJAplMklIgIDC+hH9hjEBpWTakYgTdLD3iaIY6489lETzwpXhlb57X9rZfhxamGv
mQoavYePXLVvdVQk4Ngpih5qsngIOww0V9iLqW0vXlR2JvpDCKmedhXH5OPcA2e1J6dSqXlraox9
UBYwYohAe9+ZoMYlIPaSbXilcHa7CEHR9tsCy57H/DSgAGoXegIK2DaaUpkWbIb3ouFYBnx29FDC
hxV4gTjFuB7KjAv2/ZsMv8UTiOo5s4SBdajQFF8CTIuffozTVuAlqknVleGj5QxGaUpgWe/xc4XP
+lmhKmbLm1WFy1crs7yx/Rwlm53zdIX3M6c7t263r+wBH8/GG2TXMquAlagh27M3KmTlocfMUu2N
o9vaM3QJyRpeb3o2ijRbUj09Gdfe2e8rMLu9XifX+/H08BGBTRp55XqU1fNOIMFcOoU15loW0fAq
A9S2WUD37ysLi0/AzAkLYBGJhpOwNSykna6WJmZgCVgxwlHZ0KYIcQrH7CC6IKptIStYX8roc42z
eXgkP6rVxKqg1SAOIz7ph4KokjYoMhTDr02nrcIG2EgkUfqMNUlewLg8tgjMA33P1Q3g473ruefT
nDnM2YlPhlJFCK0FycgnjkpbPMlvK/aXiqE7jr5p/txDqFASmI5jH0F3O2wxHEb/lPGdoA7ADZYN
UjKuuyCOINAxJTjaxYC02JqEDEUjI0rLNZk29Y484azKvdlpnPFIwdKjhw07MNFOGmV3+4ZWs82r
6aKWPwhwXEeNwco7GsLy3awBQAIbLH1SMHOdhAoI0snS4sCmZ6w5VnmpK9+8FvpHSmFiyCwOIPfW
pR6JP3TNSrFbkiNxZRaXd7Iq8rCVb+WqdOQusHjp7fdNFFVXVTI5Jy+4N2Cqk/NIf7j22oeGijUr
9VzZVo2UG0VHin6hhshfcgCY3K9/Qbb8suylb9zsa/nSC45LNmSVzzxlvGHW664mLlWhKBjTS/Rk
FFBsg7RGYeIf0UFIzCqg4MHMoZFNfj1ZXrY2BK8QNS5W7KBADDcJyel6QiBv7xiQzkZhc5gehyIu
jDS+fv+1/OlJadsj3BoFxXaJyHDyLoJwwI/0MApwggk5VQojtR/1MQFRg3DmaZea1YM1h8JzIj1K
U59k2PLLDBcO7acWV8naqQASKEQ9yA4EA8eOHx9HPVwdMPFYl5YO3cJa85m+XWDFu0UTlBfeCJuD
Wpg35/WYDedETwlA8UZpm79xZJTiLMzmhe7dZrx1rVZSmQ68c5yb6UXtKjU63tnWS6s+Fq5nHfVi
oN7y6Iy3UOaJvHw7NxegujhTzHjuX6VKBMY8UH0dhB6gBr0gRweozVxoVxj9f6bNXGx9w+Jd4Hqr
pqAMJ5oZrPNoVCCMVlKAWZ4BpHCHVmv/Ao1ij64BG7SW6J2/f724UAicy/hyXgTojzbnkXgRtppN
ibQpaZ5X5BH5svvvuBQB9G79mpQEfTLaS2/S9HVm9U6VFrc+paMWHMtbNhFNS6rREMEx8w7a3dDK
TpV/2hSwk350TJ7XhR/fbc/b2JrOr8cXqIlAi7R3l5urmSHV0ieGM6L7FeuVrVnam3Rfe+elwDIB
jKNS+rAD5e8dzaOXuVcc7RqaaftEN2NEFa/HewiUR/1jtqPBXZEa7RedjyW+i0HLOjiLquZ0QIXF
BxWrr1l7LgBRCFAXAiktwKyrPV2hEfcLtD8W1pPsHulEiweQE1T90StVdaaD+eSVg89BHL9gsB71
2/2fQA2x/8cSZtJOw9CuEv4tkabfNF59iDO0XdqD9zzEwFK4AAtwWLYQDTxOgIjJWuZodcPfORXy
G+v7/x1P700tLrZlRjXEdEFh9hBz8FfnEvX31RaXw2CLiVBXK51MHSkSpWiX+rRtiS1mn12a+pm+
aRq0y1/4f9TjZ5K0hpf5r7h3us+X3z6eJXtbi7xSWQCeosajwSNizkoUpApXOwlujiPTTTIaO1yx
YKBKrzmOBFQYQmWhTcfY1AM/rt7S5ckseYDT4Ng72ky4HAQHSHB1kHvKElWocVOWtpCmEAnFT7bW
A8x5e4wj++QvepEKcVuHK6EISGj3L6HDCfqdQDo4sqMFWTTjye+wrp6BsxpsxR+1/zhOrzr+QEB3
GV4EUAYtKdvyMHQdK643raOMJL1SmIXlGth2L4fcJTn+58yY9HjcvxsuHVWrVUwT05rc9M9sIKAv
JtV7lvH2jOPAmwpmdfzbXwOiTvDXS+9sLoCgNEE89I8AhIPsVV16BKUQ7BYHi0cf4y6Fv4CiCK98
d+LVhoVSGiz+JYmW8nZ5mpuzMoe4ribdLcyIrUOD7R4p6lFMFdgdjpEtOakTh0zOrrrlBkq1J/VY
ZNf0OwGpN8Opp+0VbXYmJZTNbidPRYqwJbxTle8mugXe7CNWDEAl/HEMoWxrSHwPVGWyVqGKkJan
9M+1jsp1cnVS1mxn88R+merR1c+5vke+U4jbjPjeL+p55hsaGdq05gkmeGU2ekyNY4qRjVlXl+9E
1EJukmtLjGTIpwALjak024uJy118me5zzjabweazzjmfAG30ZhAucAvG4f9Av1fI0gBg+QkJV0KE
aVR20kHkq+hbVwpL33K+Bvq0BPZCfg7JE1P0fswa62ixnf+TTd1jqIkpCwdsAmu8lLhG1E31eu/Y
lZimrjq9k08zB6LxWc1fQHcOY4kSzwjSCKW/MEniHZvwNDQPGImz8XMEG+XxDybA9lExewkkDg6t
r12kzQQHv5a1/SolIe60EChrXLLkNm7A2OIT3s7OE3I/QaaOUPqnZtYdUZeXin0Sp/SvRQ3yidse
bvCUQpOSTJe0i3I7mKxuN9bRINK2GzC50RsAcnoY1bQtsWtW8rH0u8B32fymwO3/sMDvwZqDAWkz
5B1aU+1jD5EPAuMAVhBN/HZiOvpKRciNgk/UOFizXfBJu2GlSWWxjqxkTgDUWWhJwVqA4CNoP+gV
BrSrlB15FQSUu7XKOG9itjujLh02zlgGbupJ7QIDBhEg+Z9T/xneOoMREo3UsR6IMHBIggpBO1W/
m08K2r8zjJcsQYi4RNAuAWZHpu5ZMKeb2l7zaOPT7ETn5z9SLVUTfGrVvoj9PSeioRZmyp00yp6F
e2R07frFGzrwKFSloei3VLGx/3mls/8YZRHlzuxAtfJJhT5UAZSC50nMWAj4jPocxD1L9hB5biUb
kaJaX8pqgKR+qYryHaqO+sPd5R75w5Ghdl35F7kXqRVgbBjugc2iiwu7d1hyU9juK+QVtho/1XIw
SAX64h0rt/jE4B+YyTPMYz5Y57Of6jhlAwRjHD2VGNo5j3YuJwrHSmiChGWjawtJ1b65IZkSRJ/m
kDci5saDpBit0RAnMkJPiyjz1MIPaWBqfH0dchPqY7ohoY3KdKhk0VK+F+QBH7ih2pYxhWWJskHU
tXyr2WIgE0amLe3cn5AoPyYaItg8V/KcZT0vjeD+8Y4jyZQZLGwNVq33oC+PD25ia3sAgcUNfeU2
kV42sH3WoBqteqdPxRwh+CGWxt34Wq1WBleDGzHTMPDBRtZqLeIgpK8OMfSEGCt3Dg/7W4dxUDOZ
yK1uobqu7sUoJHVApNqb2xTAmxaoPf8icNGt/EgxLhuBgQF1tCKgq6rLICU3CX/hduzXzPQ5FKut
Spgev7Mtdoo6m1pyT515eJIhE0FFXH9iWs7GVJDj+Zl/YAWGI9bG4k9N5282AnjOla4zKf7O6PPG
V0Df2+4qbjXCBdOjJVkDFo8qoSQmQrSIObnBzm+dp/vzBrsNdB1AdsP40vf4NHo4AlNru+xvISDH
SeoweN+3T2GHStd1kuLCmIyXuTT3qaxPi8LywjNNDNusdNmXBak4UZ3P+pcT4x1B+QWktciJ6jwi
PZhBXPikppsveJ4809vIVXgUZMtQ3o21Oegmr/sHqSAEYa//OjvdVdwgFiLOdKeQD0e7YKh6hy4A
r7otkGGbIQRtJIe5ftwTldVzxoXJj6zNdyObIggXaSyNmuoYibIheR6rD6WewqQRbj4OzIxKoSQZ
M5Y2QpPw1w9i6FFWF69q2s350pVqW2Tvjkt/nMOypbXQDTDrH93Yu8a6VAm7Mbld/de95PsTaFOg
WBSVrqji48EQLIsCifmT4mZ46xk8ykjwY8e7nZP2Tbj2Vxzw33BsZIgTiXPn9XF7YjhyYc7MgwCh
QtORg9UwOSeoUxrU8znSMju88feu3+9p2CaNS+rYnEBASYX0c8qd0mRMlZsGZYWd7gHpc4ZIMNoY
0J2QMmqc4C9fs+Hav/7R30i/NE6A7zk3Mj3EuLD7oRPmnAet20YSCtLrMvkXxei4rVApyZWHj32Z
aSkT8bAzH3VzRz7nCN0SbsarkSAUGw9yqRIFlmDdvYO/kGekcDcI3zMBq/AtrRpgPQAbOFbB40Js
qA5jnq2qcmmgOecnZ00QtUI7/2m5gIrjRP8dL2oLvpLexGiyAV26VWInnYftgYYfFhS0uH26efzM
UFk35S6qHtJ+XBVHrUzK1mYgpkAUM4GaA+PJUeccOpQU6iPvpfAfEJ0bIuKWXTGLSvz4/l2Dy/b0
0PC+DOrH5H7DrSZwOOlx+P8yO/tHVkrQGuIp2JDIvDVORjQFXFGuy3RuLHpyZxnw7Ecj6ccYRKvH
zShcsU7ukT9tsg9SuRhicpzlep5Kj0Ne3ebpmBNhyWknuPDVgf4y4Nms6cgPQYlHDNOoWZFVFNfy
l3Yiq/0gWBTsP24tpC/1bEEnZePUv4TSn10HirZUCPVj/KLeM/MVrk6YHoyExROyn4n2juilsLXv
e+ZmPV/dEfgW8EVVX7ZYlScWlJcuhtWhS/R8/eWofhuudxxrgd/WNuQhqpxoTEp5cmyC7QN6ATeb
u/qzq3XacZ0Br5OiOfLhQZnoIP0SchRkNUk3RzjCc27hiCJiYkQGMGb/RcT0EXwbEq3fDkRrChms
yqH7e+Kyla65Hy6g2Z6HTCB4O+m13Bm3wP2pboy3pA4UVgitwfmJE6P7G7NIzSW4xEQIUsPriEAJ
vNuupC6hixeX5Q+gUHW2+awmW80qWPq+Q5yWuIqz2+J/S3Mzbx8ucqXwNyFJrlF+EppXUB/cTF0Q
LDkkn+KAxSRPYyJ/iStUe4aFErISFNCA1RYwueSUYJF0dUgWoQIEawXaEuXdP/chLJhTmitGoAo8
XFK9l0pO9SRC/Ys+hM2oDbtx0BK37whfF+v+U16J2P79toMK9BQ6ni2I+B2r7HgEr748Y5xbwG9t
2r6DABy8yeoZYix1m1x/e/7jYtwLISchYxW1/1sLjUXNKsG8VxQzjNI5SYBaeJSH7H4GX6721c3q
MXav7TD0TeMS0aYuHZ2y2/IyXoDPqaV8lZlONOIDaiczDFhbi5q12eEWyOvn9DoDwtsl7r+aWJb4
jRb/hLMcXSfIGWV7mQvokhio482G6PwgKCE0uF3vcXjANKHaUuSzjFHnbogrALjvQIBJT8KBUJi5
Z4SHbxmOukzZfxfxeweo5QgsjL2LiYP0ozjXR9vFhARoYFNb/63l1q519uVk+szhBSR7bVJEZXnz
ouIhTwikYEPZoqHx82npOVRRgZpzH1XtpNQ1fs35GF6W+C0o6YKVJGuomZnYIukAIR+FNEIoDXZb
f3GVDPmOkFftAFNb/uklvUBrDaB55I1B+qY+bjCZEnSGRLV8KubCOY3P3VPBjrxxkqyPKR3KMLHt
+igWoj7Fn0RcKWVhomABnCa0Qoe4tQA/xWtjwZ7MFr1BRSHKLc/e0gwVsZgKIcaFnE7RCd8Acobe
fdvkejU0/DUPeV4Z3M/annsQ0QBAnaUTHlUobbOPufD5UyBQnQQk0W+W/Aw9RZgJmy2SojIyMimn
8PP/ZNR+U82by5bB7H6IzavPKND6FY2ZRKyUodk4j4hMyW9BaHi6O36KG3b4b//MhElQ+7AW+NZY
1EEZD4bhRYBRZpOorfxTBpi371Vi5MfLs6/P35Uw44EGE1jdA56gjjhuDrj55+C9HNoSm7+2J2MG
g14Ly/VV29xiEFoP5GnJWIjxsRyvAIaYNHu5x5RPBFK9OuCLOxoSs6/Ry9H8gURJm55q0GNVaI/P
CSxbOAO/ke63jA8dHgfkz8uM2dFZ/zLSEwJmzuzAOzDUoeUqIlZY+4K/wIWhhk8NBHrwY7Ns5q0N
nBAGPD/HjlYXyQYdgYHsUonZTKluxHgPWL4MZ3avGk0TojTonywL8PhLhHBF+iCPJRZas8rnzLVe
BXBeYQEKCHN9eg947oZwQbYajTsY10dXpE6js3QvckDUlWsS0NdSgfjtmmqQtI8u5OFxYY+olpAd
6WRp4lNatUlCdw7c5fJf5cYsUsj7j31cYYHYHRIhnq38maTE7MyXHY0RtqKp9XgF7PfvSC7k07nr
3PciNRiPQok5oyAfQG0UNKFlUi5sNZcv6oP54XJB2efVYpUVSlBGCqdPNhp9YxCZnIyql0UK6gnK
jjYNijD2XnZuNFlqoaZ5VB2opMR6ExAJN7Sr78x92OVbVyU3e2My58cXttjNHS5RRMwzkxDwFXPw
cL2Tp4AqPND7CEfiwvf39pzvFiFkbXiT3IDZEcvr5kGpVJX9Q47papRemsu49CRzKScTaukGieNv
2WAYr0tbUhq1Tx88u7aafSZkhyLwQNuGHl3/NhjxXR8mj5tCMjfZo/LJIz1jwjrY0kr6FeQ4Eqkg
ySTIbZeLzFSXn7uTN3cF00Txo/7mCiIRpIMUnvP+ybe/QpbsG78Z15szhVi2PzdJbKbTW9rkUqyv
+OGNxRfDcmco4IXil+nH2Eae1/miOwfoZWoMBG2MEEm4Ix9X69mN14eCDrBbOzYwBv8q15wcvJ/l
LybbOM7N9uSSePIjKeAGUgsYc5ZiM9LZHVVeAuBBsbOOa00Ne94dOpNVx0WN4Fv2B56UnxB8W3ur
nrSkRHAi9oD0Fpj30/1JJIH8TdM66sIetARw+Nln2mMbQXVpdzQVNmbXwWKgkBNDm2Mxgx8LwyeK
CQX9DuMxUhJCL+M/ZrO3SM+gaDsqgciTMA5YYdR8jvuIrX18hZkGF9wfevwktpaXuXrYuTz/9yxi
q5UvHLPYIhEoqbXAiU2Mcdi22JkTf4Vqkb+SJpKOKNzyWR7ydw6xNg5/cLpFFxI24VScYwlOHz1g
vBUk9NnxuO9cUZAzVGgUnP1tbtQ5Z6CSX28WJT6c8x2yy5EjlkWvSZDvXSNI/wo2vSIA1XP11NwW
IHioRC1cZ6iELhAa/OTEyYQzKG77mWMZsdRHziCykPPkttJCdKOjEZizzZAHuovW25F6lx0y2A4i
7njOJtCXGUXX3KRPc79eaPr5aBbSroQ1zxMRHBa3wiwRfXDkUXso3JXrb2umSj04DPZLtUTPWcY1
joLo+ZCNfyJa0QJQVSlK2RurGLzjwmmbHsG60XSNQkNDTeaN1gNr5rqbAwDghrb9rKXLuAIUqlEc
PkU+vqLdFAnIX30/LjYg8Q8kUYYUdQ6m9B8t2OPtJ7zmndjwt5RF3Ij/UdLNzbopE0IwjWJ03lsC
TSCEQC6qVRe+i9VwIGC11JVZsiGhRlMm034S3voHOAneVbMWLkxNlfVcE9UsY1DteRoDD3VRtvWP
9PdNJfaR8IfuEeZSzh7jjecEmOudaF52pPrWGkYG1hHOL38X+jUbkXrMXgWqZcf/77eyAtLmZ5Oy
9lLBr4O8zLNEYeC+86icrIhGrilQFabj2I/6ZlTh8xFPgLedyrYUTPwiV6+SaEWk/UklTe8X/SlU
QZdOxo0gsTC/y/t6ZuckP4FeMIu/iX+P4TdgK9upC6vqUjlnXb19mzo8J0geFpmc7f5NuyknVrR8
LwWn9b2I8D2SPGPpx4pFwoUB8r5HjZSYA6FII5/hHPAlIMfvPkxIdIWClEfOwQkigD7qmpQzxhsF
oqrdVPnzQnoOM04rSKH4tKIa1LAAQj/S2JpgO3XNYEYPRQYpPOT+L4v6Kt77xnJV39CNDYzbEWwV
fJMogIlrGB5LvUgYAr9FUx36T8e/zEXWwDObYeVUxchhHRlwVVDcx3sYACibmSj8AZZT5sSweXML
gempgP29tD4MnLuhxosUGBfg7ivTJhnL+RvF2nH+wAzsKvhIs8jYNJMRFliwX2K0FXYDxM1cOmWA
tSDeOuS/alMaDp1pED1vn5B1JFe77EXi97eP3wPaMtifvbg+31bbh7tSryfcBTpCrCeKgwyaajUt
Hh2sKhQOBEBUWzwQBSv/cTiKGUBBpBy3f8u+uyOav1TURoswvaq2jO/iFdqmlbXeLpvXHY32SE22
CqlgwSvOQS8yhJYvXqjbO9KQHhTkpqx04Wra5jAhnE+8N+zLs6eZOr+/AWw/GYZ4tv2OktEJOq6r
7JKTjjgVTTpiZ5IjaxhyLNyfgUqMxyReBTW0CJ00Ov9OkK25YPnGOF89r6Jp8WDCcB/Wo4WHzSvJ
9NP3zkjls99n+IiLeeAmrCE2rYvkk8g0JvQN2He7DMXhu4eLA6TAqh4SQx9u3u6TxK2vH3VLkJ91
7xHRJnJiLdFpHZpU6M2Bg652OKD+7bm5lwGRck0/9CijBiWnwfKvAyAwFWvyY/g9F2ZTzdKdU5UX
Q3fUxgI2piadgghawQ8WYy+xfiR2F6DgqjQ2wkgGw6/THzg8vYyCO5EhdIZqmhjvIK6nqLwQVmGf
0iu2JIxwT0vRtfDgoo2hl0zWDjDN1YACtqZ7Dt8ZC5u/3xEfsZteIC77gsQzyqdkJoRvy1K4VVka
1Xd9PzCSCZX0rnoOrwO7snLzGE0RsI9BWU3qqPkBXpt5A6Md6M4Wyp3GkSri355t8xSxGRD+BeF9
5/lZjHRK5qsx5Bz6lvfwMGLCpHswudc+UrQ24uft7ZugVB7X2lV/JoDRKPpwSiCH0ROh6l6ii9im
9Y6rGfNilrh2YZpLqOnSK1EcWsfCfRd17vwz3e0F1d1Y+apAdvW7yu922TGUPez9A5t7lEP/Hjg9
Z7uMvLIyBv1Fwd0OFkpTNL/uQ+zNsh1Q5ONdBHMYi2FMabPKaBdqA5wLMa+UobfvIs3WSbytc4nk
KJ6uxxuKF3Lxay9RvL7+QOz1nFOyvAwqU7gJTO8CTKw6+UvymFFfRobWsZpokV7UZRubLMS3+8N6
ZE8BkTvRUlxpHIcZu9sG3A8zR/zGx2vQXlRlLJXQjgGk4VRG3zvn6MdWjUlBldfGg86Pu4vk11Ko
WZb25KqTSt1KoXNg0TqDi/9s1BIA5JU1F9BuDlE5LwIAQw8RTsH5NMwEucXj52O0QpGwxww71y6C
Pz2zg8WWJanhbcJB8aQhNwH0QolnbuBnNvtMEG68G/4h387cqyX0lJWtgo0c0XDBtv31XGKVKK96
1NdNxC/U/TCBkjxG2/7OcJHdNvbYffmD9NXf6mJWdlw5bHlN6KlzaHL9GHxjorpk0nJcwk23f/kT
SmnG3fQRkGXuq3bRlrEkiajNDxxHzJvMA9BBS2+QTyKjpqxvI7ydyb1IxeixBuogeZ8ytUXDRBX8
ow+yER2KnuiqErpUOboJsVjMNPzBePrihxy2xe6fHPM9FaF6AaWWku3pbPgJMFHB/lxCn/ZPz6al
DNzAW01qAkXWbDdGid8MdlfC5agseH3ipZo6s8exIESzDxvnr4l7VROMTk7qjs4zvIZrcfBg6S9N
Xp1DWwgWUsWwk4w9kExeoK+/f2w3at6bhXMrK/jaf/wmsU/OjlCAHcMA1/kicTNf0WUxdBACSIyx
lVUI041qCtGRDdzD5ilfdufMi36FP/stqV25Kd17s850epZNjXhoedbOdUvmNvx1DPMf3Wvl/YEM
yXulAF2BrxYNKpcjF9bLSzFwVBKQTupHmgeqiW59Ui42rKGsjQ/4AXvOLb+a94ePM8SIWDUyW2Dl
DtncdBM2Iz+AmuDD5Gm+4GmZN0JBk8ow5WHbQ0AE98gQrXbtBk9Jac/Fj9vazOKfWXkfF0IrSLaR
Pv4ROmsUErlsC+XHqVbCn5TsASFm1FEb47o8lklaXN6Hs+jzl6VzFijOx3EObszihCZJu2RH96tG
LWEecnuJkqqTyPG8txnskqPp6D7uXbWwQKYn9gtah29UGomPh5dkaRB92eTCg1GvO+Nrcy7+DMx8
ISTI2JoFPhd5b7coA+KYgQusWONOflWcLuTy143jyiwlXvfAeq/nB9h24RO+PUWqqsmys79uccvv
QMiQk1eHMMXdLXPB8Avkyj7y5PmRSadCj1VJkrMS3lUCE/IX2a1INVhVSRDwH8AmC/xGAoZKaBeU
f5o17nFh18tCI8h8SfCLaztlIwG0GLLzwdph7hNMpVXn17hcFwgzCxrON3VK5lF13gF8nH7y5qOG
Amkax6j+kM2KcZwjI7UU2J8Rygyu7iOiIZErWldQV3yNFEnXk+R2DEb+PgaT5/biY/RVx1q0lkZ1
KFgr5og5N3HN/r7UWs/k28W/me47PKxbIiuk9eJkcE0HZTOYfhVSyYUVT1Qv4Vp5tZCPvbTTKLA9
Bo7rmqZse2AUN4I1gkCPWNUDs5BDkG7P4fZqND6lC9eWfea8lYAfeOlZqm/U1vEvVzYsWd3rCdFV
awPoSNSQbyc4rH0pnOBA7HHgsvLLCrQuHnm+94mdNwyjtQEyGZhmnWyq9EoefCJWq6hC5IVygVf6
i+g/W1NJ4A13818k0Yx1W8zspcOKYomOAAuc+/huuJ9mGY3OuBqWMKnAj8QpVSszuw8Xc6d/pjuj
yLccd8lHnv7emOjj1OI3On4O7sD1yQfFMcTHur6vFLeoH64YBDp9nnqcRfouWiO3EY61JQ0GT1WK
EmpCmDo6ItL/cOf6eQaDL5Ca/c3267c5osgwQnZJxTwZBlgfaeloaOf1wH68i8lNq9bWs0W93T0Z
DPbikvycmZx49/IcS2zPplAzFIS+EmLNxRDjEL1ja8juknlivFy9/Dsf75eBsRAGSzbBqC+zz3iN
w4yhI3sWSyaz8ZbIq8sryGXDoChNmEOUHfwaIExjGao5Z8QIFEKwpJdeXJ6t+JLiuubQ8+1d7a10
vIWX5xglzJA3/W1rAFe0/ATTD1p02TJP0dee07/zi+5RSZ4pSYkdmavJNbdcNTw/SdkYXidPwjSm
WQfTXhy3mhXTdj1J4U2vqyiO+XCj8gaZHc3iabXMze7OfRlAEEBMa4qfsCP/dvbf8h8rGy52qBZE
SnKIsTIkwbHPSTPz7fB+Xtj8vRhEcB+UcnDW8bmTRf9wae9rlIiXXJwz4P3uHwsYq/lT1r3/Nl6o
G0SF5iMXh/ybj/SSep6h6fQY9/uoacXVFSxkpd+Rj+qEuDay8QVcnVMmhuGcsmBvABPdndAeRs9y
5XtD6srKbuUAeWvDmKUFt/sl2gdijRPsSidSiHn196eeU7194+5b7OXimkO0Xj7Ewv3BNce+bJ7/
Cm5a4ibcU6HJ9W/HXshQh45HJAliiceQMVFvn/qb+WULiPvZfWklO4Mn0KdeaZKIClK6dQB0cWSC
APz8cF2Y84CA9rAbRkAVWABpmHYopduvcvexDi1HzCzg+E7keg95cioZyEKlR98Qw417psuZbBvL
asYD4jQS4kbkm9PzkaGb0C+jENzpFFrGwpNKMtBjelaF1ZKekOW/N2P0ZuHJ0fPUtoG0byPQR32w
rWfsJ4qR6YSco+W+bi12KKw0dbu8elC/wuwA0c96vjvOg+/7x2ll6SgLX1yillOQBkMdPWHmoMhX
8UowPfXyC9ayXGTE87WdAZd45Y3hoRYUN208rOo4o5W6Vblm00p1JQ9y6vAY1WYqoII0prQ7+0UP
+KCG6DEoH2C/0R5pA7GEz04yLUkft7j8jXGJ4gq2FxfqA1Sa16xrl/BkuFMxGzWJBrTatyqvt8UZ
1t8XV2mD7VQOSca+uZtsdD3+lC8YU/Vi+r0y6aje1NnJx49GO8VH1TQdTsjiOH0CRmXPtWmtBB38
WHXAQLJ0N2Ls/cDrIunX7+3308jpHeGVsnh837egdEYU3YzRjL8MmPVG5RhANA4DOI4lymutjuw0
vKqHjsquJMrVVepHtRxdGHfk+av5v7pboLRc1VdFQ7H5ELta7lTvlIB5Jt7KEA1WR18cP3dzk1un
67bXHXE5KFHFJOtVKOvJng42fnjFcC6pdyQ6nvMwZG0qCsIcIBUZMub3REZe47pPGfHqwbePXXHv
RUtz/izPzrUTqzncdAI3BtkOOEOFKdi0dnisZho5jiW71njYpkogrJtsb2Kb17g/nrLeFVenPPg4
zTzVRCWXcaWUut0uuLPZtXxfQPO8wfnC/TmO51jQfJdp/YZ9hhqIsA6ME/WdjHfTTL2I54jomY0N
Wb1gpW8IdYuI1dUhUPmNVULhJaddMh5xzf3Rj9/umAk1MnKy5FvMWz1SSJNy19U6p72WFTigKhZz
bQ2SON2/9ksQGJStzwTalQ8/2GuneM4MsEwf9UK6kd5L/S8U5JOFTJLitIZ9EbRxbGZs70dUYrZh
qVqH2fCyH7OdXRmidZWwYVxsrUyGTudPf2VJ87pkTDCgTuAl2kIwEvg2jO3MCnNT8Qjm3BDZSi+o
LgLseSl7m7hd7kYvhPesFKk1NwSdeb45OnDBNbfhDRWeutzltLLFSSgqbXj2wjUReOJjtbL0X86I
TPSFEXzm81AwT2uNxbIkl/y93zbjxddZ6UFfH54jf7sK44mhFzBWhzIBnFq9aY62o2gviIVNcoeP
kNCmxen77sVP3cVMlyB1iJKDluB5wVzyHUIJSO5YPatxZ+wa9z3DlyNR+KEhtGJFwaw/zBOGaSoS
bmCWH/hy275CWjE69lAFNIqwEtXXH5DIsTQNP4WHAogUEgFF2Jdzd9xXNKn4vhhMZVShcJ4PWgMV
47uLg68jYK+tkDlw0sxR2b2McsD5BkT5l2tNKhFgO/8EWNkiZR4FRIhbV4+XLw9geR+jPoTtyJ4G
BUftLKduoCoS0w9v51iTmqTQ6nFtV1jt0bwDHh+4yObji5VovEXrQO7S6eCJwr1Zpr+uUbcEAhTF
hjji3U/6bb2hBpUM1qZW+ucqPACY43lwjHOYMpC79+UwNV63QBEo9BgqjOenKiIfHzDcdrAcVVt8
ba4h6p7kfnLAhpfDlU1NcFOMKGsN+a/eN0C2dcQ9/ckg4CgXhdrFh19Q7s1A5RMiLNbQBQ3TUFtY
xI8jZo0BjqP4ZIHrUByaySLka5vO0ccIKX4tO3FMS+ExphnkX/vTY3nVtHWSVA/kbq4JEKLhckB+
iQ9VOyfFWm7X2LTcqO9qnZs0VB191REYzuu9AyT4b4R1F23ZYnAMudplkE26i1dfSEmk5qT9Oy/s
yzsxg9SC3Oo0if5UvoyyL6uVxFsTZr0tf7OdXfiaMFoDRFQoUXk2y3ILBvxyNdTglPiNj+p54vp+
LG8Etbj9d6OW7Z6MdDCe8f2YEs4CHIc60S1OuGvChwkwBGXD6RErXJVqGpU4N7wsfSKJPYZGrnws
hcx1KZ+FRUlCvznX6Zd6Bdut258YPlnAZzc9t9KLAT4h2Pwa/5VSFNZBy39Cdrv1akhPyPToVGH0
It9pfHgjkI4FMILclI23eFfnNA0zKXblVqG0/+WrG3CjXgjlFlyeZru/JjGXjizTIonqHjBoYWW7
8iux3ggPlQjzKkyk8eqd/eW7kluHxOoYdeaJOSFAaBMPxMfZraSTTzPMyTiuQn1TcRSW5fAGQgih
bgVkLtJjZeELy8+g5u17o88rjxmoHT737k9Yn2vOhyF7KuDaPkSVPkPJmLjSA2w+7hXr80cXlC1t
iVQNkb+brUvc2sFn2S4KNDMr58cwHUKPbm5gNBSuJhYaFO9vLT5HqMAXunoPteYrYFw9k6Jpv/yP
zg542kdTTldncO+OBR5rwuXSzOBVUMBBVLXM2EEkisOczl/aUA0H490wevdNZl5q+l9C8Sr1t5UY
QhQ1er1shQuJ6DJ6bTQrXUVTTJp793LNY8xozPP0nsPtYLQxWamptvraskNUCZ/dF/z/3kmPUKS9
zU8TrWxcOCZI8ETIOwG5YzLi9ZNvjbxh9qGq32AOvuhhiOMLMo9xnOumlWric+ROqzdpXfzcyF0V
vPW+XzU1imZ0oP4kb3poZPdcPPZn+14xl1fwQTpp7244KS5X3lSrG10DNb9q7EE3khW++PSHrLPD
wvSbrMkvQdC3Bj753f45DCIsCpXxIIEnefjJeFA0JcdJ2wTC4hXUxPw3iuhkAjRNhUiicBVR+02n
JHoMWx+oOo3wWiZSI2WzpiO3FBSbvSODED4+T5sGHUQOIWrvxVz9vZ/97b55pjjV54wPE6Hy2waF
qf05+YZXnBPL2xmj6QS+zhrTOYLB4p8EMJpQGDZpuZZDv3JleUxSEmsDQgBvIkTaVk0h/0z6I1Hl
vd3ALcMir6ytDm1clBr94Nkdja3K353VtKF1lnH5RHIYdqW1iuB8U9gLEft9auBh5O9qYafP2JQ8
giMtEypNo9CAe11oyofhgZl443jhCrmr0MXzkmt597e60jCLShOhEARwOCLzVAoa2PYptRhkA2Lb
EQc7saE0zL4mJyaRumIPYZOMj+UkBCnr7h8Cd7Nit2yvjZufzu1VduVbZqvv0MMhXwXkU3drByok
mfdVrX57Xatf1PdQ4SVD+pbHK3KbUfE/4Skua5Ees4/cN8dzaz7H9wuYn2Wm+Yj/56E78PTXY/IU
vbWEqyLXvkHcKBJG4WjYvmlcG77Kzso6yB7gHgSDnWi+itZMOCrs6y9PZZmjfPz04Gwc3sHUvuIg
GslmsFbkgtM/j9JJNXQE3QSll25F/BV7lUU8xcngzGlbIAM5qLKakjKqkZNOh9bOBEsvgHurft6k
847ooGKjD/1gCEoDubh54nyBzQuxlB3dM5Y9caYsTd6eoXW58L9ZrEGz0PLOGVqSYz4XNtg/rgjL
kzW59PR7rioAu9aKLYnSV1FuuzWll695OCaqymZxh4IhUfZoql7/rPiymi6277Go/QLmhHSUee1c
oNMwLv3925nSJulrL6xAQ3z6ckLGO4iPBZFpotBvC+K9Q2ehg/xwW3gKG9dmOKLR27yJp0Irtii7
TCB55erCBspPwp3XOXUWsGDPXJWSk0K8b4eJrxUPGyoJf8BVutKTcp6NV9dK1O4F9GDCAW1REaoD
NbtG+zl4J9fpuIkMwHpGUBmqwtL+cTnPOhaBhBWu/xtqDk0Hrt8RTBed2kn1SP/OXALvBtnTizDW
fqrBGh3PWbJ2hwPWj5o3S9QDYu1ckqLDUEtNULIfCyeK1lgccX8Pn7BVseulRfl3HsfdNxWZjxJ6
pBl8h5PNuZ2bfCZr2yCVrZwkeaZlGlt9A+DYZaoiH4Di1+Z6X946VuAjd8spKaWKcQUqnF3HXi3+
qsohCuQZRe2Oak5/u5Q7BGpYHFve+dDrHv+zvb9WF6jfOv7cLYH+5hVVDpwp0pdQOXo6cclZJMuz
6Lte8RFCUnC9IUITohTUZULJjq5wxkW3gsjlq1YQk3dASSVMSlX7gdoEI1eYvvD06npF8CRIT741
Pi3klclRhLnse6zNxqjA9/JqPL3vR/2+YCZ09eUGBqc96uVahewYmqabiQPOExocNGgt4vWKf/RA
mJUDwGqhBZVIFh8RcSkBE+F3r/z+/BDxtmnRdLJvuJgjoySly5ZgZyXQqnRa9zdeUOx9LNudhPvI
tj64Bef5tPUC/Rb+WS3WAsx+5y7Ebr+dtVB3Xp8b7bEBqcX4DFUyGQotMWcoswOI8JjU6EKjWnPm
j/uxaDtHohDQyKFxD5Jzx+3KUwxne56GIBh6r4dMLgdg+UJl1Z1gfBLmVGGKwSJO3y8/ui2lGP3e
eY4u9RAW3sOy5RODpBbQ62ZulyzXS72G+mHOwi51MegpSGE1b84ZIX4QzLdVZAJDZmg+WWvPqWcJ
zEZHyzyInzqalFcxeBmcuFG8dmHa7OxGw0hDlznOG176pZnpElZMPiDredMIV8QhtHmG3CXuMBLM
mZ+JCD+CsvJQOD8LbABqRdwV0DkJWXPM8ab/dkFlYXhT2S9TQpNvQlSEmNFmlGyQtmMZbik1eBB8
15LG/o236agPR6Nh1SREbOrcMLzFITrEcWeb1bFtxMk5GsaHNFWTD7FWXngZdV/Wmc/1RNl8FyGi
xXAZBh2kZQdRxLxW2dzUdHNfDI/WIPzb7mxJGXOya5x1cgb2iwHDdYK+tcUBCX5QBqtpM0P2Olqo
hhKYcueWk5cJhNT0PDso8bAHLrD+Nv04eIHZrH1rmRaePyk6Rw6uZMtEMt08R1EZ1yoquA2K5c1d
5apkSYn6N0pBDeEdqotnADPHnyc7sVSyYnGovMOEwSbtSRyqgr7zHH4zXUNgC0dGqAIME9r/XPVi
hL2IqeADf2WuIq15rlzSGUM3gPKZ+8pjT18HzV0Wn38bA1zzU4FpKg4WsrljHp5XxDVwdLWKKvuh
U9OwrjuiTpoAfB5Fs8YciGiEDC99Y/zg2614htAuz4H2Vxvp3xSm2ssDodN/H2Uh3IX9tvA9a/hY
Py7vmm860ByCi+ObLxerh/5TaVRNKGkNFP6LR8ov7yfvDl2b4WnkSkOFRqNcNL4zxP3h7wBufDSs
IwrXUBDhyAErnuXnbnj9aX/Ys5b6WhjiZGdJpHpSHYZL2GQaEic0gg74wRCH2LCkFo8NtalUZc36
A8DuenNhBT8TqA2w8FOm5BMMgCIwwr1z+oM6dHknvNngLt5gytBRbseqAdU/7Efy3d3WOXHdC5BT
vGersXDGXNW1oBbQK7f+9Yr8ACdtUDqciooQXp1uAXOLr0ERIMidH7LKw4SgEx6T0ja/fcpJG0Eb
+s35tt67grfwD7EnM4TNepCLeeCmcfs1QbFdux/7qH/fwC5eL6Io5LOCs1zewRxUW7rACUfo2fON
m4a1bHxFWZejCOPWHhOatAzBzd2p2t7uD5MTRb0mCkNvwIgfQXi5VEeex12xVMirCHSv5wYWQyPM
xqog9WLAzPzWq+S7zVhyb6Fq0M9w9MshIISYBFaEMiNlMIZLpA4oJHERrifKghJ9iUyclyNa1lxC
EDkitBI3Li8NY8Gu2I7u2fhYrurxiX/1poXDHN+H2/X2dofQsg3BUkzD1o1yS68qJ86RIOGGxJEx
6Vco7ta3Z5Ley0sAHWS2NVjasmObhr7dnT2Ort7dlTTPaSoiN9QQe8Zf8kK1kp/Hp2ZrdfTpfs+6
75/X18dR8sFeEf3WL68TPTLD9BZsNtBht1rjKwqQwb7OLhmJ5K/EA33owk1EksA79Svm76BfBH2v
mtdX/JghhVU492cfPG15+bWykHe6BuJF6GWMXCPx2czxgbV70imVorDT5lQOKTFHrIHHtapPinIt
ta3JpRekjelmYkqcNmKkQ8znlF3ckjyvti9hwgp3okydtaEF2Ee3e12OKUm6Qa6K0t+ScGTObXNZ
fFnr1YvWdlzRt+SwQcmG7/jyUWKHMSn+kC9SuAobL5My+ut4kQOw6cL4gKoH+hMDEQ6AnEHPYoTq
m8TL1lS2Tk9ORd5vRknV+S7cQJ1/njVCT6nM3evdQ4T2q5mr70z9mFBCQYsTF1rXXxJsxXvVHdbR
S558P55nwdT08hkkgPDbp1LpW+TavNZpdGTsOXZAr8GG2grk+r5XIXThWQglnPAR1G+FP06YkvAB
Gb/HgkTuXJE3AyBa6I1oKp9WWzfRoL3Or82jIaukfUYU+RYTjMFSEEfczzuNly/qL9kJImG7XLdj
KiUwgNxKYcrdssuVvoT5EbZUVvj7CK+kjc24y9bzrfPjTnFxv652YjLt3NgFxAhknYNa30gLwZEX
FUwbdrL/WF5kneRduS+Ei9gFDToz3PPtDLFLYv2tbEybO0pWn0O6AjwJUHLiPIQ5aNnrOt2D9uAD
nIL7YHq4hQJeVyaRtWsJ+vI8O4cokXyBZl+iWfSR3ZUN4o8YBGEx5Dt22PI89imbJl8VbWTCuXxx
AxwxgiS9WTuypFzimWp8xtii5RYbyf71SRWOjkWsg+ppTDfJK6Yf75wCnAQKkHQ50IJjuF2fDwiN
3hVL+2JfP0ppREDiPmxdtptJROn9bx3oq/nAx05SeSOjwJHUnMfgnZaIDOb/bYCJXSWG5cS8XSGm
nvZczkni44VquUKixSbnJUuoJgVA9YrG1JMZirWVlDW33cWEFXfpLekC47V6aNFkyjgOl8dlhsVk
+XG3gyi/ssmit0N+8TJxNWgP1hHSwpS5/HLqMWEv6tZ4LE75sJcsIJKyh4zcZh7nwDuPYXwOqcVq
WrVX+RQK6X/MulgMb7xG+FA4obX7n1XpkdPdtk9jm4ZBYVciL5scXUgFZ11OwEoKtyV6nsxK7pyt
1rr26joU7oyhyOdJTJQt6afGpvk5PQa37NieSMZxM73hUYlxyrSUQSaFDt0Wl178nQpdPUuHUeqX
qdj8kZeRcqd/fNpXnwCwMiXsA3mQ6/rpTi7xBIymrYLUckmmWWRpULLPo0pdj8qPAw86roo8c3Jf
S1zfmcNoR3ige7c3mzaC81UNmw11s0FkCbWAyTYD7WLu2YFX5zmsoYi8pjyNQuhP4asVYw28RBSg
NhtJsu9Xq1BAhz8Mv7nHj07baOOeQ58tDYpeyL8WMnbgpUns+IM0VU0a/A7GR8t/H7k00i9J1129
4FIxGbWrzurUa9lXyo7BzOqmOOpLeWBqQo9+Eq5EP2ajlpcSsHrb6SWI2nqIHstHHBXG3Bi+aaez
GX8d7BajngfjFEaveLg7q8dj5psywNxiKmhYs3iI6Oq9E4FAUkYTMhNFKiOA7RoQK/cQfjNgzZ9+
iVEPg1Mt4zwtuc/ORon/3jLxpESXMzg0ZR6xz7QJGFIIEfNZRbiX8ZYc+6fRZHwkQEHDHDCRJdUp
P45HqNIWu+3sQOPpjX5Q/lxvNN+ZSg3amEjrtOJaN0IKyT94glwlAmgnIC/X1qEG0TZFzHJPs9nV
UmEWDfgKnFoP4LyI9uID4SRKoqeyt99rnDeBNuoLMA622glaMvgE92G2Or6nAiuSrSNa85ZrAfP1
gcNhLZQLJMZQyucNYxVsqWht5Jgdy+8eOw83MrUK3PK3wuvtAr6+oSlZNL/gNQiK7aJrebiuC1Du
5kveju0eci7DznriEtDAr0IM1RnRWJWSNcVkCSY2KvU4HDyjfSBjGYdJY6Yt9McuEHBFd6GMQqwt
tQKPVPaloVSS/apYO7FSJRlW6+MHBTRRbK0or9BO1t6diets6ArJMDiiPWiGEbGIKrwhzLh+ZqOv
zzpCFYP5aPGfoLwvXLmcM8gv9cfc+uS29K9OZUoX91MDyDDdNTrCYNgePduS4PApBVHKDfm6Suan
vQHx98r/6Sc1RaQVx46gPxnP0/GTeokcxkD12Qjw/igsXQwwmk1ETkcRZxnCNyJWfq8QxJXCpddx
CSfWuU6pZeHb5S+6vVshemZEcjPBqN6Ka+yekMWaZew2Nmw/o/bLIowG8e9vVTKpeOV2tbH00vSY
mXV2fQEjqk/QcmKrH1gYrOwKQd1/uBZREmEXj7MNZE3qilIp4NxXQTsKl4tWE5p54V1ZxAnxLmMM
6fxxntguOucOoP5xH8bc1WtQC2NaCgtvflijZ0PwQ1xImlq4aLluJQ3nKUO1TcrdfqZSQcbdvPw7
GCJTUOB1TAwgFulGr5E0gX2JDJk92y8bDNVNIxUHPqSY9Ms4uGYob5u3i0sAezGIc6I+KiXMfDVZ
Kb0gg7NIjof2NLIaQZB3CQhd/TzOEe4noaPFpPk/m9DC+roun4shQgpju/+yXnZQlkUiVa+kztV1
s7RV9jgvSr4d2hl+YO9abu0Uqy1kDNR3Q1e7gTCy471fIEamtF8aJFltOsAD1Gc0HtmbczzXlSNS
1t7aGzCUsxq27VE/fVL5jvVfWOYVWKTKz3JHkYR2SxvWoaeitUPd1APJRSLWBq5Mp1eqEhfOXrQE
+EprDiNa5WCnyZ3ah6SfgJ1lM7WnEgDVdP+DOsYjQfwi2NxW09cHXk5BcIijli0J6f5F1kEoPMsN
b15SSFmHRXM0RO6Vd7SLEx7ETubS3h0EtuQVygjeD2EjCaujEIQhdr36PTyF6I/Co9wpO5JlNbqs
ma8ufwwBzFUo7vKNXU3DmHIgbwzy3uc8s16rgybD0rVUDB5Z42jAzj2CmnWfx0hxRhtdrlEkmCke
bGYtY5dUHels/M57bx7L+YtyYjMQdm0NCod3zakzES6yvqtl5RUqSrCK7608gez1bZarb4TrfuSB
qXPgyvbTGW5MvSsg8HF+ZB4MT1vY2Darxn/yBtlGM8kca2GWjyIXNvX4syab40QuFLTzpQ1FTmQt
aZHWrfPsL0iSDiOvJ1TCW+uvddhFXyOBzzA3fYSdQzWWTAuXlCGLR9S7uuW+FES3n0S7P302YqJN
Tx9ubHp/Oou5177pGYmXFgmVkqROq8LKPyhYsSp9XZuOLtuAcohLMOHNKmJxk8oloE3yC/lAarXV
1cSCqNkAwCbwDSREhKLUJSX+nD35AOZ13efelDSu3ITZsNdkh1pRa/yyzHnCCjR4mpt/YVPg9uR9
YHUJ9Hm5ghK0Bs8YvkC2SJFOP+vEugfmjqYjXoJ1Xas+kDoJqBNT048g6mCfRKM5lGBZG46AvquU
jbDakt02Yz2unZkmgLJgoy/gbvXS4/EYe/3HAWN1DdNfNUlGfr0VhYBEZ6WZtxFDCgACki4ISrtw
otKSVqGzz1PcFUrfHiTPnPYwLMfVq+lXVoVxY7INqDm04JemmWZjuRjbCvWGW8Y6z4zQBqHoyF7f
ey03G+7vh4v7b38Mod4QW5L1Htg/+3NayY7J4w/iq1rDuvQYsgs8xZbIeqWKwpg2F6lYUZP4xT1Z
P7jwr0NL0m//2MCqYkrkHil6jiV8Bu6r49k35QNIN8sszNNVClFFFialPcLzbvz9DyYvMcezksLO
pzjc7XPQ9Y4PyVfQhQZkf8KxZv51Un1Q5kGJ2jIMRhfHmas8muyQhi4Vfn+TAj7ZF1hbSJCk0xKO
fP7vj6w9z5FRexnMjkfPcY+UF7TlZvifbtiQHLybfIIZ3GNQUsl586XYqlqsVeL9uJhxLvJKqK75
GMxMMjbTWH9qy8K9FWBNSkcvycmkbzgu5AtK9L+PxJW9iKwaVP6PenU3fZSZ2KkzeHdJTYi4Ee4V
OGp+yYL6Jj0JGs4y9YUmulbXhxN7UZGj3MsK2ygxmEJlX9lK2AsqOC8OdP3H39qTWFDS5nmrtfB5
XhPVY3h+oYA645MC/l8NctFvX0BFhFXD618AbnS/oy9FBcLZPJiuPfibIfRgeUhrUpRrbcdw85AU
lecNtr2GWhF2bjm/s1iKlkZSa4WkWjIgf6ikuR05ogCQjrpg/a8gIioJAz0pkTmpYkU4KomEh96s
dDmb2L9p4Tb7kf+kbWnSfgljmMl1u3yzrkGDcueb8YyJrl/wa4Gb8XZ7TPd6/2rY/FUq+8i641UM
jYyk204HDK17ScSmMfyPdL9avGA0Z/jxANZ4wUM+ot7iM3UHZWMyNqN5AzAokBR9o+DIN87oWJBc
zPt+HJTpqNSwvPqHoPy/fyNR03gOS/NCM3QH+F/n14uHcm2wiTvtRnOC/tPZ5E9Xd+Phm2pf5vLd
zo0b27msLcrcmNoc7fTXBGZYYB4VnGzTOlsaY/WJH0vS6GTeDZdCxYfODS6P6vNQCaX8GRrp87ro
UZCa0WwMoP2Ypg1etYy7PFE44m6hax2pNR1/w3ISf5lnGPuBjld0tvGtJnoVnWo0KaAV4LCgQiWL
E5zAoWDlalrcnO7XgGAkEKxlIVNRJwlpVDYcTmLY98F8YPau8IVWHLf/mspwzUy+v24ulaefU1wY
SYgJ/yNYBSCtTP0zS8mxqmzpNWtJ+6fOYLVy3NERCvsgCQkUR8y6JdycBJkEmzOb2H1CMurlWO5X
6/ZY3JRq07fpUkqlVafQQH6RWG0VyyB+aBvCBqlYkeyNTBRXRMkaKcv04fRM1ZaoHm4+QzO1rcLv
0Wneoo9SiqL8GM86D6/HRdoEBDQ4DPHMLMZB8OdCTDO2ksuKDDtK7Qah4xpla3vt0xohVUp9Ap59
F+C8p2SI1uwhyDa+irwL/5rCM9oo9gwhjiBQ2I1xgnHrOqT8bdZFWCw9tinI9J3jP+VnxrNzlpTc
x8ykc3QbmQZDmejG6DHnsSDQpG2mZnpwnQbxYUWxGqT7e4zbJG8z2X9J6npLL/vGoHQcXOya/3Q9
8nM+H6cFJASjjARVzV9CAqJbyuGo7d6VaZfXlNoaOAzFHRuP7p5yFE8avr1CYdWmGUSNjAJZEVqu
JpOJcGZWA51ZaQCkA1iyWg9U1pc6eNEVBbwplmJXROXjSIvOYRkyWJIDjVvfw0GJumtE5jh0gGCY
mtzY9ZKrZTtC0fU3SCxsMRTsn+FobBexzoiyqbXF3oBEXVgXJwOnFwIMdtEmOgKhsKiVZeyj0Snr
5S3ZSfJGwzUA4hq/1WxosKZII00/m1zww5BgXpFyYhVck+JZ0PmuNSJsiU2wNzYjSx3y/M56SzIB
gMIIAOPFN7CIgz2kPYDIbIXShd7sqqoy7gUUWxo2ul3fU7FSNYMqCsOzqZlb1ReQie40BW87KBfZ
Lvdq32axETuP6H0k9cmE4nc4JA6wCFm4hgz4FTz+5KR1Rg+G+eZ7pez2DXEV1+FBMDVn9Y41JXTq
usP1LQ5Ex4ifEsiO8sjguteiV06EnOERNzcqxNJy8ic9tPvq0IQoAxRaNkcWOxw88jfD/vzAjFhA
vdznwepNQq4DF/1Hf+CJmW3jl+j3iOjDpBXtLWMzmsGs5z34K44VKN6dDEIGVIDcxAmIK/L09smk
cCmt94sQDPinfLRZ2we9lU93W2nUJ9KAm5cRQb0fK3OZzQdnC5dzZ5ppg9wIH3PUwTtA+IaOd1XZ
vim9ulNSjKL/maIhkhM3VzpqoMZzchLLF/L82b9+OaKnepD6uBfbhZUd7NneeYdMfHScv8YTSvay
3Aigrzf3ioUQY31liC2pUJ17WcPYg3ix4OKF7JxBtg6EcyPBH3IgA3dI27J7uJ57k/qWi52I6qR5
pOTjBFsPFz4SSNOh1RGlVKAfKK9f7I7DazX9hDYNeA1bEQd7el3bmv7g746Iv/vNrrtlWhzDPg/P
QeBiOFQMI0tBmqbugoBbu+YdZjXyGtOiJlgQMWJo4NWQZN/85vb9vjGLssXo1P3Mp5MfgaL2GZGl
3vf50v+ElYPQ1ShAaSNUBGYdl5eDWRWZQ6yluKfOLHJ5FO7tLtAY2IE4bDhqKVX1QIKy/FTgnF6h
2bWy7hYrQbEBVJeo68Niawqs5kOfPkb42EL+3nidQTaeBUchkRgFRlyUek6gb4Un/e/mdLtk4+Mk
dyrIBcGQDr2hPPJLwhgW4/qOEG7yJXHc7q8b9Ctl44YA7tZvjanjRalJQ/Y2FJAeO6QWHTpm3B3/
2R8gwVc8yGlLJjSa8+LL8/BN2fqu7J6aIXA3Tb7Ucb39AUBRJjaFmWzdRxdoSCUF5n+v3Cb3Zrv/
fAsIw01s5FFQHW0+fQBCK0oxWagWyOLcwgo0yo+c6k5p9bVKJrzbuC9ZkmERWRBWckRsdyyi7Gz5
v5XIHqYJr1u+7T4HzEnoikTsetO3JxvOqGt4TP23+c4NWU4umfDyNM2rR2udU12/VE+XdW/LRn5k
0D6heuURKAkk9OPt2x3vCqIlCmgGiyt2o/V+X324GC3Jt2Ao9UogFdVRaupTAN0p4k7YZ2llfb7c
4vBauizGZG5xwjgN286nD9W7/91FE1EcvPx9oW5w8xvbkf4AAi59UYCf7xfMmn96ipo6ex5A+re2
7n3Y0ZBZAE1IXDeyAc3TXnKRe+nSXHYaCXJygVivprs6qlKb4iMFzyJWRmNdasVURslAmIdGF6hG
ONmtSqdU4H0Sxe2Ay5l/0gXPjeTsrAlE1kVAtBFWZCzNpW2VY8VAQUJpVQfvEXj9w1CnJ0ZKoOqP
eBBokQqCOnZhjev4CK92JMkBR0BWPeqxrAgNtiP9KD2tWzlqFQhyYJUkPFDZ3FeJ7MHNDK4yoQ6V
MwuUS/DGIFErXnze6xjyAAcOzRBNYhffje65i2AsTh5k2iCmhQpuMma7lnO2zhBPMVpjNcIRoXEy
FsjCbbMl3HVuOCosMF871EOF95kM9B8juMJmI+rvZnwGtLBt68NW5DNgIgwmZc4GhhYX8m5LIOv3
EpAELuD5s5gfHqYYpFQtjnIJPpTjqPwMdOa6LEESEngMwa7CLscNiDdtykctQFsz8ULRgtpGqllk
J0iYyp+2cqvLpvwMz+0gtnm7vF/J4+amoA8jlh9cuRMX7qnUMpDYW2iEDdiTycrqSSr5CpAs0slt
ND5c6RXSuaayEuvemA9neEIgnZvJoKRp2lfXJLK2kwxkyB7PsPtmNkq8OU/RpX4PJidtR85pMDw6
rli79QOisqDgC5E/cw8T94F6I22IbnurGve8OTCa2UvuRpDoriG7ogmI5v/E/5qW6lt0NWqEa7t4
qH1glk4FTl6HiwlAsQDhV3/PGFVjZyyQww5+bnDpuflpmucrlTLLzxWUyaYqvOwgm6PzFdua+gu2
SoMIfYxiDbOQHZ1xNBQ2cC2qAcz2YSRKrDZ3U3HRX9lRWRX05oHMu734nyUMdUBLDBttpRicO0CD
ThCRjuLVIydPujb+ov8TcibyoDDGSzdS13iyRJ1cWuANi/+rBLR0fkTnoonK4uyou6EQdcCImON0
B1F8YlhXO6zHhNrmt7n5B06MJIupWs+cPUROzRm5iGOf6BExAbQl8YuEyD4otbt75Fzyk7idOKCK
IAYa9q0gxMmxySgJ3aziGJ27ZR5WN7qw2APl6BzjUT5MNUcNKuqCzauLfTd9bjAIUuOaA+0gVSX3
HMhhz56ef6pEDi4MeqGHu/6d0DrdZPWg8jC6bJiqr5S39e4hrd5lQcHMXf/u8ryLeb53JAZXnZ+g
jxKn4o/PMXRDoMYKIRO/wjsqqQXxx/00DzlTHj1o8g2y8ro1agyYs/DSF72CDjZ486z1n6a+aiIG
GDp0b299IPveLYxQmIc0EjWvg0hKcu0Jfitq9M12CptinAi7JJ2WUxf/810rsRA0y7M5S6GMsMok
ZzJOfvz3aVC7sZKRTtFDdyavQMTV99HtYZs2wEdk2/lzLrcg6lyrFSPLJyrOHG7w0GK75OKY+Ile
/Jm/mvQJqAFoSnqapCGcYEO3F/hdI/QjccPSD1CHvS4Vp/32OCt3ryhERe9Tsa6/ZqSFiQmF67fw
51gI/c+UeB925ZqDCBHEUlukfRGQS9wziIa6R2QBxu86iPXYsPJQJzqkNrv2CzvmB4qO3R3JWWsu
d1TUwYK/ubKz0k6ihyFHYYHdeGgdrJUE6zt+MNImjc9OCzWENXV1k7I1ZdShCweJOpScw+TYTSU2
URdcmCJQOyHyzECNIRmxMalqYZhsr37cB/PlYSUu2nczgF4xqyyrg5Yjsjx//5gx6L7LMEVzwIgZ
UDNgq5Mqrdid+T9A2vrj/mnF9Pi6UNmDh1RtobM+NqSXlQv9Kj0EdzmgkW6XLjTwS1CQHtDDnUox
RIJ+FVEzHR3Rdz/AioOTaHGdgcRYIH1sjlgsHNXLxl3lylNWSmPltHAMDXtWYjZoAgpYxUGGGwqW
K+rgwu9mBPmi0SIJdSbJD7TEkRwagI/eLrpqKfRpxUyStbsbm91ReV+DzGHdvIPDsARKzf4ZM5cb
Mk0mXBxsajVbymdP9FuiicSZYQp093rQk+FnGFX50ULPWsQifzWhx5gLRoNs1erVINBxyK+mm9Q5
nGrNKjRFR2CMDybiPOPzi4KXuiNREsYfY0EjWZy9T/WNzGs1DPdI1sG516kIaJLAosSKYpxbZ4+2
5zusXQ5v4D8rTAWSu4D4gVDRkoXF6s1MBW9FayRiiyN/2tEBHuenyhs9kuP+DftJ4jj72yzZVC6y
THFWzcW/lRRVIZQcNJyzWs2nz6b7m6UFvWXA4529Bp3rnvhluuSdHgllngjkvirgid5NtCLcZGng
PdU943TWSu1FWzsvTBoQrFC43iSxas92jrEq3bxJZqgTUCn3d3c1EK8Ne8inrGSn+ee3CXb8Rajn
A4dXrcA1UgvcLZoXsEBXa3lE6LjxBnL6eGFZxy4arbIQbmo31nrztJpbm7/YYHfKN0FcNIwngIOG
81c5Zad2VW0mlpbwG8N1+D6OjwkOE8tkFyvfw17C7YdNzGVvNwZMgbzUkQRB69Bvwax0DbJgXibe
oJthIj9JqaKT3yyTjf9Fqqf7Olk98tWznLqf/zxPpWDN+0FG2nhXPhgBupqjFuVuv2UOdGk8sYX7
miQwXE7jCIL1kRPzkUSDfWHxYg8xKghgaE6HS6XWxhUrJQYCPZMnwygJcJDAsx9ElNp7FJlF5vsy
uBnCT+DuOawP7hH57Rn9Kau87mnX/d07V18vjfxYb19f2+C3xQoZojuicJHAYkjaw+t00PM7hGj+
eoZUZa2L8zTWWQtntRWbCmtR/L3HL1VSGn4N7S+nVlql3lvTl8kJdEIHe5QlOxzstBnzXpSyGRta
Gg7pTRU48bbOt5HBjY/uTmCNYnyMtHA6Uewp7DKlQSUfERm1azeDSPCdNqw+Id5PUnLGek124hvl
tNfJPUVgucszivGfpVghbUz8xWu0s83vGrWX5nDp5K5ANOpgILoNdN6aMG2CyzZ+1MxuLuk7HKRI
yq1zIVqECezAwet4hhT0zRCt+CfFmfB+jmkg0QhUEB1igt67H/HRsZYJ/7fdcp2N/IxIg+rx1Ogm
BAcRobErh7vDHMNb77gpE/GPs8m4wZg8t7tsH5Ka+I53aFQZcuSi+V0dA4u3vLSmEdwYS2O3JHlz
c4axX47PKoFGDnBLm/ZUCHKtIsUNF5ksFgIhiZAYPlwgLQfjtvUevOuZ1/C2kqeZwaFEKaq4ApLz
REy+Vy1MiuQDfU01yGPu9/SqeImCwjYj8vbMv/uVGAMHkQZvvNmYJ09Ui3X5GNm/MkS0br9Dr1zJ
cxBtGmVcOZe6FtxTB6Y1Mi6OgandF4MuAC2wpzjvFEHyRF+jdGMFHuULuGGqAYm2rKSkIejoHYvI
itZ4UCtYzqNWpz2f6EF2fCXkZq6eGSF9KfNeez/aHiD7uZkCrD3x4UDjmJRCtTgdJN6L51A4V9FF
nYhPk39wEOx2Od5ilOEMn6oXgqxb2dP/KGm9RuTkmQuPEFoR29Fr8ue4HcNquagh4rSSB8IVy5DY
FAxZ20jEGE0ESdix4rjDN1WDLyAuezrCQgDnk4V7la5/djcAzUMJEAVM1HNr7+B6DycGyTY9zQBx
Uz+rCSHkCQixY8wbqDYAzPioPU3ONU1HCogEaM/JXt18B9Lmt7Pz/rgCTYLs/LDOi//DjPVfdgzU
hse6d7uuPyeVxCR7WVR6jTnlZrkQEg/m/X/mGOCqUQkiFhlm/SBIre/g5LlXI3/vdVKipbvdSIfp
SxHPgssYCJGylM/nLo9HQVKIqfxR/gbn7aNy5hINP9e4T6oDRArPmijqRCoiRttsE/aqapLM8YUf
SMBVv02KB1N8sAABO3gdbIAJfo0qE0t621HxQN9MKsqXRCQpOqlfKKYRXwSzAiTGDIjdOpfCQc0Z
LznVYCtCgoDGTSU+2BH+EUtjj54FN0w2bYn+/5bgrEQzmr5Gha9acr1Ah5+El7fWmXCTAdC/l8u3
oT51FhXJwmzlfRIcZ1SxLCU6VGq7eYcj2tsAi1jR2mSvoWHZTivLbwtV9iiUrsbINGiiEz+Pa+gG
OeWrUATiTh5gjhesUB50FVjBKfN0uasFA3VWMgcPL8x/mBTp/hQfcaRiDKDZ5TZ9I9+iUta1sZvw
DoNpZvd+B37EBiU24rLV9Xv6wV/gVWbLWFRlu5BfhQIamPWAXcu0mBnowyZRk2MhuHZjU5d/EZ6C
Jhzw4Ve58WD00x5hGU8Pg3S7tvYq6BwFKCOVJIwEHtG1RhlHr/lGa/kOtkgL1F6l02sZOdLJZAvn
YHchZSO9fIVcE6hWPl/pKE/1358Fy0jq6A5vxmej5E5X4LOJe4u8a8svkH6iPH9vxDCF0HnYpynx
jE4bRqA26VpYuwYQKmwEdRcdNQmuL9WrJC9vpNsk7SLrKlCArVs8fRwOyxzjHumymCbdOiiVaiso
Inb9Sp7ZQIs8A+h5SiApVQX48QvrTCsENFaMWLlC2GQY6bkp+0G21k6rNfErto/I1FFUipVjM0P5
8CZUJlT4y68XnKZJAwQz1eRdT//zaFHNoUcf2j6R6RXlgjuTMMwCfL9bUZZpn1VXa/U8CnUXW6eu
905NJzIL/23tK6WFG/lAFNVKvPaYcF5ZGmd0niNRl9SSuLn9jJ1FSUMFayOzUAsrrbhmx8CdwsXu
DfRi4h99+9TboI+C4dH82/N6DNGdcXiBMURKR0FA+kzX6jh9BCgXgsoo6g+0joUpTc8aCz9ZHoh3
qafOAXqhktR7xCy78XlPJYKd6Hnr1pFNYmNPfrJrsHeN94AccWD+cPFyx0BZLW8rSBxDTqrFpCrn
BMfFLbLlbSKbK+ueG2GmtNVa4fMYQP8t8Lx24eIP4qjRTgVKQmWerNwA5/7/600Ww7qjnFu5XXPQ
erJSc10T2Vj3hzlzxJ5B/pq8y7jBadEdgrqj24U6h+zP3xWHz06tYLgSqBd7jRFeInqC0G0gLxFo
w7pHlwOq8h4MwCr8VqhXpIjLs5pcOQH3t903xPJIsRy86nlNEYrpW6iNm5Ij3skX5irc+0zjJMXx
C7by54Eagg1hlul9xvjkIfMscork+nuSvIM7oRXwZQZiSWJ2s5x/briwZGV1SQSJzwdFJD54lF+4
ruu1w41syfAS3CXdTMLNDNNmb6QP4JeyyAtV9qKNCkj5eI26VpyrTYyuPj5oNrcpe5APQrGsPopE
dpuPzrGMjYQN8t3O6CnWwI3ekBkmhoZJQfNg2iM4ziPsYfTQNQ3Fg0/SimSRVP1jG+eCSu5afPeD
KFFmGIx7mDYZa9x5Da6Mneaj1UQc+/P3Q6k8OQToFBajWsu10H8OtmWfbZkX6pzc6ykZ0m+Xa0h/
+CffXgGuApKrya7E+FItj8JduGMGcair7LR54fyo2ALTwEx7jv2zR5hQ+GHbhxsvjo3saXf79m+a
1CX93SYZc6CFfA9jZ119Iw3wCMxUPqpI5GucQcIhql7J5tGmCZxRxd8ha56GV94IWI6LWSOZxeMv
nI3PCSGWA4URNBSuRmoG84ot7bT9x797w83CLYug2TwSAxzOCzrh558fORSO2OvSzihCbNCvihzC
i2EF4575GstcDu6CAcLnxQGvOE/XdTe8b9fOEzdMox/2JPLaHngiAWk18kDKscJSxE87mkM4xjqP
A499I4ewCP7sMQprgaJbgbFgoLhaTbE6vt+0gU0IWnpoiQzmvC0mTswuJ4SIE34IiETF1dwFUtyS
DyumzH4q6gdpUy5e9hen8S6BHC8x/qLbOOAczNfHCS7cOhtoXizUyVIoqnkry6SsgVABo2g9ueOA
i9chXskWzXecjt3kV5aZ36FAgwSzaPVLWq5In4pq+BgTwWoiiNPetacZb3/zQwbdWj+5dtIwInUX
lLxNPhUgC2aF77/M5tZh6+Nw/aXUy40jPLyWOuVr0PQOqNmScxxSnLEHBpNceWpd7qS7GZjvzPnu
WAcFHbKD+vumkmLcydQXhgra0MXhbbxIVZ/VwyCGjgukkuAnGTHvpeo0KAL2xWYdAo+ETmEd+6Cd
XG+ik3HZfocKGkaLvaIcsua9vi4B046RBTEC2yCWnTw4RGYUxi+TCGbvs5npp8TSdthBg89aZmp2
ZEBe71WcnGjJ+Z0FyIHzMF3wTJiwtqdic/kKEAUQVl7Fnt4xPhtT2rQRJc0obOVMzyr2JokPYUOZ
7mEKo9RI3h6leVQjpbqzX/YSghz53AQCpcYjA/GYLFBP5zVuwUmhDF6yGnGddCCaVyjQ3/H2QApF
HuM2zHHpnzOxb5ms7RAXXkvtxtSuSwUfCkOCxLPH5+NVR6SAxrO1rSVRDIhovJx7F4NzOjGECSRn
ylreW/Dwi7IIS4HtZnQBAPqn0MLNW5U1IN7xV+n6w5ouWYMdrfKilQHvp+jz/wvpszpKbihFVS+5
iCkEyBUl5NDVuFUm5ztze3UOesFQDy7obbfzgmYuNaWU/5bZ/y1pTpyz3rVKgPW/HARnPpJz5e0d
GybJ5KexFPOkvbXh5xy6ifh6QXjsnNPjVAiuT/vS2CCsMG8RTMAx5/zFhCuz2FTWLurOJ32uznoU
ZIVbS66SzrvmL2vWh5dTgul5ZbZCvfOtre1NMYaIe7dq2KhbfRPwQPIcWKJqcoZvaSUnOmGHW9vm
aKzokVURcPyGWWIIZAzPIEZqMuqX2ZB3jQCqVhuw5ibWpuw+dmVoFePOoSpi6obp+ex7k3sfsR9O
C0DnF1AjGFjka0u59tcp1TmGRpXofpHesOQdXkjnLXSlfcZE7CKJ+xICOSVOXUyaza5iV+hHxCVC
m7QTz2oxPomduiLu5jAkRMxeLE/nJQJJ6P4Vleqr47gOSvcm9ipUgOibqq77LCMpCPjPM8fHDQCh
yvEfQQL0Wjx7mPfQQWuAHRaegXId+aRLvleR/P1axE/q6pb0pert9nF/eMdypBcsRvic3PxykHEq
hETt/hAbA7bixPy/KzKISmJ4SzS817D477fFT9gCjt63hSNgBDghYGSKS5AXos9Vn6Al+tLUI7lQ
0Rqbezg4sSsHByqMrYSW7hJDPKgvSG1DmtUw+W9T/YIDztqc8uX7Fmsb+6uvT2PmWA6xQsJHUKeP
F0CMAoFyFeGu0YvZ3Iuz6efYnzN7YKwcs5qp5gpFn8N8lslhVYVG9NgB0FO1jkHLgZfyZ/M1rump
i3kUzAKVWa5YEQKa3fdhknuR52aWxWc6OcPc8JmxwlYvl83kuRC4nzJlQHJv5H4gR7RXLYpjJRjL
6LRYCy4IyHPX3315SuKavvW06X8LEQhAp/a4eFmecEAO79zBSuLDcdAi1a+eH9d1QhTOmoNxYuRp
7iHcjE8iawbPEeePlF3FVIH1KHoHJw8ZnQ7WXUph6bN8MBLlTr8M5bSm+KseZoozo1Hm6L1uJULX
6KVekFEBIJNLLqt7BE7w8rzmyp/UFRxwGfFeqEJyBEmDLNiE3bzBkuVe+uo5h2NgD+6R5RdKBaWS
o22ccsPeO1aVeX/T4Mls5OpUGF6rsVHtEnNa4Ws+axQyQIpDAF7idcRNZEjPZziDw3Tig6+cq/1d
uYKIY1cqP4N0CNfOVCKgOHCy+j9NNmJ8TM5QxgqkScSTBjM+UwzQola85cThlLW/rEy6m8nl1qQx
GE0SJpwka2Ymxzv7wZ4k7zdaN6MK5o0AECBFWvTfKvSjm+PZP2CejnJyvxnSOiiDfUZfrSv/va7D
w0s2DUiVtDaoZ8huyfHn0JgY/NHGmCbL9auDUK4mJg0YzkcPQMas2vh+/Zw0alIJogez54U7kq3k
Gr8KoxK+fRZvzD+1gM1I4kgGK4ONcG8CIOwFrSoBVTOB6/X56sJUJO4cVmE2TCKMterEJKxyDo6I
7Dodf5YOGB7JcOXOTxJmL2S5H36sa8WLSqJvZ0za5yAlXz5lKw56ffNCnQhdopPu8WwOXd6OOXec
lkYp5fn7Czs+XXLPLLGAmw5U83/Pq5/BhlS0+bmzJ+VxWDnXovI2KZwsYeemkSIrnhOiWBo5S0eD
e/Cux+vsVJ8R3/C9nTperHq8UMX3+CY8Q7zvv2SrU8koGA5nYd3rQvneEiclkpL9ALV77ltYTYXi
k3hyX8VwAdl+TE9md+xiFMbbpWcDg8iG7JObPZLaHmqTCLzJPNSHgLOjVQZ/k8a1MfgzjuWZKtZJ
zeiIx3+gVJ8Y0yDExKvv0LgNU/LFRk29IuZc6JBQroOPrVxzMAKG0+icVNbQOwH2W9G60o3E2HVo
NMdFXM2/KAwapfjd8hb3LKncvv+5R+4qc71CpglEHUlE2KnhGeqt5asGmKIEumKcu0/PjUGn7E6N
Di1ri1IPWylpyf+d4Ad5bD5hVEbXbcf//KuSC7U3x82SbbkqVpig5m42H45AFUEM1GgMWuwN10vT
3LGyY7DBPwxbU8rDnIqRzJS6xQluzxhCXk4qRcsPCCNxaItdWQ6jLtbKF5KHT9fk4Jo6SAxH2xoP
GsquqVgYo8ztotmebtZPDLzMjWUlb1f3VEklpek/WW+25vnQGRAp1ECV9PVbQvl0DVcWDqLw8uOY
LzE1N4qeTVcRNcwujC2IXLougaaqJNuU3a5Z/xsgjHJM4ubxmp/u6ffe2SrveRZmEt6T8USKt08c
manZCASD9X0FBhAwpGZiJzQ4tQ3dEqEo+x9AFQJ0Qj9uS323wCaewfHqorKOduySUN8+Jh7M28h+
vGXO7IVwbgwwsXitYeSjAsdSIU0v+bEiXhcl/OmWOPXuJPbigBXaWuGumu5WiO/9tZ16D8/iaxzu
53xovwY5od3+bPyBSLziqrTiHTL0VQlt08jU48f3W69LnSiD5upiZioZy8dT8cnkW0bcNGxtPtN+
h+EMox/TaZ8RiuIHD8Mh3g6f460rX9M3+XPXF+TI+E8IXH/hKf36KkY8Iz2t2Mn1rLGHskZpZK12
GbrBG1mmMoaKCWcV3TlyVRE+gk5YjaFJ+8nf5fAazn6t63OMuoDVmUfSyFAUtka+pCivRwArwVFg
2TSX67qhxczgCByy4cSN5AdaQsHVr/z7ojVmT+6MZls3r2WbnaK9hT7EWRQaaVwhbSNDQWNSTftO
wjNPkUHQOJ0RkmbIP1lVTq9pKEh0CR8HFuep44o0C0hPj5AEEGV92Jjo4H+iUT7gFCYj0bDm/t/D
ZhzdqLR9n2csIzEXqckLwSAce1jKYiqzTOvqfOYV4Ct9tECtLCBNUzmAvtAE717Z2Z+yFDi/cRZl
jpSX1WoIrlO54EtS5TJOsL5F2s0kKJkPw6kYC//IQ35N4vF7mcSsYbuuqSVmzBNVfQyDzzjVoBWm
cGO9e1UV55yhW22OfxG35dQgCwTsyeEGPdwvhVhI+RGtHn38QUF+zl3k3YlxuqA2uJlsaXJmHAmP
4Fnq50Ik/2+sA49pax+zxzblCUL0X6ADCYUOMjMKI1BmzCks1RSt/yw606orfcYk6K96/pOELcGy
eHZm41Iq0LiIrOEMgehVz+NAdKtwo4QrLXkNDY0P7gWdgI5q2r2o8QeJzmXZFtahluiuivbrC/+7
flizdJv2tbkmW4twnYdiNxB2Pw2m2QAZEjE9B3PaO908Ebvc6mG7hL7+ebI1anUXNfhsjMW7eiIM
mtc0u61NF5PZQ+CorJMPt2wg6M2QREDlSUwzFqGjOKx4x7m2mM1+Pjq764VrJhPSnRlZIO38w413
5038LgXCEF2r0rYZ+6/il38ZMBl8BP7V5QtPBY4WlpbsgcZZHSNeFEFVa0vD5CHXmjyVhvi+YEoS
yXJfpOJgLAubrQaN0DNRBUeZ2FArmSmlqgF2cCZyPLMN73345+G3WlDZi68HX6Syzgwx5g2olkwa
MC035/qrm24MaFQFyWUsQM2Z9GGV3pNrT5phlG7x8Ca4sZ1ALqy5RjNuXKtvOyimU4Jf5PvCwabZ
01zLYLZ7WHM2bEMnqrZtuF26d/Q3hARZN87RoURx8PZKEwHh0LUvOGwnU9Y+dulhyKZL8FSJZhC7
VqPmMdKxfvN7GlDQZzoUEpN8G62MXYCopFgtCUVFmkXNm/HKnh2NytJP7dQJg7BG5OF6gZ2lhpIs
LkYg3GnxklkiNJ3au+90qbM+bcpUefRkzj/oiZZgHvolkCs7owOwbW23mMAGceHyV9QLa1beonWG
ii/4di9hsmAHPlciOWxVPiCKjkLVWRsV+3eQR2ruxdhSkzspP4A3bpvvicJG6P3MiuHsrYoQnk3R
UpiiEkjsSTnd/02fy1znFHTE9QlxsPoDoRRBY6VrlIz4M4b4BuE07aIOFfLoaJHLe46ZUD7cZZsm
XodTzixGqQFoTTMLHvCQLuwkn5NPTi/TPzCwUZFrDwW9OmGnDTIHQ7BqeTac0FEQAt8jiE1yE2Jk
MdX22qv6qT41VjLcPw6CoNWh4rpgkRWILePZRLWJ5JBLjKDQLleiS8gGaldAs3o+e/sTSzS44bv1
ABtdGJB76zNjQfChgEoRHOggzibpfBf6tOEc1CDlMPUuwhGtUENwLhcKYy3vtseI7YHf3Jy2II8f
dUyeBOQDv2s3KPtVehGpqDGvZnXV8h4o2FvX89ngh8yKiGlW2LqkPyp5T5M74JZrueugorF2qNtJ
ZhwDa5if1iHv593Fq8zF3VdmtkOvL0ie1SrcIhViWOZdzENzLf6TouegspX4GWv4jmiBV1Ji482N
JyhOtbf3USJyOvUk0/mvqHy4OIvk3OLy3gqJJzGL8SEDKb/Ty5sx7VoIXj1FdhOr7Ne4uYfUd32E
GS3eEz3D0Usk/OrNP5tySam0vhPWHMMFhxh+hBD+moi5FBkyuFuD/V52eiBWht3rVQX1nEhYmiva
q+SziF0SrqHiiZzrfpkObC7Y2ucSuGVZq7ch33J+y5YVKtqPApky8ud+X3CS79PP4ZDXSp9nGlO0
O72YaQwsRnMrVnMIYCVRljux075qlzZrX4CP/VT3iprIDERtwSOsxiAaCt5f26spJ2z7S1+tZ4Q5
adgymaPMFZtsUyaAYpaTexw64VEwCY8zbjdv5ZtNCe+IozLNmb+fqO3vJp7AZmYmVLpAfVnmpabT
RyghcYIeE3jT/tgDI9iyglsMEg089puJbHJbxRBiRF23ZUt/4rjYwFo7aZKXjjfYb5OHAjecDZPb
yWFeex71PS2JgIpncPxklureQKEFMuad/t7hpGKDT7BbqhVX8rvWP54DPUiZHZrnMRBUpnZzQbSM
fW+a79820CjfUvkpWvetIso/cmulP9RUKBcBlWr+u1nOXo0yeq9ROBhfinyRzZSM/iQ9jRs9boVL
gFgXS+FaXs5m/ue5h0gflXpNFubLCVsMIZ0lXltr9RxssOOeS1k3/OiGJcd/oVlItntYBSjcg5nt
TU4AMZiSf1zzpu9HaaHD8Px7yHt75NHv3xfVHzUPscfO6KU2XY3XiNQZLQGYm4kg5ifCC45gNWAP
aicLp6gJaspisGJN+fQq+tg4x3s6BbfkcIXKCIxfI37hUIDBjhmNDr+jDMgBgNZFIj5AIilf3Fy+
/1m5bNpCSYw/YWj3JtmGuc2khTT7XbFqFPMGChsRJQLVOB8SxV9CS8iLT+WUZ+rmxZbuLx0YX61V
L1KYcllxEx1HP5mtA51TDoeMa+4L0GgcYnWzEeqoWW+h96avuibh5NSGJSKYXuqvVkPIbadKCxNq
3DE4jBew1sEYzwNFeqU2HbM/as3mED3jn/p1/DR4cr6X9xNQSj/LwnfdA9ehfP0z+Lm9WiubJtVJ
+KbKin0C5SkhD+oPpsQqzEUMCKHCF8pKM12LZILSsYnjJKqzBU4RNSp4fYIEKCr9sZeJ5XC3tSen
UbaiOtRh6JB9r86yc6QfShUgpzZwBe1VYbekE/VJSopr0SsWPXRvvGBkCSz1tof0hSesr6Bh2Gxa
smhPaxDf+8/zuIbX+rKUZnIZfJfI+zxH7tbh2VrdJzExk54REr5Wd2HyUG64c7XAz8edEOC+s6yX
FQ18dpzaeKimT70VeHl8tGY1f6GpqVY8rWmY0+29g3EStB/9ZADp6mOV+iM80CVLJd2ypg7pjuai
cfBc0X1vrctZb2Ph8OtVyKagK6B3Evx+SnGzjsxHpBHh28xLmUDFuYl2c/SuZIWvhqBl6ge+4ZpS
ZeIRNRunf0tI62rFVGbJxruiwSeOsMq1hpet1/gmHDrTqrLmvRRn4vO7WmiZF36JnUnDtGcmDsrD
2wneBuKCA3YszcO88MIg0NSLjAL1UsrU8VBOj0ivqNUEaKIqLLDkEyZf+uX0vNMZ8rBrJ+bFCPtJ
8Mv8xJvuVk3on+ZrlXQL12jVpjPaig+MOaAGmHJH47Em1yq+igM6oOG+3mqEwzmOUNx9YonhbB5y
aVqcW4vI5KrbAu5OEtgys/o8p9inY3KdXgV93qtE3VqcRiHYv7FrqpLmDZkDzn3jBt28ZYwJr1yE
7+0srJLNXSN51jLitxuNeEnRR3WYtLBl96AdMY3KkktFZ97VQ1MfeLyPeja1q9mHD4mHLfzTWN+5
jEt8JaxojDdrHsGW7vrZJb2Fwgn17Hc4cQqG1rf1FFkl3hGWgRPqbEDInYGrRIqWWr77kgDNCjgN
yKv6ucnf8GYzYdnEEsrRekNC2x8K8W4c27Ez/FBScCjdve8C+kYlIS9iH0dvB0Mbnd3LNTLFUsGD
MHI+PzyVLeZfs2fVrk9HJvy3wsCTwa8UpbbiSOjCZZYq+0EjBlDCJfNC0k2sLvF2rMhPP+LWad+j
BvZEqzOVCQydHn+BRXZCHb1ulraqpSw02LSj+CRBMfEVc47pWJZ63YCVZgtd5vgpg3R82k+1WrPe
HTVMFPnRJKZ5M3ItzjLRGXF3bngXdkjRfaobDkQlBg1sNLpziBEN5idw/Hx3RShuo/EaLaCHxvfv
Dw8bp6z8QnR3ofDv2ItDoD9I14u+DH327q3FKJzo1/4Dj5PUHUf2595LU3SezC2hdre7RoOmmZii
m3AsO/uEDr1nWDHEIMZJqtUFAILMI6wy0A7MtivMQ4wG8ao0AqH6nAl98IxDjYm0q8fvTCHK7V2T
Vv+yghl2t4SmEpajToCclJnzsr81kj1P78aW+BeF2ZTFjk+aCtvaXFUnoNEdaiCp90m9kVlBGdYz
k8JzhLORtWv3z9qRZ1L3YPfJvIIWAq3w7y0Illxn/NFn0CH9+P4Q5t0wWfrL1krhRr6mYml5Kybw
UUD3FTrF1TblcXQH8K0245ryEovi97WEorR431CWoyhRiGgVk/t8npi0+SRP7kTDTkhI9VAvWgpw
jxf1xKCxxwRHpx75i9wdk/NJWqWG88xCgxenxOAuD3qjnAOI7jjEnvcWRT/mJ7M/GDAT5A2bIA2t
JB282MHgEW0rafZQQtIgcB237eTg1Fk8A2VkNrTZ4i9U+1XslT+y+gdrpJmtz13zKOpRRJRFGLk4
dCV+RzI+zb3vLKziBk+hM+0Mziwv4FcAZSaU5uc3MO7tcjTZmtlk0ckPX8Hh9rwb+hYfWqkychQt
3RXJs7MhkwjSVf3sbfo+x/KA4TZxu9/5NMEB4Cdu+TCqV/psBcz3LFhtlBoHFBxURp579mVBeekp
O2hUCt6t6F0iziQM8ursUx7sU6ibGfOZUDPwQ3WO/cut1z9eh8dZhYQpDH2XWV0rZzAuWSNYzycb
SO+uZj5yKoHGifXv/BDyEI4qZD6h/pB93qRThnxCX7yGVuUpB+UO9AKhfcGqAlgmGLP0sdEBQOhm
A2mr3ZXQvIoWZWpvOgJgyo0X4LTSHG/KadEd8iHcc/S/9Qg9+zkFvXPznTLQviMpSYiD6JYyT25f
X8ggX6/aY6h2sAIZmmSHCPsPHCgpbrd9OjNaJfeufmeeZCv7fzjIExhCVioH4aYi2dVuXCj1oaGz
yc3m7sPuqWOeMaS29pjn/HkW99U2LgpJ21HcRoAGNucCIe4u65cKI/EXphZdcp00ZK7Q7VteHS8w
or9H8ldzvWYqVtt7xTTxvEYAJGAmgZHgip8HCqfhJ7ASXTLpzwSEQd9xylekN1H4kDIB0x3OOSUu
h09RDj5djzha5rs7Et9SoZh2JfZuKoVZFkrJx1H9wb9uJNoAPtH7iGxcF77NnfbvpVy4LtXDEeYU
E+hHiPToAOCNsUXqSDe/pxSWG+hPNUhPM+9qfR8Cs4qJ8nsyboYpDMaWYPjnPAY97qqYCKaeq9dU
BqrhzmncHPfzw4zYavWpXSJbGf43G27ziIgtcJkrnwj8yot5MkLlLQMfzW+6x1xTHHyQXwPpg+dm
+bOshHYiJ2+6O79hAYV8RS6kK187MEQjT1EbyVPI5MU+SigKt7qsoTtG3K2X3nIzj2rTWDH9ptn6
KbW6o5OeB5irKmgQg7+4/03kLiy69p2Fx3esp3yddUcvysDjxGEZnsDuqv2HKrmOYWul+oyE94lh
Y3t/SUkQRqsndtoI7nMI8ZLN6KGfuRAfxFPm5IPrWgkme7i3wWaUHgnxigy3w425z3V7fq8sQ4eJ
i12g9aGFqJUC+14FqDwW+KDdCmku8qlBqHPwF1DTP2D75aesfAz00rz917fisrSQWdSUVbTt6HRK
ErObHAXwkdyTGhoFo1yonHkr9uhvyPwRGSxiclr9NMXBxIkF2EeAr/H7T2r8BxuAtPKANIREY9Wk
/eEAc6SKqS4YuhBGrvzJtv6vNEqOKmajoIC+56BT36wFnour94qJKz2NWTUCfRLLzNqNhLXMSUY2
kI8qmbTsO8yrAHR05I0kwkHtd6BvXIWdnhOkhhhXtVglqJ0an9fFFtsBjTUnXGc34XMWwd6EsOI4
IPvAysL7q2iOLtoAHHAVk9BP4Y+mu/oPQZq0WbDcKiX6PIaa25pieRGLFSpef8ZAfK7Gb4AcV39g
Z10L9Ybb3VIuHB351LEIIY2AdO0GVuQDv4x1tmUaD+HgLpnp/2yOhc3XKIJNmAdFC6wELHhwelm/
SS5WGpKvwEdfFwR54NF5WHqOw2t56cWLBSXjsCsv9yFP4ordYkSihww/26kTMqcO3UXXX5icJIdA
l7bjbQOiKl5Mw7JM7NeCsrVmsbffZasw8Y+c57fU+ze51524lfQd+sFmB6Bu0SpsBDvz+gWWZ6vS
8aWzFqATU12BH9Y5dGLUAGKNnZkF3OLCIGLVRAMQuJ5MBa1tQ+4rqU80FAF398CQka1S7OWmf52c
QAIoVnHZkfDt2TDGSHFN+gZLYcip/r6x4mQBgTZpkJmSrGItmz02PQUROGWyk4OLgIyK9jaWnrj0
+fjGR6n7jGfORITpWi55KoDXLLGkfufftSiBgNMVx94F5vWGwlR4cQ+UNvrmuslmzat6w7FEKpyY
7UsaPdFb4Jk2EOE0aG2NDbdtiCnv4ji1XUG4mNwkmX80LhYUUhG0VyqD5SaRY5lJw7ity431HP8H
iqbFQQJa0vMRofOf2KgUXRjXqDYlGJC1o4nd/AJKcS6YlqRWsg6tloezOkFd65dHfabGgSpKWhwg
6lR5bpRDUse5ljCE0Qy8icEpl0WZW9IY0zixFMOK+HCh4MLpPmZuj1WXp3JKsKu3RXCLQOawdgu+
aV05TIY6+sexvqUsr/FEiv72ILrTwRV9S4moIY91MbHIsH745kq9suoiAxZ1HnHzsEft6KqesLsb
dDYUJOXC/dvLfsa2luVfHIySlhDVEarpwnFJxIb+H3757q49AZXrqaJtjkMdah8dWvV267t4wcti
miXhW3PjsOGGNwkes+U+cDtrCIz0eGGpKaw3uTZumbGefCrmeWNCFn4vpHWY/QcmLxEvBkTlPaJG
zk7DOIYx+asfxRyuTTMBQ+TASy6YzJ+q3z97jtC3eIKQZZjx5W6iZvmgFlBYI0JrvpL83JUK00ng
UpQfsO7ova/EhSQGGDFontddQe7xn7IWM6cgm8vQ7MXRShwlvAwYCH1fHRqT9QTlzvWEZ6EGc2hY
61tswfIzoV/syc50Z0xG+55ccXPDHp+lstTFgWpoe60Fld75e305ovwGGdzv8Ue2E9OfhLxxz/Eg
qDrF1AEdawMYjf8TgwFnVWMxf+ii+Llsg6B9Uc6eKJCZATLLq4IL4pylPWnzpRqUhapR2UFpr3DG
z03kzsvVGgodSZpcJPX/bbGYhaIVC6zmfepcnqaSZ+mVPODNAclJTgdVDlSeWMOQfA5s0ErGjKgP
o3KMmbXwvKtLFRO/ESMBZtAxP4tMvWHfOHYkGwN2iCVDdJWd23nuc6OQSmPOSJyXanWUi0swQ7Zx
A4XwQtSEJNd1l1n0OMTTu8QnkFcATCIEpASpvpnvuF9QpAk+7gtAh3xonp7dvuG1OcWylkbJrbmz
Yo+eCo7vEIkzGSk6SfzMvFdDnngf5GpnbQgSJtAckMCi5f8ueg4BZL2q9mqtOKn3tK73/ANsOtXL
B0ecBg+5fJfd0XG5cGu+4KSVTIhWUcQZRNHNG2mtwQ77QB+lTmOwu8An8XqKDise/XaXDSp9HE69
ZhTf2hk4VeUXAaaN/DL0f7uLlXBWD8mvYfB9lle24WhaCv5lZt8oYKXYoUzaoPxmubieEjaFtdeX
5/73toMQTfOQmYaDdCk4ulf0I5E5WkSG6zagRnbzjo7oDUhcar3EYAbUZ2pl07mKRNBh9UZlXsOJ
Xj20L+O0RcDZwE8Aa5fujLEiI22R5qGEQyUHmeMob00PYgg8x4SUNaHTzZoyJLrK7kXvawrRqJ34
UoaHywmNot3MaITud18iFeVoZs9xLpM01+kCl8iT/Q+EiniesD268/wIUKEKOdlMoETJ6FdtfdS8
GpUxRthMhq7TQ4YV2BlFFWd3QykL6j/n7Qscl1MCohwruc4GGcO+9V+h63R2OIFzLZnHbTw1Pp5p
JO9Ap+ZsiknyN5KiuRXdxUH0ZuICHQaIj2S/0mbvlhwfjAEfnqLJjYg5WJ/SW8ta6HIuWWtHO3zu
L81sfg3gL9Eu/rtVoHY0B/szYMfEFnANldlfVX+/rGJeqyxzQETctkcDEL58JAWxX5Eosiz43HnT
gTxgLwAwiD1puKCxmupGCSq4rQ0Q2TblkU6AAXdUhMPI3qdrkXJZHDeU8cajPvM6Jq57iiAn/dbD
jjDuosGzyok/Adf+ehqtuBCR72S9tN/FApfbDBdfwYtcwOLlLQFpkG0tJn8gTzBPke9SxQADX3uB
FWSvAJ+6UQgt56YPFfx/glPCryUHu4RvLfroiaBtCClyXk9h+BwoJksqIiVLnURfk4HSUaDHziHk
27cVY8DP3FSUUn32zJ5Duo/JXFJ0JfJtLb0hgecAercFNVpNLcjuU4azgawaLerAraEXMfLrwhP5
ocmeg8+r7nUeHBiUPSA0n8zEqbQOGUji5KFvjDCRmOhE+QCP/gsSNkSEgwNh9fZtnBV9gd5DLVrM
i32oIWgDbhB5frv02M27d2hYywXV2sUMclCoPFTXeQbVFsU7msnYvb1RHkeAaDT222fY8g/u9muY
OIbv533YYsGfH8nJAtF/IZNFD65e2geeZ2cgg4uFkSt5bJAwA+nHoGcwjg//wcQmvuk9JT1AYox7
D7gMzL4Z6OFrAZmvNKhBA2mSawnaxyiAp1pmEwT1Y5oV+TiML/DO/xZLPWjpqNJEJjsH4EdjQLcU
R85F28RETMsoq/ARc51fuySVFnDkUpX1Ssp69OWDzcFTym6kDDsTHhTuyObp8So+aivT3ETms4lG
Q0/MghCI1Y2qgLRgszLZ+LgB7N9q+ckRH3edekyLG9Rwc4g/CLKHmk8yaQ3QaFt/V9kOgDLto1ew
CnlMxaE8nBNDwGcaJEPIJNwExF7SzKlicoyJtCnOIUTNoWtSwd3OpPGeRfQ4uXc+rAdHiJKjf4Yp
y5zZyxhtSVP3Z+YtIOPFqYonEtnNFkZSd6ivL4FrTOwMDWIjiH4VBEwtIyLFmtwP0PPpM1MlTIQ0
zKJ1WaDpt3hCJcTjWzex9XCn4cAkV8+hJuNtBmHGVgIgh1MlAXuuB8hByM1dliBOrHC0GIr2L0O8
DlLQZbUcSy6sC6j8OeuPQLt48xHHfFYSZaioR/zdiwRs3uwqmPvOj91GulBPP2YYl4wFELleZ+6b
UfkOTc/BPuQeg4kS8GyGeyNwiv2X7XzAueyi1JIKLKKPZGxLiu5gvelMikRJ9FpI86swc+S1t4O5
sctUGC00gYBf1y/lqSgorl4TP+jd1mV6XCn/CPW1kBXXfAb1OPdLKQSY/aBRMsrmG+lYz63zX3oV
Q0+f0iwQqH6TV3J4C2LEj6dMuc138NdiBECAw/STCnYtMpMigH1QAPC5rb4YeavfVa9mydWzX2pI
kcj3losldks/4goR525PjV5+325f1OIOrRMDLQ4+fm4QHJ0zbAGhTiucX+R66TrkGu0Vl3g7oKLQ
nFlEXBPOtZiXo7l/zvtR8OPgcInXlptITYydiGqlzKqAmnLGIX4N5RhZPDI12t5LlpH6hmTZICS0
Zni4ImqOKU9FPnG1za2weREGg1whGr8m97g+uFPlCUiU4qZoNtbFKLLZ2t7qrArj6XX8lwEPZsiJ
3GD+KNUgTzKhPE0Iz7Bx5YAcZzB6ZTFcCp192jbHMaMHfW6v23ivJeI2K/hluzPRRUuyG+M9ktQC
ZmriF58GV+z3Ri788Nt17pzWE2XSEG/FZvZzQ0n060TCaCslV6fA6AjyKRxILwN7LEpf1GA0yRq/
ifvdgpy0dLLD2Cf4eEsEIt0CcE6w4PiTMV0ApGdMY5KZhITNnhlgNntJQbrKBnQyMZvuAXhreh3k
/5OP99F8+KxOhaWfRLF3y5A0XtVuNoomQbTwecxy9Rps1b0ImAsCja8geaFMLE9M/NlF9BnUthJ/
z3svl29irVwafyXahWqLoLasrlXyGYlUz5O7whWshe77NQGLnq7NgUIs5jiIzWowFm6bMrDQBP8S
XLreuW84id2IY/rwvtlDJC7/mJ7W0cu8gkjcByDbTw9Um0WWOHZFR1v04DHF/E82hnFYy9ZrpN0k
O9EPRljw1VKElJlmw8iEpfikn7fbthB/XcJlilNc5kVMqOQVVLHnpW35Niuq1d9YjFhk6R0Gh7mp
XzltdhtZByosDUq4oVFiGkOclrYMm+8Cxkk2W84MmAkzZ0qIRXg0pZVhfZPGNHn68VGx6oplT4eV
HDhcagx7TPPKTmFoWaIYDZaMS/0KMsnQlklegfg8c0LAX44Uvtgbi9r+26qRAjYi46UKM9guGCBY
P6EnvxvS4M3qh0dBYeEsGqOC/hLQH4vO3UV1p4PuOvVAph13UDe4DLhCb5od85fYqf3Lp7TMJFQP
3piTI9jF6hrL0nY54NGTvoSOq4DtsxTw5G8t6APPBTGLRr/8zcy+7To1yTilI5BQvUV4WJA+4UMQ
cwTxZqz9xlyApS5e3g9KXdae+BJ6R5N854JVOeBHPaC6cbdoHaxT+/26xzVEYbbnHVERmMSSqE1j
Ms5zTaB3swkSlJ0sxbXOE39a77xcHb2mJp7wlnroXqxlFr3PDZUMUQKPxjAaLX+Q4jG0/PWzlYLN
KehQxSnunn6A1nEH30Ir4e/OmR12XWstJuTqnRO7iMMiuLO/ErPal8h4ZTZk65OjuRylRLNfCukX
kjIRJI8aJsOUsVasofe6MJ3zzWbyZMFCjtToAWH3iV4X/Zw8lttksUiUGN35H4Q1+rduKqLwROzH
GikS45K7sXgdhAu7vc3eaDo6k3ZzxHXGe4ogQzUwSIwS5skkDZyqXz0+jSSwAgKmZXZsNQ/4aMx7
FqysAPUHTd92LL6ZuoUjgSENVe+BT6miaTVNnGvV4tc4yoH0AOA54sRVze+UPpUKMeUzrP+Ptj/w
MEiUC3gyMtuhm5mogXbvJ0Etx4zYKYwTB8G2RO8emzIslPAt5jmTf7LlQM+E49guDXewLHaHycy0
sTKjFQIw0mTlX6o9oBg5Mr9VTQXyHZo8mjUc3PL8OcqOoRqYW8UEa3KTNlG2Iw9r7T6aBuEfGDSU
Lh2fTmshET99SvvpEa0nliO7QRrnHgLuJD+rbQwr5ZjjWayMjcCnb1Vw4ornxZwMi7rg0vZDYNSO
ehdnFvXtZ688FdF5DgSEFpDmQXzYfSMdJTZfHMBQkiWQQMDSVfY7JOI95M2QzL7P1NXC7/BTMzJv
tWoz7MO85Pzj1qFvCkkLIRXiT7qTYV5Jz+kXgV25qat7V1f40LQ1yviM9uzl3nx3ZxeyRSdq0BD4
ZB2Fm7ZO2+0iIEcZ1FzCsvsoO/4g+FtFJXha0XSS58JkB5mg5bzyva8CDIXS/9e1+oJ2xhHMzOEO
w9cucuSNmx57etWUZ5TB8vS+lOgO6meIqORHsHpHzXUswLkvTwlWeuFFYtQ1Tunf//qlkc8Ayyss
typYWyWnxFEnKwBn+rpsBQgv+uDh1JXwcBrP3xrLyKHJzsaVO+HJIK6Lrw3aI9LVw9WBEUOZIEuu
ydNMdJ5ITCeRNmbr0hsmNKfZddeX85WMkbHO9f6tiD868pjT1ONHMtT0eieoGkttZXqC0osuS4i1
vir8h5xPBaJlqIIcl0SifJ1W09E0+JXlbcpcN2rVtiGa6FpETddC2/j+7xV2Gu3Z/lE2UUXhyzEh
NwAaGvhFXrRgpN8UPmHWOqEWYhSUDqOIuHALiVhiGHWZC2dDeTFeoWxY2dGjlIeEhIkApVwf2uEE
SWbOmyx7YemcAx1T+5SUxyNepmDBwdBL2mSFDgb8MeAgPICgDjenHRkuAXTOXDHvNYN2OqVQBNSw
v5j+IoBHudSfIZwBj65Jz8YTeG6WYSpvTCmYb6X+LIgjjjQzwEvwoeTpjx5QPras2rn/GKurQ1wZ
iCpxqHZ8TdUgizD6qk0Kbe6wsM1oLg6BZ11WkKhpEF7hkdcq3x7MelyUfDfJAeNvdWbTN4TdYkJk
LrWUl5EnJ8pfX/1sxASVVuLmaG4DjEIdl4tzpF8z1+ejK6/42E3atBh1YCHHxxYxFYuQ6zEW/08i
aYeSSrDffKIPromDsDke0Waa2EHuC4RuJA3gcDpVIj5/treWJ+IjRBcBddKjazZbaODSwSy/Zvm2
J2JyUR8DCVR852/Me3g2dtxE1JfF7H5uKr+z8eGBq8muA/8xIm5Akivuxvh+z8dnf+rEmpZzJm68
0Ygh8Wi8oDHWHOqh6MWKUqT5lQn5YtdH2CZBUH0wfy95PpoCW1Rl3yDqN7GtDNCVum7MLrrTDDX9
tLJD2b2Qdq4Fyqqu0FFbYg6PnPx/KKrgW2Hw1dA9J2EbO9ZN0LFp7cHX3a9XZLynsJDFDfHagSbO
24au/veN7f11zkmJBCrMfPDY7c69ap8vXKFWIO/i8eA6E1gIlMWrv544Lvbqj9aZtJOAefcqa2Ne
g6UJGcf5JUcimouBy4GCgRlCY//hVyKwOEDnZFPzl9fXYb3iqLwaLTWVDmflNk+3tBDZRpuUkkpY
oOHlusU0o3TMqhwJDi2J6rdax2n1baQqKpBRjJI5O9EruL4qDv8W0074VPvnn1Jc4KGYlzbxQPQN
uvf6MVfoUrmOQ/1pFiYK3bXJ7Hwy7fOV1hNffdNN4P7WFI01nIGnIphI1PoNLZA2AU8XWqkztu/M
wUrGRvnAy5/xOGunOzFCMMPgDJ6PP8cR57BSKuONzKCcqxQUl+wiY13cN1FENRWhQ5KWlkkyI0fq
mmM4hfCDFOhrmGoabhVXSJ4EYwwbKHflMI/Hs6Or6N3VxbUutD386TMzYb7W3Y+ttYOjqUF3R0fK
3W0q8gxzH6r+vSDFiaCMxFYIKfw/UQQHw2tj5H4zY8guXJ7/xtt3Q0WprQTEKKBOPXR21sqQQGw6
dJe+8g7LraNiaRMZq8ZtDdtaKSMcqriJLkztM5As+3lcfNkAqn3DG0yJcHESjLgr1kmzRO/n3Q6o
tDGKNaHTYWorF9PI35XCEDIEY+agCHb2s8X2LlWn4GWACHmyyT9jlDw3E37ndz1vIUR+Opf/QkiO
kruQVFi9wBrFv0cgotrTwpuJeGPibmlmFbQnVSZAj6fz6Cu3U1uiMophEGyVPbl5QK2InF/rcPYb
Lf5SMWGsTr6yWnZgUsJeaAjQbPo6QGGBpAprfxbTrG+4KHyVdNwLvsWrS2u8wUKCGpOyPsb+SSD+
RAjaG05RBgjdfxSqwuuXqQaRBk7kwmQBsNM7m6Oe25HgzBPKY2XsSaTr3uY5kGJjmzcKjKe3PVHI
x69g8myPZVktxBxpFrs1R/X69fZZlCRTgeuXGFrOvzjrJ9ZnqLkXvWR//wnQCggWLuo/WC/4XrzE
FQAxy4X9hMBKAGz9rVeT2vFwO7rVSaXSwQlIhVjyTHu+4UuSJaWPZKmJ8PR0UkfUDauZM6TXezgL
jtq9rCI+kXEw9MMz4Xs34sL2AbMPa/YJjkmry/IErwIKYHPdbiBCsEza7ELYPtdexzVZ/QufgUfF
t2NO5xDEeg141AnM/e97YkJkApGXNt0LRzrGFHVqnws5yPp/EhwCJinp7yaK9IsSWyQ0eR8SejXT
iaYdJjghbA5FxIVJwAC8tLTyeFqGHOxS1IEZCDwgXH5N0bXjW0YI4o0FPfIXDsiZm0NCSJiHjr6+
Jofc9AZf/SC5zH931YG0WJrrYVaxNOJUg0iOtllzJcA3Fy1ccpxJm3+59oEEcl2YshBCQOnR0wqv
wTsInsSHEGEhWxtchNGfzcyaIsM93X+74k0K9Mcxs8IQrAD16PTTURZJ7r6FQKHHs8CIKkS+G0p6
bBdYwyeRLm/ND4b+pEnFVldvbq6dLmOjL3irrhftj0Z+1y/Hx84uMTNILBuW0ePau71Nw1qDmRYC
N5ijjhxKgmO/pWDxSGMAfvM1NtHkPuy5ptQga8F/0o/jppZNg1P/5NHYUL9ojtRyUofPcTO70flS
mMF9HZKjIUs6HhiVDIEZ9alpHe4z7CmaWxPTxUbJUhZ4D5T9g1nFnD9XipxEYKKVfjEsLiVz/dz8
7YkpNRGyG7xH56FWTKHsrXqx6tjlrqcQLM+cDEPNG1LYdAuWGDRD/vPKfPpmLV0VImylJCetoQSW
dTYKz1W8YkE8K0QpsslPC9UO7rlaf/ZEElHLOYPkhXqk1QygX7G5XETH9KTLzUgrnIATpf+boDlx
I6zSX8wslvYfK83Xll3aQYFeJVE+94B2YJlN9SG3ILrLUQj6T8P5ZeqiErC/B8hwXkklo5uNOKmM
PHlZmO3+kLy6RyvoEbM3HM1UD1nVj9qc3EyCbLNMF5dQiKQalrtCoLZZSZCyyN60OoPq+aqxBLBz
PwYAhHn6hPHam9EvaHp8DXWsJw7mEPw4jA8ialC12UaEy4NImy3wkOJH02J1vfeRNMdLAigBfYm2
g6HujFNNwidtFXttRMuqt+dJBmQOU7WsbGhwvI8rXgmhX9YMf8jBXAWdh3LwpJ8jLlJqkSuAYwTC
+/mJcIy9KfURrwjWCa/16pqpg3Ho5w8pOs8EZVO51sB2hHaGm/sy4pByfQgSBUEZY0uJ7UG2A8yn
c7Vgk8TDOWlYSa4UhAfBulcKMKKdlA/h/rOXfmczB766JB+1vVVxvGQ+25NYLOtmwh2TC/LhMgI8
z2UeCcLm03fFDDjH5MS/dgPmcvjrhomwuKVcr7iTk0aXOwhUdQuwXFEKlJJPrPu3veo+nLv8+oai
uuqxZ1iLxNGvNpdQ8bLg/7q04p6M7vWriSlA8NrAC/B10gt7LVbAq7miOPI8smT0bt8DjgscJGFe
ucpdQRJYsx1euPnVEEZfQrgJcmvrNdgZ13gPGTGw2x+Jw3rXPb25yQIMPANl4TnDpcT4TNzDDrZ1
N7iK5nE74Gs0aU23aZO+vkAGkcFeyPJcZeAAUJbNgDpEBHQHX2I3gylZGySdnP7WEiQGXK7j5hd1
nJj4q1ROnG3+SAi883vBipu54wdlIiQA2KLp5lODckMxABC3CqKwCIrAo29bpijl75mvbXjlExhT
AhMQaDNjmMwdVGfALnns9P/DUAcbay1MeWlXH9QAm9R48YHN96kji6aPHsQUDCaDON8F8zvU5C8H
brO0b/7MkkC6VNompCDa8qRK+aDJdtX/uZp2FQRTUWAuvb6TkaiuRBB693iQ8IqhsgtfcXhVMt+F
adIIYkFFSYmF8Y3ygSX+Dz4mvSEqEQ7FADPndUk8r1YurITqf0PupBiZQyf7gZmuZ/iLi2RlQQ0U
msWa6IF+uTZe98Qiailz/FVI09fqYoIZcp+egAvai0lPFnBctwf03uQI2/W1ZDtY2VwKldOFhhJJ
N66ET8QFvvj7yjDyThv2bgFvA/mRHFZh8GA0/+lBB5o3Y8gU0PBheCqwk8aZif5ym+jdKJN1o20M
dhPc31xqJfzwyJrJsw5rB9O3D4mTvJg/DsYSAtlK6e6nLYucOfVYxF0jrccgGgXkyZjSQT+n+S/I
4tHoQnp2agvjiahlboghAZ1RIjoJo3KhCNJr7EtMZZs8TM0E7lTt7rPat9IOt1WrHWf4MDhFLhY2
8DJ9Rq+znGJDdPr9tYngNYnpWAOdVp19No5mrQcJKcFy9au2B2uSxlNgsm8jvF3E92MROhoAh2xk
9Rbe+lieXC8J4pZ8+tuTpsZeDcgr/6r0AlDittD2To9cyiDaDiho1Rz5L5yR9uEdT+NnXd+OHZ8R
KZP3Bu4e+0avkJ47+R4tGlanQAMN0kQR4IXcitLexEwnbTB9p8uBUUAGpdhecPKpSqzKGSPlH6Qu
hCl1ZiuEXnXjgU2TSrTQkKV80PDn72qU9UEws/if7+RDaP4wgpABLFmJhXJBJKqE6Fyfydt249qx
ML+RwW0cEJK+UpY1hkmZZT/q1kOnXYNA7Kv1iCDiflI6rbIabjwegP8DZQB7wINZoTkhaULDc2/Z
8jlbJHsZMAFrAFz4zug99FQgccq3WGhcHxB4AceK9XFyag1Kx0OUFGQ6i3+dt81S9eigqw2o8kew
6lcRdykpXsbhI1RLtypkpF9BVW4K/LmM7r2tLUGgB3PPVEUFlkOlVJI9uijrBcNGhlDlgCEU7EPR
Zz2y8qHFpk3Ge5KvJgVa2APUivQ2VAddQVuklY6PxCCjT+DKOH+bzNvW1XybHbQQOUbEXAoL5FQ+
/8g3iPEfaHSmOnyKFG3ANMah1hgBxqolOtlfTGm1Lslg1tqTq/Soc7JwfwCF5eaDqZm/DK6Tsci6
saEO8EdVcxVs0f137IxxTkgEOsJksSJF3jfw53n4Y9TgUjTk0x4m6gF/eRJ0ZA4LX6cbz2rprx70
II888cBTSEaeEFD/7lL7KeOQ6EcQPf4J+yjacOLNlJm2CNLBXbcNNpgw/yLBqD3+t7SIVxgL3J/p
H9yDSM6WirxVzcU2JFBE7/pQECjsuXiCWHPZC8SpgACR8+UNqaJAjbg4kbMD/vWMYPJAVnbzPfIu
ZOzkWQAz5j0CtZ82MtGtk9g+meoD4hmUwRevuaniUU5mmIRwcFVKkXT7zttiFbLdUArmKzqcd56e
eJ5i+uNKjy5bbRAKzqK66nhxaWu2p/iSHzngvjct7vWRLlGXxYxyE5qjXd8vrQXgKqH+istyjSkx
PC0WKlkZ8UomZnJcpgob9Hf1kDKseiPi6mYWq0jJCXSow/+FRdDJA6P9BBR7s2YICQ0iuk5lJC6c
hGmiL7iKkwkW/xHQQemonPAI1x2xJzsm+G8SrZ4njVF+toKzN4Wfoqwa6IweWlt0epWF5wNPP9pr
aaVDm9k647wOZdfTUQ90w2kpLsX262VD7eLDHhXrlZc+O0V32ua8q1kJk/R1aCEMe7U1razGfyeV
Bvl1Y0HhQGPnmChooCrD8zrJrsa5SuqP1HTV63YvAAWAwpoQbHuo7cqJzCujud4VsGYMNWJwBCZm
stqtxZLs+NM552dmJ9jvT2LBISmF/MRyykUtBF2mMjAOfJFfPyPRGsr0RN7DD0KsRS21b3ffwu5J
2wSPwOpT3xmrgR7KbP2jLz3iXxoLm6IMDPra0J62mWq/Jpzd0ytAUw/URt9/Kug8mfk+MgEEQvUe
/l64flGrrlAYkcitOk6lk9AkI/ZoYUBW5BtP8ep3zaVOeRdm5A7ZYymtetGCMvXb3O/y2FoxH/+j
w4xi9kEuAi+nw8T7g/+F+oI3u1ERlvmtLG5al2up5cqO3aOqSQHKeXXXs3RCKoMVYVnH6+Fs0qdd
jsFB9yai9MdnLndNlxsemiBbbxv48cHhoDj6ZSnOs6U3ocjiLIPRxkd7fmKh0LTOfkA+9fPlF51y
BXiKrP1oj1F/AG/ed4u3sSvW62RFj6QH3W5DVgTSw477AkSETnGVAcdDJZ1Un6rI9a9G8/xWAXPu
RKzyLRK+jqUYNDVcDVzWjf9yb+UP18ZUNn7OeMvvutmWxyfGxTUnyuFJU0afjj7zpsQcQupORyvv
U2fN0NO23ACGYVwKwzsU78pNJCBHI8ef48f7nyBOQe0rNy4QFUshzky1LhT7qLUXxfba3EuX5cWv
6lQy2KakD6ht//nH+Nbd0ii0MqxKzmFQP3wZQb8T7eu3LImQi88SW29PmVenLYhTVQxaudEWILDY
mZsN9IeUewznE0DgG+AAgo9GdSUGbE7q4rD2u1WDhyyU+GHJ9YxiCDURRIZkoc5hHL8RzM786wNc
K9fsnVgTAcsIPs0VSV+dK5LcH631zACIr3gEfga58v8vwd5ghnlwZN9S1/G+VYPYCt5/iIbB+TqK
zWtb5pVzFfwYKMEe+WBLzx5lkdfcHou0l47DardtE7fHUVJFVpoZS99Pnu0O+0w5uBJt2N2Jkb7+
UPpr3U86uZzSW0ZR5Ol2ducA5/qhYb/TKRDc/b4mkD27CXeNqcoUvXqM7rV7yD0rQ/mebVYXU579
I+d7SvhN8Xx5DXAaTDg2ymFwCpjaW5mPqCVWjIwh6nEYMr0iZT3Vf5NZh/V/gTDbOguaHNe77EQO
fqCZe8AZkYSRfqi/9awoFKifY86X/DRW+ba2NYbsclgUoH3vU46j5SixDzCt7zmEqtF5GUJtGEZa
RMK4UKht/Cm2jfozknodz1dV5Ztwm8y8VOH1uP4r1UCJj91DT1qgsKbAhal1Y7pI9wZTRfQxN7Cl
38liSztxUG1YdmBvQ/nAuVvvSuKYdgEx+yAEKC9sM0XtIK3Wnd2fDjBFba/6+5RA7uQn8jrybBo/
4upqDuelPOw7aVqofYwKIZXA6JE3ypYMrFLDfyM0f7FNeVfFUURiJVR+fL0tchI0vQM3bB4bxeNI
0r9AzgUQjCggXCDhqqRzDx9qIb29EBCWUMgyaVB3WeVc2hzmy/VEHoSEXp69Z1jK/sqRs1VGGw4y
DPNErLzz996iN4V4lKesp2u8OeyonLxBTtTURmDUKGRiJB7462EXCj3sizSMwFlQtmFemz/q/+2l
7Fr1j7A5NILtfkvkGLFODdBJGO3LoB0l0waf3fpTEqElMNvT9OACF4CqXhlSqFjsA7RqRFKNrKSR
g1xZEv7WzDfs/q2RliSTO58Kh9pAdP7fgAGwFiREleVk5SGqMevdxRhIg/VuOqPDXEbcRxteQrmy
4ASgXCouSYHpRECjLvfwRuAqG13pQvEKIE3mJ/4N1A2tkryKIV38iON2iMzNbtReJFwnJBPntvWi
rsjNDED+pYFXKPSLXJ9pKzSnuiP/EWYmWnXrol1qDxi869NH2nUDHeEc12fTOzxKNHW8TaoOqwN6
uM/oQ4vXPxCSkupwcjgfK8ndwdRl7sQRYFLn0hX+FKtXFtzW5JZa6i9xcc27Qtjc8Qp0di61f/eg
WGc1wkaJhzTHu00ri+c2+KsNMWCSpiZcwa9ky/amO+kSvZIoGRLIOZl5YyehSoIrDDLZ9uQKKB8A
+nuOIWEKSE1FZRnmSMSHXmmkPZEud/btKMK5gxV/7NkJe9zWQs6Aztdc7th45zkNuO1qUASQ6T7J
+BexHDnug8sJX4264REDtGVyYIyDHH/nKodlxBhfdsFHBPfUKWcO3UR+NGNw3ig6oABQtysahyPS
ZdiUXXfZH6y/iz/KtYGdzS5Ydpuuf5ZvywLYkae9RXaXaaOvmQDAjdfto0wKWQzB7JaehyurY12p
2tu2R33FWkQ+nDLNHjm9k/rFutDG58LaQzSFCfmKUpbh+cpbibP2gAjPINiUOHD16f+xTvO/PdCn
Yy9wkV0+lQyz2UL3I4UFJ3MACEPFc0ycTywxkNlkwdhqbZABXQ1nwwBARQu/4Dl/JzWSGLVjbFad
OI5Ot+tVTvjdJuHvbh0SOKB5fDo5DsmcmJ4Rb5DZwiYQ3kfRSEf0zf51FZQNc/EE++nqDMvEohQu
Sr56XdicQ8U7MEgakYGaADbdSEtQ6PIfqHKCidWIuz1z4tPB0Rx8WPtUsN2jSMcX/TskHLW/X6jq
idkBwndxiqT2t4G8Cdka1dqbZHwbzpaEF/yzbvQKzyR3MltnSxqF/auf34ehkMGV/x7LsV+dvazz
mZhBnzt8hdIOYwOdGEdsfTnTXYbiiPX1heJPe5uwl9lUKrne9mKRdHUyKZsg0bc86+rshSuaoAZv
7WYmWYNFmoNAq2Kl35xq4An10OpLHE/3LOXCBZYLsP8UWtnv+JOasSCGaF3C3lT8e1D+X14CoeAF
PwnG3pkySnWPxOrN6MqSFlveqK+RQxUVQBP61rOYVVgCHQT4cxVyEmBhDjhaS/m8wnMolT5ZOGro
cmoKLjfsggM1AOFJ3/RhOc1aL/hB3SUGeWGGR8wns542pg3GJuYi0ZkE/lUYEg2iOrfS2jzRU8Hr
WYi6vHeGaDCroFxjOCxgTW64EKK7j9FuHMk21Fh2/v7VC/7d9VF2rPd/fPEodPsWOg7RJc3ynFJH
MgCpnkddxotMnjcosXK4QCMCeaoHCrzHQ4ZAULoDhW9gVMoHrk2zA9c7ODqnVlA52sYbMZChaT4v
nhVnNSAB0wJK//DMtVZdDkr1ShH/eM2YzVz9ZGXl5aQ+xtctyH4fTvPgbLpvrQBYbptXB8GLH4Wr
gecUFkBZXRLx3z5dUIQq9dswySAto1teU4ytl422MD9iTOSvDu2NVep+/dhp4LeDj2ZrXPsOs4ka
jjA3yXxON6oEHyYaFM0M2LDHiPJXypcgtRJf3E+Wt3oPBez5rc/RjQMS2GTPVug4X1JaoKtjkiL9
KYzFjjn6FXx77htK6bfAF6HcH39LP6jcIRJG+joWp2yzRDUs3rHmexVzWfM6hxYQuDLYlC7VggAY
1nD770LNdYM7Q+VSNqfkKTWeKManptc4mQ2Swhfv0+5ov8fMKE1y/2wWn9APsnc+FHDWapwWo/de
xr9RJjYby6ljkC85vhM33fvoWx6VXqHT7draoceGIUVPYiznG9nz8vRQWf86vcXIJ3JDPi8SQCkY
6PIAPmKylQIvBxf9Su4DnfsvXZp38R3P68HeMv/ZB6KoilW5+kKFQDbLma6o9s3tmmM+YlFn+gt2
6iaL1Q4XNIxR9ho2cmhZ+0jfb6G+mzvuPlAVyDC6900KSwudWmUSiaRl5qDE2CuPC7VRaI2fP47C
3SwTzLQyKcoLaV2lyIOkywwqdpJZ03qlTJC4Bo8KIo3K/PvnFF3v3ncdV0tuBArfc12Btf9EpD/F
/r7V0fwmCa0Xn1W2+USGFt6rgtuEoh5Nk+0Sj3VTzKZ790tLICvdedKYp9UU8pYz2O/tVJClCpA+
xzLQh6Gk5VHxu267KSYM4RzL1R86T9XmesxoBuba+5/4+5dCVdOL0Fs/fy12DI5ZRysf3v7CLZgn
0vyJuhsciRY32gzjt/4QFhU+rEiifL+PbfpBnHdtn0h9nV5ENkWfXXa8s4HGavC/5MgSeAMj2Cuf
82wMYrIErV8SYPPu0iGk/K34j6J9Q93d7Pzr51EDb7P/7eHvCcGMZ7Jc8I0yfZROdhDgXiA/AGoR
uEkiKGGueZfu+tk9/AqLvAJJYaxhkIRjGOtGIAsogmZpaWsPjZlxZjRq13GJn+Sc8Ya/X3dhP6h7
IzQePL3KfRwM60oQQgHK07Qm2H5lA1BFhDOY4iptv/CPvU6uzohh1G19v1IHKM8FEm6CjFZF4qjr
Z5JY9S1rIA0HTBKlAeg2dGXPsKWTbFYm3oGvUDm+5oVpStFY8idPDYRiKe88xxtrdFhAtn2IHPB7
lKoTbAdpLUny3n5TzCGccHOF482M7Py868uu6zuxAQuI36/mTY7j37/Rosr4DdPFEUj6dVnJUGLJ
q1SoajEWqgwwdQAmi9gSCwAfEdNritqzOnNSDa4RBKoAMO8+IhaX3ULL9fPP7IHM78WntFaM63BJ
Q6TT664pz9E3IfMEw4fG8srXXofewzYLwHtbIMLt8io2nnQcpwMoEtDIDiD61phebTm/b+rzo+08
wnrtyNToU+nk3nkiux8NaTaSz+uZZ3ewMdqLNh/L/BM3SLtP9XSfYNooUMEX2WJuXPCd/N1MIFAw
kzopLkx/RK2n48y6QtcCu5KgpqPQ711fq1E1cSnCk29I4mRULsyRzJbnWu+t2oMJ1cOdIJClCwj9
EawqLQg5y6iqzWkr3rT7fcOtX+6Bfp+roQif4oy9blgpNP1F0kAooX55myNDBA2K9UDBGAKILYaA
1meOe2ip2I6pRVW4rd7xfqgCajxs9ImrJLr40AUzI7WxsQBMFz0sgvm4VJnz83ZrTB7gaFQmLUyC
W1MHKpH6mHrOgVhf3j1iMoP55gWQQwuB/gCjh5VZDvBYVpI+TQnvB8tvQ+mLvo4VexZgIKgEkLTG
snde0f43iEeB4NKshP1TqSjaQQs8oUQ/TTQL7wPZky1Ql9Ws5bO0qNXoC6JDnxfShJBvU6uFp8BU
yKPNLb1KCQpn/N2GvPp3VSW0ZBxLiGPOa1wFV7Aek2zo4QzORW//GmDWg2+ciDE7VCrPUILJql01
yieNSFf+MkXxisZDhhIMyRKOBdofJmF3imwqgD3AiooHfbdjLZyZhbUg+/3cqMmvEywBFB4UEyuy
3b+Eft1keEsWdGXulnseUyUBYI8tZeYG43cjAJ49yoHLAo6vDT7kQD/YlhkIQkJqfaYAjPAcosEO
lkblaJf/VnlInQV80BMhwT2pQRTnZ2IFVBBk+JiOakpJVzzc0j/8txDwunHj8EtHk5g9fHRAdFDb
GMfANnVctDWDRCjUKDdnJ28GFAYTXkJZmz0TWK7UmQ+u4w3Yssik+JOzLP1NzHSpGxDzT7OWqkSt
KgQrdmc5odbjXuYlCtGVgLfMj9fqGxNUJmcVCYXDk3AWuf2tqxDESB9BaeAXwMFqXsU61BzciAAs
9AVxd4aqwHPZeZmd6dxkCAuX+CUa3TDCvkgZZvL+UfPQxwuGd2mI/a7MRur6QDOo+jOFFcRrYiMV
AxS2R8cMFoqdvMUfZBZ8DXLPtOKgcLGf/8NU9TYmi6bEAQwfu9emG+QfbgQvmkphLMq3nUXvQ3A4
RuMSJjv9ADXPf6KMmQycTOfeAikG8BV9Lb90O5uHR4GeB+Eyyq50xhq4laNHfKuFXJB/gzix0ROO
rq899Pbv6Ue0TxCzCSzZeIWkEliCGteG5GirBiZH2bYIZGU/zmkQ+KbAnJZgKy0t/y+kJQbU9ZJD
TzUPPHx+wOXtDAogvhWWoOeZfKW1VGxmJHCxXsw68DRTtHzPqjrokYpTaQvIrecY3ubhuatPQlUr
9IV+yR5pJ9IxYIiBM2EautmgMb59YGGiopaLiKYrcY19sWlmADqPwGKXWcKVkedLGNx5QMIH8mA4
B09ChH+viYCoYrXEUU3rBu+bZ6Eh1wsUNAh4yZ3wHjb7efwo3K0M3+MfnhzMN9Jgs0ynilxO2U7t
sB+jHctkdGOieU69e9bEFmkkwy65Q2SWRSWh4qFdB5KfhFAhzU7KQ6zcN+bXX3ag8KnJUpBLH/Pr
WTLDQ5aIiYupvm9VUqul3Xg0tIW65EzzapRg4Q8SsqlDoi3GG/IPpCW+2RSZUd2f7ZWAVcMkevYh
hLInOohPk7+R0rkwhIyzGsFxJTUszGmV4Qg/nWJzxYuviSzLIzcXvk1RBsfj5j2thaUGX4Z4X9Ae
EAUBvIkeeR3RJWtmEmYrp8b1UqsbOO5BwqNZWjxiQqHyJuLdHQNp2kLwCXDwbwMvQNhGEmIUnGKt
5jMUd4SShrA7e0KSJznbKcYR0TQd6pNOZ1E2YQAA3mw3K40SPKJpHDGxGhjpD+EWKSKMii0tnJ61
Ux22RXBckyDW6uexLnT4N37+22e+9QDxMSeNcnQxVM6WP/pV09h4xAaJFxJCMpeEBxTtM68fjb/h
n+/xuAU7xkj3iJrhiWTDey+LcDI0xhwCkWnTNlvZPyuzWzIXbtHL1SfeeauOWKfEn/mOqAHLbxvj
ReXrlY1bxRNMNd0OTZnX88GnqZFTu/V42njuTEztczGzF9XtrndBhOiDvYHkcr/QgT09v2/h7Z8B
coKdEAwEcrTyqC8yeo4LCHq4Rh/M/AAcCfdjbtzIDAibzW5JmKvpoa3v287pvhL5DXUVeIq0DWrT
ZsP3pmGckszs99+XNdHzJHY6B2LAObWjFOKBR2TG+LD/Gt9rntnclsAesmRbYYf/VhWgr/AEHzC/
GIHQsjwG6I0+zh/CMopXOSDoxTN2skFkqEyIB36R4Lk+zIBgR6izZEcosle4DFPmZE0dQ6Ovh1E9
Wr9MIpZzW9Hca4bg6sTMi3lEwUEOx93/ZPYlIv455kowz2OT3dZYVDHkDfmeIvRzs3WW+Tf2td4M
Q3sREMz4V8TJdbxkHZbjVq6n3beMrOPQuTiVpjilGiGCpPhiVvAJvWRQ4pXpgHPDO1enX2mD4y2F
ZvP+adPfPKjvSNB7kKdgiBR+7HG8XpN3hWN5yOyWrMAvnmcRHqmseQyikBYJ9Z8nuqUe1J+wqaGJ
KbQCK1ZlgBH+A6eldasmv1mKDsaZ03zBkt7rNi5fvAFrwI+nIYWUlkF5a7NYAxhxS/uV0dw2TSMi
t6TtDAS9GqeTo1tPJ/wwCEyepHkYGeLQskkikPOkXVpVWH057W76z5tqidD3b/Y7q99LnlgVowGT
cHB1fL8j3Eevf0dm+QxJwqOR9JBURykyUbHtmV3F1gCHHI2K14W4jVcqhSKfdu4xO1vlbuvRmM8x
nZz53WPcZAcq7ilcqac8k0/9H0J4DnSNV+7nEEmZY/ehklVMYW1jvXIIx2+YUYAecHO84Trrhmtm
mwxyOaibWp5tPlydXYKawr1biQJy85+8OtDL5iFSk2GVkFlAIfRs6EL1MDssP1OdOGmNxzSpU1v9
zaoYh/FIAVzKf0IC99ldJt71Z1a6N/zD1LVK7UVXit1Zoo0DpLkzh8lpllaN8zUA0lRqn1wnaW8h
Wp2veEiHqjJuZhsnk2gtFS+Q6VwfuGRVjlRfByKcjJceo0Cb68PvLtwm6ybTsV9GjYsFOmNtU4EM
FaCXOA2BEbvRvL3Y7OSWrfBp/WVFHu4xmSJIQr5WrHvre3tWHbGW+pkVz2rgUL2HUTpJUtY/Fy6L
zoLg3J2tksroKE4qKhGBctVJ4BCKzo4OH1Q2vG8r9LN8gUroW3cAdGWx6pQfN4oNZt10eSWyh4G7
FszTRM8a1FyxeKDdYPGtBybpYwwKWOrILwxlkZPAumkEjLGtAhGyAJCNJ8Q8T54XdUifU+XfoSIG
96isRtb+kcCEVzsR4GEC8qIp0MCTaFi1coDkBoSQNYyuaJ1MyI0sUbOaSx16pdA7M5cljnK1ZMcx
cyNwFnk2YXiC0Aas/m0sT12D3otllXqIr8E1Xs6U6s2RrgfZC4alPpN2fGQzi7o5XAPmWll7y7rW
IBQcMQrbF7xlZyxIel9KA/hPCRoHkvEWrvedtiKdcdXeYDP36gjoYBtEDH/O3mewi5EXnWKA3PQa
5kuM5fHhaFqh18fsAS6TQQjCCYH6o+RBxDRM/ixcUE5jJ2a5g/HX5YHsqIpVPFS8TdtMYbXON1/c
0iIbdaK+hWUVxn2nnWJGZVlhHV09OO6fpRS79LwhMvOWnykXzIpc/n1IysMjZSY2WJFJgTrJdhRb
CPz3+aF0RQjIK7FOESf3CVVIoZl+iwOoC+B2ZDXOx9Hj2BlycPJ/3jev3BzIXMbjawlW/66DzzOt
6FsyoStIY0Kp9DvDaKMQuOP8yXq7Lnfpfy7JayVzKXixtIQKI0j6jEcmW/0+2JtK+KpgFhvwGuAS
l55Pa7hqAZpTbtZ4oj7sec9xr0ioGjt6l+P+pUk40y+zGGhdOKhSpz1Iv1nBCH7p+sAElIChqYyS
gXfYYtw0swa5MsI0UtUPrRhFwUrzb13fJF9ywAPlG69Q0EvFrOEaqp6JTGtDiZNfenpowiSuUXWA
1SJUNtwys+wPILtsh2aEbxSE4cJ80amlt2fT5RokGthW8+HN81nUObs7THaRWOAsATtvVM5x8s2S
UPuDwp7oUjbVGWrmG3pxYTFXQzLm5kNq+gfo7qOmj5XeX2ZAp/HS2PXWvfIgF0QpifALEU5iU1OA
GSiEZ4XiWDGDnqGf4jcf/D9gxox9oB6Gh4v1u6A9WdWaAWPMG3RfO8aeenMhRiI2Zhx86CPILE/4
hvDgsB1XVbeHDwJ930A+dZxsn2hl+fbeH/JZ/2+hNB/5GzZ7nAWCZ+fORxma/+CQDvEk7O+dbE9y
ZafC6RLvseGwPZfQ7hcXM9zK/xStuTgHf1F+pHxkNP01b3Hu/STRS5SYa948FcVNdBA8lUD7xyqN
xUbd+/C+z/85CWv71zIoJrY15XD9A1rnpnD3oGUiZI/7z3CwPTrFDxlw3f9Pl3xBmmzP/XLJQmgQ
0FngfJfFik23p7tz6Y7veaWqClWbePHJjGXnlo0fvn84PZqaoXzaIN8AejLeLjTlrAAg39T109/K
G4DGsqU5taJMWuihpKyRQ8B2FBZlTW1+s4K26tgwMO2pgyxpHqdZN1NC2i0ubh4eAqyn8WjdKcsc
1c0ReFCLzmv9ba1tyGfvCpB57GOlDCmG/7Kk53SW8nSZYBaMMMtXajVAubDuUhyfr0QMAIpmjFTC
mN29+OgWmpNmGjlyTVkGkHX8273aBnCW/PHc9L/dAaWHF5gqRa3ZY/FswJMacBZPnReRUBiaarCG
O2ShpvLR70wf4WOvgaTxgms3Kxak/5hmXhS6pWYK1KjuYTzymM9nTdQ9olGpwU4Pd9j7Yg/vO6cv
v2MiD/hsQlcUO8AIBAeNL/y4W5qa2VEs7caegUMFtiyQYHSKE+qE6tT3KGlkCIoPvVkdDxSAe2u1
nmmA8H3USwIo0BZicVq7qbzfoe4dwPGfuiDFH0MsWmZcKoYNP/O0UGS6ASu/WfD72gTMfrT9qPE6
Akhu8jJ4oo57nu/g2SEJkd2d5Cq1w6cEXO83flleiW+e6mbC866YEJEVIGbYeW/J55mtFr5e8OVX
bD0HElqoYQfnx0P+MZAfD3PVrg8rnghX5zFNeIx7nRkPltRaDwT3oaDJEge5gwu2/AqcIcDPWLpd
8JyyOLUQNGC4DFtWSbpWYq8pNIBN0jXPYAzmX0tTJMBI8W7A2Gpzb3ON6CvIZFD9F6KXAlbj1J06
ISeTLMfIuuvTIeS5iJJ4M4wsK0bcGStEB8Jvu2lbBe0XQdFtHsGlyecBeZ8sf7+5ebnUcDvtZLCA
IV6abxZquxwoz+hGDuxFceTmzL+x/BBZkQD8xyZNc7Hq11b0YnTMNuG9g4ZpHMLwQhD4Gv6d60qj
xLdKMgWxegOuOXxAltl6Kmnck8bRl0voIWiimLMZqkqKM2QjdoO1gMmNr0dJtEgnbD3ZInMN1uvo
ElKyV0XuVXQ5tl3tF9vyaGfupDNTkLSgCC/sVxTby36JXM/jdzloby9SYwl0aNf5fdlXUHLhqYh/
wue+dd8rewBxLjDzWZ/rjCALYlc2e4f6Q4uJWwuyrtoSBhUojB+FLdBgrBFEQKFLqzycovKCKxuL
ipVaai21AwVqbyYeHn+zxCbEFHBYm4ucEJjpctPiKX+O0kT/ckwilVVedUQe6EULFsUjb4N3zY8/
XGjvq6Otg5gvHX9mD/iOmnGChychTCsBmm1dasu7FL7Tn8Ahx0ZZ50bM4g8xLcqB3qkVxfyy8vl5
K8Jy+79uh0JcThStSQb0QGRhLWcEHCW9rt3mWKImuShua+gnt2T8RnuAk/g7mSjUQZuvxkHs6n7O
AiYHFe4m1fdPhaUrDwNXLAUH3PMwPKmfmpOKyMEZ9Q94xmuA8NJhb4Vp6GqoLLHI+ev2BxU7Hz+M
iZBhC4scD/K9cRRqSX52hwAdsVLQbWUyWsZVvS0FnIFabZ7kvPiT7A+l9cNTx3alw9Yer/ARPJkc
oSwqI7xcUpv57TRyGbyQnhDZqysy/26/VG9soRNF+ZxkKh7F/w1fe3g6aNa/eMs8LEmSWB/NYHH+
ui/Mh+PRBEK2/d27YioQhKr+7+SRNScgurZSDA4pueOHryNnyrGqiDc+edO7vHISOVnB3o5iIbq8
FJLRrFcCR9rffsU2GiZgEIZrnVTplDbihmCTRy2jtDloJeLlk2mnVegP4LB9EDqQaxU2wEK2B63M
TjOo3oLw8lsmCBPxkwVfou3oFGD44pyRd/khdVlXctyS+rc0B8IdlLD8ehcVPcoT1+eVpGsQRqwp
4+GLk1Nrppn6IYEpHRDKHkcZk5eXp3innTYeiXRr4LxZ0+3j7PwZTUojvqPChXcG9NJ7EigMIAUE
ADeOFRXJG2vS+0Xn3WpSZshYaSWYrZH5A15je7c/H1WXJqHABSnunAP6cd6of68Z3s4RfYdS8TDC
YMEvaUQJBlXwsLki7eH2kPMaBAspG+3XljRViUELgE6gam8+NWddsY8yjIca5EWa4WXcVTHkEEzz
7ciIus32MRJoGXbv0/XvB4b//HQYI56x77Yw1UDJwjNtEb0vy0KRJr7YgOd3UkuNp4B6jWuXx1fb
tqdWuPd1kHOa3L6SFXpojZjtduJ8f147yJkHW+CHwGlqnxjrTLV/09+RbV8mhQb61xdwhzhbLG3J
BRzsaSfQDzZAx2fD9akACnFQkjMBSAtEwy0lqpt1JGF/S1w0iKN2bmlT5VJThbgJ3Fl7JVwJERbc
wfRLFN8vR89WllArfYOdAfkSf8Kn6J91qvtlwbCzg+24NDZQEHB6N/tL8mx19OkMOob6RzHxxEEz
FZ29oiVnnKfdulnEJSJE8Rf38UiVmdYnVHkmQX9zNFvNE1Vpq+T5MAd7rgXGwNeEJdpsSiBHfkvJ
Lc/ONX987bju8PI33gM7EbkxC04ny9NGJAY5GaWXM1zZucmNTzfGdUo446TbbkPw/H8FKV/WvEgA
GHPqcSE+f3rKow6BnYOSQ6Lch5Zzjdd/8ilsUpOL3z5JxrLJGFCfBrHmF7kIb5q8rN1j3AA7NdKc
SWwKFc1CpVFpq7IF/6q+g5oTUbxr7GQKcX7LYXHj8MZAspAcLthyP/1CjqgWzDj4psX2NFlQijjW
c7cA8YVGO+XR5uWygI3ceeCJXrzvvMzXb6oClArZPwI0xYTxA6tVbeTkX6dkdEnPoEkNI+0/vguN
Rpw2SxOv0lxkdudSA/fyaa3kwmjZPNQUZJhX9aBFFhkeH7HhoKj+R+7FiBXxPFPkbbaVKmv0R5MF
pFnaVaGcOPtsjLKVJ5lI4uzB8ItDIdJcyKmzzGEHwvVw/73A5a1xWB7vjqxvw0plnHePWY2oiNCz
gIxCJNpWU/Souo39jqV8ltAonLU+9z/PsR+tF1SZStPCAezwvYWUvrZE12hIFRcj1nSol25rzcQc
WRjitFKJUFVHMkzjYoAZHfhxloPnCT+ZXezJ8rE3JLh6IGdlql+pfrG9mwx5EsH2daq6pQVSJNqu
eA8CH+TqgsbfRaq2tMu0Q7gq9MPmJa0Kr48U2V/jcWQyVHLRnrRta4PmDdAbC2b/Lkp2b9fbUyqq
XcONLx9bA0VvMukoXLBipbiYU6B1jTfuE0hr9Wjfwe1ZaWNxal0AQfX7998yJkVqEYhOJTSK0xgM
wUM1uzdJJXYiUlRDAPqBO7lbPnt7KR++DX8faIjXw4S0OthZnYaUsGzz/e74oB37XoTcvahSTXIa
FqHoHokVyvxNXF9gIvJLVQ8fYw6qqdtJwJN6Qomh123n2V9jz7xOOl378un6dQk31WkF6WhzT/9z
9rsjHNbCxRWixRoK7VcOJlL7JxqE6AWyAEL14zmYVARyi2HRfSscmH9ULdgRFTNEF3/FB6O8mL9x
m3lqZAvH5UTEkcOe5oUpM04rNQ3WdaiMRqqpnSC5nxM2B3nO33OeWMNWbOXyqio5GIJTmQ0CqUMW
cNWU7JCeLQMBKXL0KVRi3kI4EEvqzOkjm6E0kGgLqPlwnXQe0hh/Ek+RUOtrM9cPqzP4sO5IqrKY
4krwd/TOMJMKUBco/6TKhDbu4DyGqcyjeJDVu+ZKArRA4HtgaRHw0nv/YOULzgICc7wOH8crpP6R
6+w3NAQvpDaDaZubiq2hg6ynep6Ge1NqjdUN/hZbdTCM1IYYvXnTGRZd58DDqsvuNz+2yTuPOqJE
VD8GOfVciAn9W1A7hTXVQ5XRitZ+daq0kBJzTSexkyPiVADwHtbSaISY+ORLszsJVb7ce0dhdq9G
GYYXIMNNAFE6bOistSG0inT2J1mAMI67W8NA8Q8irPMbj+VhhQg1Wr4dUdLUu50mWcKJCNG+IovE
1vSw7E4h13/UySKCtfG0/j9EK2ewL1zJfQsyiSLBonNy71H5XQlkDb7bg/5JDODX5am9djHEKDPj
ZMHRLBOmefKgZf5XR43PdIJoxeIZqjuy3D9VMVZrfFsh4yVF1RqRY5dJferNFVAi8uLQ5UXssfIW
DHdVzfJtmA3Wu5wIjLZhQg/0Pc+kix/MDATxtzSN2W96qNO61RPQHZ8be3TB3ZLFGuoI9YCQ6/9p
eXnQi71z7e/77I8nz3jpgcjv8RBe/bMzIrrWc/S9fFaC7jw+PMYLfKjhXmmtOtcJMLgIn6wfUWJb
CvqYE0xq+FkPvd9mlBOBjl9LV3leeJmiQOWcy+rfhZxhRX9lLnWA5Ng0esbkWAlfvkGlzRkB6kGZ
hk2EUk/xlEXnWIpNk6Ep0SFTtbOPnAxsrbQmmS/hjAW0N48OnKDTJG6QxqRk1aSLdAgz5WzqcM2E
VwxrOTe8ViTwh8RuF35Xw1Ehu64m3NiKJKl8bQZF1misnwp7RTUDbSCRIvdKLO7KIxhebjmafgPU
gIo1pICRQ+tt9BDiBbJ+sViFqSKrAUmueMXhPlTF7K1kd65N4KJ2Dcx5VuvTtckuIVyW/QzKijun
EEOLVt76NYbcgKJ+MWCJnIuol+FPBguFDhPKKSXvcjYpUbPmMNvKso5TvBu0yLoKmD31zTdR4GtU
J6XpxvSpoiwxJ0SVDKhVUrVWXQ2mmiIK6asNobhkGlAOQMpB8D6AHcRdloISDixhMXkLoc0C9qbz
Ij/nPrnzx4z50BH6OzvPAuQ/Ri9z39FT3XpYMh6fHKA1N5AknOgb93dBYG1woaYXlv8s+D0uSJtP
ln5yinto0724GzZpIkroC1muPXtCqiioENn7ATQnaJSuokRNeiHulqR8Jt/W+RLWGBAn8pVcehjO
NoOlfgRMA3dh1VQ3rbNcssDZjwg8M23IIg8IYbveXnok49Ulc1A/QgMELZR8dFFhZRNuJSkPjZGX
7j85cRz0LmwxpiVJC8efOpazeHD+e6uI2K1lWHWlQPShTbnXS8GLRppjVHFidPRqTjgGxhtCovaC
nzja3t+Tgnqg3AVIIeVY1YpcU9bsU+sAMG3ACONIA65hPnXZiBSwSveTzyjdB9itMJhpOObbfsvA
F5Xlu+44vEUNY4s6odxS4X/uqEQUvMtrD4u+w37N47WShPNvQ6H/rOGqPROT7t5QIrb5mGSTQeCA
LjQiVVjJhP8bl85oM7lroElqiShTn7ztTKnl4DDlNpcnCsmYfyjZsJcjSb2X7OYMZ4ncJv0f7Zws
bzW60VZEbqRtwFDlo7xb+FT7uENnAaCuiy5XJKqYyuz/njt8pLWQ/DP/JZkF85PTSOkyHTtp/Dib
4Ln3UH87/JSZZ20Rns6okvR2eIVQJPpD8xuTxjXYXnQKEj6SzrTt7jCRZR2UjHRuLuF01KwXv756
lu3QrL/eqSgApNAUr8v5CTXTNa61ODie6yC+SwHwWUR/RRQ5DuMqH2etrMigHSYConqoqDeU/7VQ
bi3eyGRDs0AHMm9zpIDhuKbeEIP+Vdc44iiAhrEE1XCf4afsDD4uehhvu48CxFq7QT+xH8Fvdj22
y69sYEOpCOmD0b5fpOP84N7lz6bt/x0kf2DqZDjkQrNZdsc9sy7uvApyyVEc376ncjQUCT/pO8eJ
Q7HKrxlEBJnUYOxDEd0rhEqEAWRkDv3piFTD3jiJSMMrAR8GQkB1YtGjs+twqClK9ukWIKpcJWME
f57ZmO/F2j/j7YLhkNirAixTmD24VN/wVwfiZdXjzyEDGhiwoQ1o9V0pEBuq7FMlbLizFJ1eyo6J
fhZNKpepjXNbXAcoaRCg04XJjxYZb9ZM92WxG5te39iCJF3T1Z5I9amI7FYIwW416dMgNe4C4m8g
oTCPCepXu5r7LqWbYpGRk2ndJhdhl759O2T3qxn2GshkzjAjqyuLfizlhBPR2KFXYNdRyehcA2Zn
54HexI5T5TZZukntUwORPanANq1iT/wR+COziOpf6ovSouq4n3DFQ1jr7BADHrB0utzR9nGU9djP
vXbN5P2KBlheEseK7TCU8dl76iUeyt5jtoROM5E9H8qONKSZk+e4R4xWF55vjRTViKxF7pD3qnEx
ljvP5HODUgTGZECJ4MNq/VLxAG+ULGc4HKjlygI+OxcrCwl4bgPHXi3GM32ewDH/FwGyJOcjsVIk
rPBWEU6GQcHgcNLCVYa3l3VnAwF+ychJJf2hNl4iNK6eeZcihJ9oe40cNsODiKokLFmJsiMnW9r2
GVAx7Yu/zrsMiTtBO0INp/x6p7MlhY3s/megpzDDrmaEwsRwR2Am8uzg2zzuQyewdnFJlyZjs4wc
mGyoFwhmEp7PypC0HqhsyWKWIykgWAddvPK6AU552GeV9l89ZweQyK0Jn25dWco1NT8n+EO3r33v
lt2i5BpPFAIpjyQVAldHYW3D/5G1jNr4xaTvEIx1FFZQClNAX3WQtlnVfTzxeawk/qR9t0E2Q1lT
GXuqvzeIRFUrLz8g1dQedL4ZRmUnfmISnxkeQtK0PhXTypGws2Dr8EpSH4XD/pE5WOpg5IoSQimE
Q2c6x7kxfy/VjrsgEQRPW91INN/KDO9gi20zdAFOEhdtoRqumR/0bll5b+4sn7+Hm7u0EWxznEgf
zIE9H/jHlqp7pB8ez26o+ImXL9JsLm7Zah5dRX9u5yeEBPByf++oBIUGVl6sIQ/Y8LGLb/EDd5oO
Irz0QSXQFV5WKlRXp5/QxU0kibywvY8dfe6Gg10XpC+3FiXWsdrqtmWhfNvlENhKG8EtK370+Dmw
XDuz9fZVPBgHI596PLfXEgzBIrdNOGuHK+rqfk5gL1g6QkHbMvhbY7Ycx0Di5ibAYMcXX1t3Eruv
CIAMzNlvFjuB+fgPkoE9ih4UVLluMqUrV/0tokcDJt31sqbVPIdi54StBUofkvBpZysje1KGW/8Z
qXAXXXF2cNQwf8g+MTzcKx+/Dp1udUpuAieOUQbmXARKiuwOkKCdAdo0nPaHgvnNf24a0W1sZ9no
+5VHZM2wBSxrILDn/1FmDl8ge86YK7AZktwKjbpSypHD0PTBZN5CXLcZnGv9X+dV+960xzXaGaAz
UMbm4eSWC+rpLhKfn4QwS4/EVnSVgy64sHnRx7QZn9/Vs3NO7TVd1Jw9Qv6z63Me0C59TvJNtPgz
TUwaEkLom422Pcesiae0ZStzkGQthpbzbOjzl22GQE3WWt/UNHO7Cni6Q3lD9mWBuqR7WQSQj8ek
L7s6qcFlVFpntUbepMNRC3keM6d/RS10UJFDBx3fCyl3za4MCfkIfwIMkVtuBZpE7q4hp+/eBvYO
ZQRXv4e4OHPbyRtce9KC2xVXqr6TgAqEN0wLgHnWWsSwK6nxkH6hBmYZYS+OkqIWPYlcn2jTNHM+
ifnMyF180d5cEyK+1RF4XY5yHCu8PoXKk2GzWMS677EDnMv7XGvYqPEqn7lCCO5gaAHyqoI1pfoH
WkNwok1IDs7vJCMDV07bqJJG2Liyl5WKN+tnLo+SiGMMTUiOhQzS1WWr39tBKZ0TxK9IOMrhGpC3
nwGAcbrdZEJxBhKQA+L6zLMrtKjz+peI8xnE4m+bKCz0WQYNcrsj7+LMcn1CDMZsT/1ENAb7psO7
N4CsXrWW88oZWnuFMMB000sALntPWvJhiYTC0l81twOvFC+ml0ZtkBNrgCCsjeymkXZFcoZ5DbDW
uGS9j8raPVKxkhDn2TbLRaWLl2Sp5uSaBBYWa79w+hlzJzEuuSjpPD3IuLQ415jYz2TuNFn2FCC2
PZPcxe530AIjSCmfrgL0H2Wuj1UjL+s1V7PL6+UmHt02rbiPaweajcS8PRlBju2qewCbZsGELoiB
8peHW0xA0C2hDVemShKEN5D8kjYTZP3kMWMFQRPlxiZxkEp/KvvvxYPtsT9TlcuWC5oOW27uu//r
sTcqRvI8o+EzG7lpwsmPAVangBPvZ7MzdNb4k5Ain/7MQhsxjQMs+cwB0wjaV31fEBMBWa1Bv6yQ
gMsdUqh9nG1nxOjt20PBFhjnrBj/7B2YteO58CPj57Jc2KHJ7aQXFLtBv5kL8Quu0yOIXWgHFqHi
wWfidVu9i5y2urDe+7ezf5wuxcxUdbBISBs1JBwPIy8KBrSezjNangYQxM5FU95/S3ck3YLAFJfE
7sH18zRmrBjpGCuCJ2cmfQAtlP0ompd2VkqYcEhmyLVN8qU823T4P4xvNoNQNqV/VMS7Ku6VmuOs
shn1dAGss0v123ZQppcxFArtm+509COKkvWjssVl1vEnVSJ5AEvGiCM5+4GevTfcnbIXe/RXJz0P
NmQwAKY0ys4oH/7CaEkPA9uXKVGa8kWh3oRAN4Zk7ih/fiSwQmPE8VCD5grtug+aEurpE6ma8cCV
v+TNFxl23tA7LqGYkRaTM7SOq0ccDo29EGAt99GyfqymuW54vqX8mDQQrzXIT7F6/T1nOFQhQNxS
wdIpKkhVyfEE6IJ3Xo+SRCOdlQkD273kymZmhPqrxUkAMALwq5563iEFYqXfMEmmizyM3J4FnapJ
OXS+M914V1Dkv2TmkkDtWdly/qE02kaKDv5eB8eLMv/3xVN6XuktjfllzPEiYxHQTcgx3mlvQL2D
1F1ztbv1l3nbbbhzLwxpc1GEEJjRjLralASN6X3LTA8Do4RE1sg6qKapVyresru2L8si3S033109
4e7cm7J7XWP8vPR9skUjMqGNMeSsa7DqwEYQ5ch0EbeiwA97T7KH5plmWDt0OOYJFg/3qjNCvkvz
aPNwjcnfdy6o+pR+Lf79tIeR5Jp71PFtniHRhlgYmdukXqM5fZclPL8Vor4CjDuKszyjC+Fk9Rj6
ndgReq5UGn2EAfc/4vc10YumjFA6IeIh0AYAlikzrluwbY3UUnHuN1p81qTXpVn1wwf2RMXhpkH0
DUl5ODtr8iEjZ7352ZPfxjgcYdyANuogoB5mHjm/gX+VIDiOrfM/C/knu7uCn2+Gi0gq4SjAOnuC
ThHGT4w/BQIEhYQPnxi0AHhvCpDpuNQGLXR6aJ8M/3Yc/8katCP5F2Tjq0IuPX3WUqPu1hqsKSQB
j7O9HqAcrXGdglSAbMGtHuWaNSvcW4tVNJhsAkP1a+q/3Xauef8AnBdvsaznS68PaPlOBazlBGyu
Fm/N24Pk2zPQ830nkcVT/1KY+Dq6LSds8NUa0lOfljr9VNCjyvVPfqbyOiUBC2Uqd6KQyfZpnV2U
brGiKtQrAQQZT+b0y8G7kYBsKBgb4A3iqGL6Drx/SpCO3oo4O867sIj5ZZPZIWzhkB7gt6/FyZwO
BGpls2Igyf5FxuAmhwWTsIDxjEffTzHpODyqtV70VjIcREX2k0+9h36LET71408eJxfKf/3vWJ9f
J1pgL+aC7MMbj+LNayBemdZj25+wjui3G/wZFSAv75F/ZLnGxZrRGhn10FsVAXY6F91Y7YusU2XO
2SG76EO+VGoDzpJMvZydVkUXnz4b2VXUVvsHdpGSJcfsCy8inY4ZfzuWIQVAQxNtURh8iaJSBOqM
flNfYvJ7hr19RzIQeHcdpYBY3zLd+sLlQSuLUPcXrwTsYN8J+sbEcZR7UdA2u5vUR/FxTrv8Qn+3
dEzbzyhxgHTMFWk4G/Y0+qjMQLLv2jyz5JPlGtzCTrFQ8EzDr9ARxSdHZjEJX4RX2Jlx2ZjwFiz3
igGMf7exhnpEwqX3GMTLObw/U9jhqlIpwf519xH/ACh85Yngj2JSYbE1bhbLf6g8qvUBBL3HmCzM
hf8jjRtvB2HkF/k5y97OmKKCQp+wM9k32y7GsYpPtO5fG90jyOJKr0t1fCC8M3rpQZUBwbV/B6EY
w4FDTDEooSaE0KTXjp3SSoJ7E5819pkc9Zv1D/jN25cpfyfjZWWzejAB13RYJ2hV0+ReoCA4RhFk
x9lM9ZmQElCTtTQp9gIG0OQU99ATnQi7UzYbW27qVNIY9MVV12e2DvsKhBxvenH29rrmEdizruGX
tEayU/Mflyv+GDO1GKmUbA3qqHwEdHDWHhIy7go4VBKxHUS+jKAlvsDpLJ9pWdwQ9iZNI1GN8x1a
qJTUK5Q0Amdy6GIwBSPatmRo8mljk86/75+BpBruLrd6kNltaoj/7FOPsiYvB1FguWQg7EW+2KMH
FKlsdfXcIBSZViFabqdqIcsvArtX7Gw9BpGbTRLJKmRnxs7iUE18qbtalqiZGuTag+6xUubRNome
AOGWIaAmOn5bdqIT1QSYFJN7nduqhH3hmLl4n1N4uQXoPwAN4DwjAknZd6nNk1qbbuBdMp+MliXK
v5yNlNQ4NjvBckcDwMkpiA4K2NbHmkTzpP/dHcqz/AR6Y3cPmd0gxgjEYJxrQs8LTifdIpaGhA4v
KCJ8SQB3SzOXdsqAeH4Blg87luSPsrncfZlgEmS07xwvdjC/9JqYnftUMvWvzebX52q71+Wmd6tS
dh8T7laaQcXMZFg9oBL8fwSYHcMJyqvykkBoiwmHiHzSKqbbUp3RKYSoEHGJvkZ9nCv8vXts21Xy
TfanF9zkBULwHIG9p6QKneb4mQj44VVIiWqaNUWvTKINvva3em/JnHcz5QBiGy14pUFwBIF1Dxmy
tXUhZ9e7DjnSoY2BoD/f61glsk6831lDibB4+wB5Brmfecq/O/K4Q30BPrfATkV8XxCFZ012s9Hp
d0T1XKKZx3v2OZp3YA0gaH0bY79drcfRTRTLyZKK4D1c82v5B+WxnntFf9NCbnp8a2uAe4xS+5GQ
MmmlSXJlVat7xTSXbnEcgZOS4PM1NZM8INmtA9b2uw//D5PfgseuO4K6bIEA85w2GjCbfxdJS+hU
8bkP9ue5y9mXoBWc45Of7Y9CDErgnGzoKhrO+Vk5UzCCm7daxv8D43TWSoJHsiL+xSoQsBSkij3P
O5TDniBZxplV+vYh4nWn3Cd1piDYxBrnMPPXUzQ+9B6h4lxSsPPk2qPO4JwjmGK8QBhhs3tQ1yCp
CBD6IqSKIiom6q/uebpbK9PBNJd0rGFFShAWAx8rBV2ThNRLtwo63L5LQJHe1r0veIb+Om2oLdLd
Ut4y7hox4DiwIsUg1Ypr/dH+xt0sQvkJiksVrg0INpvlITPUo/atxbHY++M0jB3lShumAyYURrTq
Ett8GmmZ5zzlXqE0ReS4AfIQuvSY9aEx+U/ZTqeS9GEx6YYqQQk4LA0C9OmfaDlYFZLuUt4mGsgN
k6qENcAhz8ax1afSVLLBdUT8M7x8d/h7VLCNtXCNfkkfd9IUxg3Xwnl3CFcXWAcnOCDkavvGHKc7
AB8LCua98mU0aGG7fau/DusN0sFqe0fYueVHk1qlNIcmMT+u3IeqYO9hF2pUukk9T9lmGO/m/5pj
TPWEbkVuS4lCEgD/ZbdyBHrv/ksYyE7qWZrK7fX/y5mp8JkPECHcVvZzP8ewy4xYNu1cgrQSo/Sz
ZFiMczp0aUEyWU9g2m5C0bZzTjVzDWO4YvfCRfcXODoakbyz6tLjszJetY9ONJpWEonEK209ivYt
5ncaIUGaWWHakydInzM4uQseiFZ6wBcvqmzD4MimiDgGnvdB2bz6cfVeR2YVlBzKCIx4zXFEb3cV
SOcrZsQnJ1SbBTt/DwHuOAk7V5nYmcHkNutaBEVkKcX1644QzLP57GfIRUBdIjnW/J7eYVVb/M+X
y6l+WWuIMAQ9zs8ea/F4WQY0Zkly4rAoa3fPmhBnqCo/DgrhlBaUXELDWHtPEUUE9cdkaZHbYUji
Ooqwe61NuKQL0qDPkq3HvRBDAWUcEBJeCfYUrHyBhp2FH1ldsVvuzk6HYlcBRTosYrbWIIlavQMb
apxaasTo9sMAnP1/JqMYf6+Lt7eRC16zQSpnSVgHtmUQMZmvjkfRDP9ThX2xwTZ9FEacp9UiybBd
iP/vVPvKOAokyNeJkk1qAS+4W2Mh4IaTYwh3gt2ZUlqhlcA+e+43dkvKfeQ76x0FK+Sf/WAnUjjM
Kz55KRLfiVoOjlM/pI4QuOEB6QeRgwr1cEkIf4uU1Smay9SYGHKtRg/Ueh6vpK3tbn7md6dNT/dX
7jeZMsDkNqZx8LGhI01HMJaLT60WGw9QZUiPQL2SawbqKtTu7WeBpWY9//NscA9P/Q8kQO06vCv9
vqdwr6Pq6aQXWDoRtxN2xwGlspNVEqiHJbx1d62juLUSltJILtyTa0KnZauZa6TiPKtCrQ21jM4J
6htxflz3I6v6+OldfoXsaxWswQFRXzg2Tek4ET0Z7See7M8mB7gRssuGuo8NsqDhJuZYKYgCaUob
wEOffh/FETVAJUQUxzi9m8Mbq8q6skMYGYbpbB98ECdzrGoGTiDmOg0fMhVmiLzvg+ExMvlP6cPy
2g8TlKJa3Qt+LSj16slGFFzoAndhQeHnzbu6diw72E2wRBuTJK7J9UhCXlbPbXo2SLQlbN+wzdgw
w0FLKvNiiGzeEu9/Y9IjSBNMkB2ebIzewImaRXXQKNTqfVguA9HKR9nclF0cL20ZCwgbFSvxpVr3
Yea6umjIMI5VCUwbKITXh+CO7IyAlk2kkfVbVAs70LwgCx0gGApMUf7clXQ9DAR+k9tep4NzLyax
YuqAcKE4wD7sYRetuyzAjBZHCPHFgAOQfVO5KDALsp9bcJlAdNTzBRJkg5Qu2skxusHSLbnQAHOd
Dfg/w1aEbXK/TYbAJFLVyLiGqLgbHNShqPT4C8SAqgIQYx5JtY4j8xGmZmQaaSOIh9uxI2Bucpba
CXlOUgueKsDfCiQY3Gvs01gwcddYlznSqunPJYblfVugiEY1aub24cSGuXz14JfEI1CWoyiPe/xN
yWRVKg1d3gt8EDMBwYTm8uYBhtBl0TuWgiYlbauMNDf6cTpdvPW4eBZQQYYnYCXiUymjPn7SkkO4
WOTqEUp785CYi4jGHaB8SKmw/34fK6CslfB7cBxzjPvNyyBadmRMF0vSj41HXZSNONu68QJrRbQe
an/8IY5GJ+v+2t+YW1/MsjT8FHW1NHMBwXdtWzCPymNQBQu57+bDvMi8+OP9qEOoqH+HtAblhL1x
nAX8e5yCwwdmBEY81uHeU8/+FDV2Nl3QrEuObOmbqPDQdjg/wFNvptv2GEbeieYV6mP2z/LEVvAp
O5OmblQFMmENLiYXb0454/herbud74Kd/NatZQ7kijrLlZvNs+6IF5UQOBNt3Y60OQBh3O+74q6Z
7lnQQbchOgN0WzrA7U4kzcyQkx2AfBKnyjBQKI592c9E7EyhZU6pRiwpW4QwdQdz4o8lTd7klk5K
tLpoku4POyggFwUgULNpoyPVc6LH+H7z2sAPq2fPp+ENtkHKLc7p6mB+PbBoepOtaNNvpUlUkppv
XFnFv7tMHXidHCqZ/jbCh0ZpRRzPDIkCzHdDATIwjI8aVUvD0Vm975pCtWnqHfFSWh2pnGIBcnmx
oQus8hOHHjDvP/2Bp77Zgdukt7cBDSD6qridRB2IBuMSv0ngySbi6oEO8MZBX3TjGqUXn1/9CSvR
POKOhdAu46UYTN3X5bl2qMkgn5xrp1vp9KtNjk2sBjs2tiL7B9NYBHC4F+ZsUTCyu0glHyLTFm0W
Re7rnmY4uuhu9FkBpFKIaartFZShcpAsM5iSaQinmur5PQJpld7PtW15yDZDr6/qqtBCM3QQ0ZZo
PBFoM1XtbZZOJ2VLfTXQwQZrZUXFpS6tuwOB6hByzjUE7UJ05oVGdMzmxrNM7olW6TViWqYbs5px
EJCxthQixNrrpHtoPVeMAnDuoMVkZ7OSLo3AmKogs+KmGLnH90tqWz64oPYGGwf1pkC/eHKUapX1
uRZUB/K7d3aLgI0LDuknx/CU1TgywNVIRRGF8WRhA9HTktJrVUKARIDWoAAX/wl5S9sTMamKx8t/
Mq8sHsna0CF6bpoiOENHLfPeKgl5266jzPtdEPhTLO24+EtKqdqSRFHSryOV7M0hL274jlalE0wh
HNLuQKfDU09FDDWuU3WZ+5mYMBAtFyNctJGiZyuBeQunYSdjoF1dDEPgwWl1Eme40nXEa8XBpOat
uY4KTaz4XNYU/Sbuc78kPy4+zCz3n6jPAFfW7WOAx2Hn3HVGEHkZyJ/culjwIHzal+3KukOLnrj0
dG8K/TVUpoWfWxstJ3Ewi/LD09UHHSILGkNSnKQhI/wtWJ15F9LLO3BmtBMSqebsU4nfX6iyUP7P
tQ8jAxIcan669i65KsAi7/kRMm1QvdtedK7arWbGvEcpBZBO9EvDY9wdEk7hqI/SqUNsFBoBnYGA
GgRSqqqg+glmuV0EMU25+DRQ5NWTjfuIj9YR8cOApBl+kUxO1MtfGspMOAHOFvye3CdZLn28D+/m
CX5VOASpbXpth9+qxr5ilo8GXn9qYDv4wo2nQjqsPew6B6lWwCEPrOIcDElQJryeqbz4QNN+T7lG
xcRY8HWn3EiFs33OgH4G3RGAAK03fFyTQU/p2uTI3cot4wcZ+2Wi60YqDQEvEPP2C0P1MUCC/X9M
ZJdXYl8Xee/f+MEz5yjhZyBkZhDaYmqpEbnb4CLzVe0LrWl7ic8JF3ofwKUibsVQJHuyTMrgY4bt
stucmZfFZfX7G96Dawd4pDbDO2v1acpMotHboyp+pXyLGECdwKO/g8txHXEJzWQfYFWgjE3Caa+V
BiiDRaOGkS+hobKvSTko81FnmmeHINut9P0eO3b7Cj0ziSEK1MxRvEHfMnbbpCNLiw+M0Auz4Nml
CXJe7O3fy+8mfQy91aNXwJJKci6bTmAwZv6pbS12qnxtIheFV8kwATfzE/D79IhpxrkUnxcgkuVC
d8bZl+HW489oIJ5O1R4BX0FaNy7rpLY1WFKDgQ7R4tDALQTYJV6ERWM0bi01JcM+rEh5KgZ1ZH+g
h96jOQKLiZDAA9oGgTjcI5hL859I6IoXLZYj/HSuwx3dN8Aopebeys3J5mlCEpdaocAkI5CO+hMU
ed3H7NH7mIgxEknrkIojiuotVLwrFVmaKZQhQhhCX30FnSoBbE80SjJlpOQ42DjasMYqbQfkgx1h
Yn3u2NYH9qX86jA4TSDIWjZs198ub6QX125TwiqQ6a1Q1OWJKCeeIZNJcH9zOHi3A2bpx/13xbjC
2Mu9CbN6Lpw0yAjHwwwMZH6yQ3yuD1f32e/LjulLkei56SnnNeK09PH0+V9+11z/EAZS3gOf4cHT
e7VQSq8JZUdrI/9v0ONNQDs0XNeiHYcAgSvWZHU544oLE0GiqO32ERNgrBDzUzFyZv5pVV12YIi2
CU9CYsThL8ixbcb5I8+FwsBskSrD1TjLUYm/wi39/cxtjX7f0nEklE55u8d4V5vbu3Q0Yqu4+8a9
MoiYzOJgyGz26g5YK3bRsGCpKtI0dNHDp6OVf1Y7I7r32zrxr38q+0voN//IG/GA2Ees4fpgXEIp
/J8Bh3bhSRlXDJlAcSm1zz54OuekTdT6vWM6vQqpGXW6932izYBPJ5xFRoGEWhUnPJdHNjZsyqr9
EPNa2s+n53m/c+UHWAxGD+IKgJKLzPQSzcBE2NamuYpsmi+sJu77uNmGD9qqAA84nUVmvuYkSf+6
XXBkla81rQmewlxOvOJdoyHvELD69d/LmxGfqAvTkq+V9gC9Wbn6lijubG6//+J8DLV8vnhXJ2t6
6H6Dx7A255kVfihwtDY5OCmYZow7R5ZTd4hxAQu0Ny4rKhxawTaNKjs7QxleyjDeYxB25fEZo9ez
4UmLQJNzzLMWGWzxNphGeMlM9OOIjs2ueRUdiKrpfX/pQZmGI1xBVnbE2hUDsUKpUDzpa+WX8unA
Uan+gwRz11dsWyAHKCMQVxLnfUDfn4KPxDXf9l5lWdE/RC+dMQyZHzpEN4xfI/Ma/YMOA5R/Rs3Q
P0U3C4/Xuiz5mgRxEUpGfMDVjXbPbZ7JxHj4FEw6eJucKW5lUjT99JKIYlIq1DjY2exb0fzjdnfB
SC2k5v4Mf2ZV7QfizTqc8V5Ca9E/pOPXMJDUYtA11UHONvAAo67yAbmWAi8ETPjzMFoZM6rhUVMd
CrRaLOa6CQvSjE3f7CROGc3wE25ImJYFGLzQANd7gqnjzyiVzBV1uNFU13pkTYETDVawmnqNc+1C
Kp5GOadyHoR9fiI39uklDg/l3Ho6OUHE7iuaTpi3SJr303Foo/Ngz088/5Ce1GCTzjfp4/uyofVG
njzs1n6gqVwOad2bqtwy6el80guL+HHhq68G8oUP56KnVfBul6mbGjGXb1F5l0gS5NUjXxZQHxRV
fni3dPLlV+eNc+jCIjvOtbzLatcLZC6mSRJPKPJ3S5lB34Sls87iv75DwW6Zj/xz9J46qvIkmgO6
zY39HMYYnqcvMvUXLBcnJ5/NX8N4uuo92KgPvBclg1DN9YDjMnXpHQhrymabUa84/4xBEZNW/JeP
vrXMrvfWJXEZ1Hh1HbkUg9+HK1lc9zUPut2ZGdT2QueURfB5Fbt0948Nrk26/eHGZaBMC39MI647
lWHFIJxk6/SDisaKao9ZjxKu2OdCUhtYY9hl/JYPqfaWc+nMlcwkPGi2RGyRS6LISuTdZXxiakTZ
3+5N7k2Vms5782P8Je6KZRw918wKyBQQ8ypZD3HwW/2yRWzSqgBt9J/Ep8xxtw862UFkhk6Dot4E
dPDIBP2lAhY+olwZzuCDGaHYMb3gmhdkT/3xPejzViLzh9CpxJx+dA0vCmKhgnPv1QyFze6f8rx3
HCSj5eO7gGDFfmrEB+Aid21vMXIiUBlb6z9/VuPC6f0DvD8WtfjrcRBA27pofDvH5mSwPQ9urs1n
UvS4iL9nG+Rgwb1iwnTr55M9n86G6KJstbVWCf0JRc3/o/uGKo44108gT7GORNlOaEVPoskcp+IE
7eA3v+S8clE5tZQcPwlefq8oCl6xR4z1Kc0mqRMeie2UEGkLECDm3uNY4kAQUYuLc3wGCR71YzWX
jWEGU9lggxFURY8Babhe+g3MQew8GR6Ss/Ej/BoqKhrWFKq6nirH+Exrj0V7LRLuX6vogBl83gex
fk5a8/5Mtcnov7RqXnzWoUxw+fZSi9E5ecygfv0ptM54SSkqm6gGE3tJ80w1ySm0FGvksxQzsagO
Z0AlmbZEHYwTpG7GqergiP00/USBXQRFCs/HAv7ftOTFfS63k7jy2d9gpB5IWYMiGcl3fZFJFOMF
f7an9Ndp49ppHn4A090cADYl5XBxOZqlZnnW2tWOWPwwD+HxC67DTAIviDuSsoKxNcLKGWOIPm+D
YMPCwCjvCVOTUrhXTme3Ab0pmy3U7Mjhgmw5pYb0tgAn4KA0es0VOK8GWTG53n7F11ombj/j53UY
tEtFJR/AwsLb7XwQHevKMhNHUQ/cEnLNbG4QB6u4YeEwH0EZ8NGXT7nKTsoVOlZBQaTESQsQ/EL+
UFNHAoHsd4BSQHrhyMici2loZZaN7HHIF4UjRuyFDgPDZ6tA318CCP8naUZ+EIJj8dv0Vp2m4q0h
DRPSpr63HOGxBEFTHNMR3tlyIJ8urzAo1G5t428nLeFKFZD05vbWIhQD5FjPSed4FSOe1o6cS6o/
6e4UNukl3x7BWozABohjzmjhNi9GVL1SwCrXWuptPQblKPIwOAcJRGEtK+vkhCwC48K/EoMvWsMz
VYWV/hUrFG+Z49Q6pBKogvFRJPtioAmu2HVb6BDrYBQaa2/5PscXAB9i/HBqk0yX1ScUm8QqkXXL
ncE9azrHbDrtrvd2C9G+sEE09z0oaIg4ZFWCKzzg7TpZ8598tQA9xIWpahXxBx7E1UZQAllbkfzT
PWGJYQteta5x+V+UsPlk0DBWmqj2/IjcC3UN+0/Gi8Ebu42+uUi31S7YwJm0Ocuu2ainvNf6amCM
2mHi+aufSH9P+DswqFlECANi5Njg6kbeKRnihW3i3FJcimywBO7n0K6pgpqbVhD1P+LiAkOyzHaa
2Rgsguf8NtjjCOZ1jLF86sujyz26RtpRXwqdswpFaJ7JJlcHmHABkWpsb8+BpNdAcEcBMqFxSGHY
DQCS/XUbz6leGS1YwydHfR8AN9BBOoC2y1Sciu+LKhTqISLYpKngJBdkoziwtn3YbFOUMl3gLsWV
9Zr0NKfIoA2DUjWXvP8cab7XmAvsl/MX6dWFCMOLbBW9nLhDhZHQ1B/ZITOJDFq/vAcUO7UIeCfW
y+R6MLhh54x9dWJJKr7ecVFO1ZRR9XcEUZmfr1ySiJpbjfSHms4F1leOaXAKvbSE2gTdlkcVVkld
o2iydkgHLosnpQVAAMOkSTVnczggIHfnVNlTKPlXzENKqGNOTM2EJVAxC9sTbjEqpv8+GNP3v0Ak
B6t2WYrKQmF6c43INFsYRXPyzgdwUJKkTNuj36tPXblKgC8BG9xjXzYB1ucwxm5sqmlPzchx06j6
IZFwOhxGGMMNFfE8etYLaCMxOZqUSi25A76seX6NYyof3rqEMk6Wv+3+9+H8K8wMD85IHRdVhXxI
VzZbQCbbxr2b4ex93QcWfM6wDWA4y7Q4aT9Anc8SSiWQCp1h7Qsrs9wls0r+FQswYGkAF99jGZX4
ADwz40yl9t3vlArdQJE396uy0V3Y1Tqv/f++F+Uc01AznIpKSrsv7Zc/A0Nbe5a94RxAchmnhb+W
4Kqfokct+2LFiN63D/Uw6tRJwrkzARCyAziSXlLae7ERA7bLlbvTo+VOr4Dz3aRt2JzoLAYv9Xzg
z2VpqU8M7iJw8tBaCpsWA6r4cOFMBzNDtuTTaEwsBJDQfE5RsciOpAArxGLRb6XoTuZE5gt0Vhe8
UxR15g8Yx3W4NhHNGEQMlkoBqV3oDo/J5/UcgAodCenUlIDz2g7IcnGGiAtKk8FPbw6lFgY9wnY3
qOUOJ0fdL16T3CBqzI4/3TiiHzchvbET0F/J5WnJGmEGMYtWVXB5l+BF99XqIK78FCzgDsTT74H3
hc+rB/1QBHDXsGO2fYwEX4ckRbsKHoHsk+tdpEhn80akIjAeDss6qHHK7spMkdVYC4z6YZ3OrVxQ
e7M5Ry+zx4McSA7e/Gmgfqp52H4FYx5ddBttckrczBIS4oydo4z++rJb70D9fqVFlMM3Nt9NlpS3
8o2vAjNIMhnNuIVTk02InRfn2B/eCXZpkzAjFBsVUHelEKfl9qxwH6Updpljg7gU1Lm1ATjXrtqq
bSpwLyNUgAW8s3tgI5vLrP+oLeVpvkZKKwqrpCrHIzpnR6PXd+znMFHfyU+OtZB96AtVyaHF5dMJ
CkKyBDnMC6d+zp7dz8JpRAb36TwdfpMGvVh1Ux86oyGbhjTLL8rREfWrU88HkaRAqBuSFUghdtNZ
NfEYORlAaIbvBIHxMPqyitOyRtFCpiXirRqeBN3CuD2ylIA1RfmDAfhTDbm9ZYEXkSmH9P/sSztU
Bt1tBVKPMlXxh8PitkN6QpDNEM77r32veW+RkPbrhfJbtvfueK7bJSW2kNswzVMCyd1gnUvCYDWx
SSawhGRMkh7SsfH+ykXcE/UCHLX2s39akqAj71JDDd3vqos8tdJhXJu85fih6mvj0bXDtHOMBnrA
5dNxLNgilBVBRFsVXnB3gkRGjVwlrlRwHNzmGP1TnbKu2MZnNlgMCxRWzsT46DRZWj4+cZcPldWk
bVsNyn2p5vK06SPDRh/7SpQPTlLsXTn0yvD+Ns8rpAdYdhAyTBhNqK5VtW0uppHnwMNQ7B7hMOeu
RrxS+l8ZOeT0JDvWwlmSIvKTVKFlDkQril2eGncoKzwb5vsJKQdnwBo6UIL6se0tPz2hDsnCT91/
TVqC7YU7WZaRrLsQeWkN031egqdIuov/q/uKesBdseummragEKE2mlCU8rDEmH5Jutfi7aHbCURB
EvwLRjZOASC4WJEgaq1KYfmOp5aJ6DAfKqcm10HdN9Y2JKTgk1PvzpxQb2SL8l8BQkl9lSPD3qtd
/MxFCUCdkNe9nc520p7q3svzVal1ujGtvvuD/+2oGmkllnKknQFIIJQykWteHlPPat5xwtkIqXaZ
NQI5HpbPpK81qRB4v4UGcCG+jvS8QawD8b1czGqr3FKQngQpuIDgvp3PmSWKdruP2a1Kd5JUmFcO
YZdY6RCsHzB6MmHSvKhcCe5q1/1pvkK38eI2QaelAdmh0SPzTNBFSdx5OcvUu5uBYHOVaXUMVUG0
lJ0Y7IXgo+l3vRWtGluK6kTbOqWYCWGVkV3KKPm2b4tz3BmPLfgr8NdFCyupHxydhTQ1ufpKGWIq
zXerhXxt9wzj1XouJfrhlpwpW+GC0vAKsh6FZiJhD1bgo7DAP6chr7wzHq5diLblRN8USF/EICnr
PTYlrruTPLKQ/ozzU3Tk42ju4ijwpaWJJhza8QMFrqVzNEATTnCx3ctEZJqJxj6rVm25mvACV0DO
C+DIaVo3mOc0w/2N9/hdQzjGqHqG2m4krnwjRBR0McsrUfVErSGGnsWtxmqUTXQRg87sByHs49rh
7bUvL0KP0g6+2qVRi8VHIpHUkofydDZmktX1S0oSt/gavmXV9u3DGIdRYf9+sAewE2BsNRIBNmIX
cCyMcAA0Q/t6WMi2dnnIne2TAX4e+d1H/kpT/P/+NiyET7Al5n7xib8MFA/aRMP0oadfwNigL426
3TP3XeP+6Y72C65LlfhQ+h+11I0AjovhysDFU1fwzPpEf3H4fgna50zEiw9v9N3as28VNTS9DkV3
F7f/d59WoMMvAvXN2nHfIJSGXIDkF9FlQqMeRz1CO9QOQEvsfdcKmvEkJkmtmu2JUf7oIfo63jNg
B/GkVefOBHLiXF5a1/wu94yrYPOrbZFOJl0rQw8FrMNwNyFe3TwUD+7A1f/NVGq9dlhwVUSxn7vj
r04wuAfikMveS2g63TMnSs5IeTbhaDv1B5QFE1xzSgfrOYIts2xVjyA4VXap0aUKxh+0LLO/wMnO
i679FPuiL1aebK2XSaukA6cEy4/cKzqnm70iWDpU0n+uNQIdttGKgU+fFD8M5ZhqpHCh8kfbHqjc
V0NNYeQUyYKG5v7gd1MyODhVtT5xAoPg+l+m8gPz2cah0CSdfU9H0HUw6ja5PCLYZbPFzWC7m7QQ
aLDjQK6MkFPZ/mlyUaC+kwUnX8EpPDhSpSFMR04hbLewa9IAdtZZKkkJtafyO9OUFbAgxt1uHo6d
j7HqXyfZTA+w5kbmzdSO3Zi+Y4V+HLDmBw6L3h3SDYqdGAtGEiwWV0VzetniX9r7bA1daMg8l8Ll
L97L40EnhGGn04NBeGOSoQqXAKThvZwAy7CKWwoNXX0l2QDPGNnBZE4Tr63ERmKLGgiLuV9UxQ7t
t4lunKnQ2KfENMVaV0QSyxu8Q4LUd9bgmO+JqcLdpqIVj3Z2wYHcJ4uDTbFEDP3+cB/Kk5Jckfnh
T5jqHhcaXgCBfKraEEZVDoFvRosQhnd64ZEc1NhGDogJBA78RjAWhervBn7qbHp/kjv0M+pj+Zis
qZ4dvOUNUvxINiYh1bPq5aRKO6+7dP7h8K4OtWsp5Gzmixt5PRh48MlrM+brBng0RuCaHOKERyeb
kKG0npROSsbIa8O6Ogr4lyoZAadRjitRdSV+Mvu7+FPtrZYiEgOlv8Kw4Oc0AAAk7Jh5/6IIzjrV
GYC5IGWOBWqtbV6u0GDzOUPdUw4P5Z3MQNUNkyhXTMrPfVGw/L2eSgB5Hd/3VE6CVg7Ypsh+yIZM
ESmRJ/FUaqEeuEz0rQa3ezvhEGN57QnAQzcIfVe4qiotOihmxOu3ZrxgkHUXC9ldcfXMq4+j201p
mnyR8A8cSiH29LL2qTWA56InaW011OeuCnNlMrke+15O77q96LGijZaPM91jVD+eE6FEgghHdivr
QYnvrcH1gVlH1F+S9EvQKuOJELHlcGKU6tYQ8KlneiIxiyTUcusrcSvjk+sjzBXf9vu/qMUgdj4k
xofVgW5x95SydB7yzgXh2K+0QwJvu2L/QjZJaeMaSjLrNMsdfEvJzY4nAnZNVWkMx5t+JhhjwajY
syuAxbVd3RhxLbcL8479MFrmLlQhJpWMlSyGtaFckAPW9sP3Ac181Q7BmBiW5Jhh9HlQ8QEVLa6Y
WYpiVYcMi3at3Bgfqf1UK3o1pXF2gws1utkxbzsSEoqYCI/60TZqFCaX6JtMD69D8YxHrumOobXT
3JW4d4sUWRXK+W70hq6GeFXUlW7yG7hS3y2ieoaF5sIzxkS8fvASmZBm3P2ERYlZMTQOjAxpks1C
oxKIx2sRAvRxVq/6qUoTrf+Ep+nw+8yFo0H9FoTnKRMnUQqohLXJJQ7saMgKohvlTa+wXnOFIBPe
hPAa4JK2ZWujQNkUnINA9ild4v8TTEfwC7dXnqLLAjwTr1weHVlqOPBs8lKRsisj/V0F6xzrX5Iw
AL2r3JaMQNkUHqrV3yLNqU00G8coFpAnZlu9rbRbx5yBxqmmWQ1eu7zer70Ou/A8SYR+elDEq/2J
dvqJz67dvvTBWghDa4WJgv34vr3HvXOiOiPllvm9uT9c/XX5yGtpGvnIWPbjBfYSC6lvfSTqmI7j
y8R1zfYnXX67Xqi1RxiQqkJO4ABiYJCpoS8LNYCpG8XnYB+ZV4FE4h86tJENOFRH7ssWckUFwYjC
1+JJx/wsmPOVCUE1rK1QqY0tIPZO9KdDQjzxSYrbfor5OuawI3iks0XQWWeHw10YjF3CsOcwdFMa
Xqm8Qe7w+m55ArYLuUfWk+J1Acv0VK0ZnjnRXHtGR78sT30n1ydoLLW8ffv/0nJNtGJ08JXmOl66
cUG2B37EHsEV3OnFmF4oI5PR0xNv8LUn+aJ1/i5i60ZafU9R3BvoliKhkYGHA6YmO3BDwSt22haw
mTvxdUfsw6zgdF/hiAYjGXvIHGT932b9X3BMjB+R26lOoubsX/2xVjQ+Gu8kUdmbhcMfpZ0SA/uN
to5jj4DyXpsfPBXYUyuilJe64UVeyzR5P6gkEbTs485r1FUWvI1iP57PmT3WrbzCkkupe8TqvPtH
LvFgQu5hwHPBpUd0TMPq+QfYNKg6axKbv6loXNVb84AoRD0Goz9Lt0hgLg4y51u8UoCnH5ghhZX4
dQ/BtJ1pY4zM7+J7/4fgTBhtneJ60sM3Df5VRMPLvWfLVKiolJfL/5oeSktjijy7/48sSo/KItXn
5i3ui+Jp6F8+e51x0GwFG2WnewOJCZP6ZsD1xfQhgtyZrtwuZr+bMz1ZLnxNNFKu61Ro4yZS3Sbv
8ZGse4s7SAL8iT72u+r7a3pyKOqkiOCaOfAhG4j4aqJPiLzUm5uy8jrZLSw60SmUHcAtfUomWFY/
BethL3cH3JC8iHOgn3zHHvZ4pZcY9/XPqxcPHSrjJNTZo3YDefd5S0wUxKSq73YiVJjyuVXM7ISr
kA+wK9LvXmhDLaqj68V9CiFPtgAvimZFERqHF0AwWBLwmEZo21rwmZLnCOgu3A+SbAOBAD0MgUyy
gFG091LCne5W0RGK/qyp2wXrU70f/afKv4hgtNXIR3zMWMQc0TnrZFO5mo3huCNhfkHUrQcl36Zt
zw3iLXomtb8ZmdJ4U+eRQBCOFYUF7UICNNXz5Xf+G8AS393CQBu4ZIuRxVT+OnPjuBTdD0TlDk9H
RlD1FdgJYhoKCO+gK25rmjDeAKM1iILp/T5o0m9YoG1VYUEu6GjqKu+5Lo1v+M+6mzJ+bjiRRdhL
5secs4HBa3jA95DWwdc2/AwZ4UOdOQYQq1SyD2RkuPEheHTrsecd6MEHFT+PNPBddUkbzjqHKWgd
NZhIAy36e98btQQ2NQi72ZThziB+lCKLpqPbtq2efVrfBnMTY97r3RUhQZTiH2tb+miUfgEp4Wab
2OIB0fyZyGlc/6KfQ+uC324GjVvNOsV0kNhN69mgVeQAM+haL0DOOZzqav3MElBWTNoJ1aTCviVH
FG5Fs2jUPgXun+cAH5xQpZSLeNZo5CEUGngiHUNmtTZqzAA8SBevvxJtK/I6Ldm0emMXBK+CHKFS
odBIYyK/dF7Cz/GogslFKLC9Fic1kuievL9qyh0ezgn5lfgYBWqPLETo85XYRTxykbUX12iGfnpJ
Ow3DLPWgC3IcXJusZusx/LP6OzOchDA1dSIpwEAM+JT5H7OpFudxMFoKtbgh7pOwwNYTHWHooPMH
z0tkSWawRzhD5pMOfEMOsDzC3JoO/dQ5wVYPL6VKoZMzo9Wurno5CqZp5g44DOzFpXul3Kb/lIM6
aCsbQBSHFZQMrF0vryN2fQW63YnkseaQiCLPKLR7A9DRMOMrj0/5uqzJiGVxu9kGk1H3j35XCG41
N0a/+dWp1ThoYwxmdtPXYxqRvZ+feePkgzc/ZSGhN52TjFlZK/cDG8YHjUoM1C8s/m2JEw5XWZU2
MX+av9DpwkerN9biJn/ll+40lN5Jl76Bmk2pqfqMqkyz+KYRaRrAuiwhFYRws2jKVmSMaHQM3UjM
8Uq2gV3aYOrKhaT8nkrHfEivpk6Au2I321C/6rgZhQokc0RgpxI0uWREBman5t0dDPDsOeO9EGwr
e+TLEq7k/g9OKIlL3OgJP6gAt03RC7nzwwgShZH0Fz8p2y/LGrVvQNVJv28Jt214fMM8odkNzBUG
mE4qzjEa/NLUnqYyE5qUyB9C5eJl5QUWHpOzcCN1+6ipAiE1JUO2AsyyPl6a8h4ZvNt1rXIomH/N
7e/kKsTo54o3kg8nftCsC0UYMCALEt6oA9dqgFoV5DbE+njrhgNDvtZZXbbJvWly7eO7T5zg3QW7
vFU4R+hRKuzYHq+xPlp+1p8G88D5PKvrsaYEY6+mHEAE6p9OfdyrDDuiaUPgKXe23TTHJ5ZvSlJH
J8JUXWq+nvQQKpIZxGth2nnWNi+N4T7zEzoro58Jq1HmuUbjGXc/bc6LvuzGCvDDUXTP+hUenxgL
MH6XIwq94Xs2fnEqBEEVjmFAwHj2FxcmvjVeQxMp/JsIDzIeW33IL6AaJoUqlMUZ0UpvRXzhEwd4
Pc8e+pknDvx8m7bq/6M7g4quESdj7dFixtZ5L0xMHa3i5K2rqcoeKh2W9c/XZvJqLXku+0e4OBMq
8saUKf/ufZbcq9cc3LELrrIPvP8VxWd04XIGmfXwLAjJZmaDut9+xRhpq873r6igNlZ8V6rCo2sl
3zzDvh35gwPSJ0lNsyf0YbiQ2KWSFNKz1aTtwgsvVpTOM30iYThRsSJHpJRyIjQXRwxKwAmSt59A
aW5GV11mv8AZxJgB8/vcvts3Hx76w8y6ldr7bCzQKimoQA5F+XiZ2tCJm6T3m9cSBeKk35dYN9YL
akoRW8oXhiMwYuDtsTHV4dicZLKG0bFa4Eweg0bZ+5FCRLinT8IvbO0A1epia6tRmPjyP52tf+d4
ABn0CEBNjoDTqC9IRaYKiIuEQwu3DsqG4SxrixifapbcnUmN4UtT9apYPFxvGX2nDYpthwxCKCUU
ThJzfA+bVOu2V2oEqo8jALenFBo2bV8o22ht6TFxBFZo1yPb/3+JbAU8+6q/zdtaJhDoLDvHK841
OzIFvXO3Xv4rR+lKuJxjaljpLbFROH1jXsdpx2Oc1PwT24+GVJnbync6AQ1mF9WxjYDP2HMgI8p4
KckeNVtmNJqTUosEUNhi5+MC5j4hZNj4elIVvLwfvmTYuFkcZqt1q4Y8KgRRSX2im/A20MYvqNlL
P9yatMJSeeLXQIO94MqzzH2PLsvMckUh/vskuK9TTPYVSeMHLqe2uJ12/mIGjuRSoj9LSFDifF/C
MzqQ3JALf7MnfVcsxA9g7GK7GcwXcg09aTAw8mIHVbEaQSkJmADceXobWXDLFtUnXb2uI+jmdeiW
7rGBVviPPEIPaEQgvwaCrlW1GLDAzOYwxEdePzuBaMd4PXyDLR50yL3MtHZA6/0fWIAlBIiHJt9R
cP8rf2vQ/qK+luldDEf/CTbU9cSlqcgn6AYkkMUBvFzA35MVUxJHARld5hZNrc8LHgXf47XMOoSi
SXENzRE3v7sUtVXqmGKYbYuW5k5xd0QXLiMOEjPl0RrWlYhxLgcXbqo78W8xvTxH9346kSlWffCP
gtAOlogL//33I87ntvCOH8l2ajpUvJQHqK/T/apaO6bWe9UzuKpDCnaNd2D13X6pn+hzhncA3a6Q
F4EoFlBeBD2qQ8TsnkTQaXd2mfEEbzCOZCcDQRE0KOAQg4G11CMj84WEfWLM4FBKGr6hlnTnGJma
VrduVf5xz4uCBe3kdci/XRZH938/0qagsAJbO9JdgXsmVi4hJHkKBpyAg88wiShenwXQdb5RoGx/
YDQlEWFpSFRDqs1Sd+F6cu8yw5RKEzq1ykvtEY+XQYV5+kOhjDobxEdl8ENIZBYfJG0y7cl0trBe
0ljSYkU2/gt2YayOzkg/jHdlBN677H1/eG5q2hTCt20mggOZgLqfNXrw0LcfgJGA5LgLak7CZ6bz
3gX3fhhUlbsRTIjGydRZqTBuyE1/hgnr8aw0uAWHGPwkiUOjDTjKUNqbV6GCejmqB+VlTjf/UYHA
9Zgsx4sGe5GexS0PfSkT/gv8FSfMqWyfRF2kZikeJXgWFVfFs0g6EHFJJ8mY4qGJlFt/QWwWkrqi
A+OBZDkDtTvSbLE4UmcOl6bS4EUIR9zsDvzXCMORGerJtXDIFRODZ2YO5706dmfoh5e087gaUkux
wpPwJsTNKGu5IfEzf9nyibyauzP+2C405Cz5mp5hmqrjAxDVAATaiM3vbtWA0vQUTUemtEIyD/GQ
QvJKBGvEOacvqcHKic4f86jFBV3ethrZqZFImcxRy4vtaqDCGhu6ymsVQtmh1b57h0CEj4ddXZIN
c6jd2zknREM2cCRtDjUXa95rrZqWOExfmuntXCUKuZoPXodwvAx6ozg8n0z3jMtZBMeH8piTB31d
gNCBiSzc06dc/DlwesWktZGLlxhhaLwigigKEzSHZ0yRJi+pjfq8pSn25kbSaT+rN0tHHx1wJZQh
O1sjPH1uHBVntP9fy0p5ofHvcYRhO6h5/Z85S6A4NDdOBvABKwzylIjbDjmua4Scuh+m6hgUHORJ
ds8pKswyZ/hT6HhnS57Kaoo9YyscaRSIDCBUpjJjlYyrpS1ZZLPO93SwXI2/ts/MPOenwNaR10QN
8DIGqmqx2MkdrwKICHrF5YMQ8PRxZXvHbTLeMalIpkzGWo7nZBg+EVWpt9eEERHx0VeIb0XN7ODs
pl0glUC6BdJHEbOjiGtD2hPviuV4dT3c1bwHa+4VW1tQseFSsEPdBo+qWrfHSSc9T9/zWtPCIBFf
uVaG85lqk9ZzQzcNWU5LDnHYH/tP/lTtIJszwxm0BDSi14mLqLSwZAxL7UykrCAO39pikAJ7T/IN
W2vyJRVb8atay69d+HY4i3RzjsrAseKJTgF/8xrkxXpWJK4qpaqYlr82dzWpRug+QP/1BPvUyHmu
22PmPVbCs86woPv7TW8k/7tr16jZfj/8l8iItKbgyv9ArAqxXvWRtnBTphSOb9ijclaAkiDvM9l8
eZfyxZTZa7GVbKqgzqdfxGRkjysApcjSAF+rFeQZP0vj5GlI387vRSROqTSxwqPkw+m26lcq/5hV
xCZ09ihiYfpZfhWI1FS0Nmpmi3RD32j+eq6Cxu+r9AgWllUBh0wKoHoBu4ydwQK8Wq8foEyNgCux
3JMrQG7SndwtW6Vz6xH67NQlyv91qaRFczO/KiDyTqetPy+182ExTmc5v2AQoRzRpJJweh8mJJvE
NDuiAhf7pH3ChtPsSuUEV0dM7/9Gt3b/3wpfG7D4J2TE+TPtbBBve+6q0ZQcXjJ/NBAvrBbisvoo
sO9pB0N5wGmmoOgJZ7bysBJAc9JD1+Fo8Gp6XwianNP/MAB5eVNn2p+KpdiMeytoDFN/e6oGsY8/
lErLv4dBVDTHm+ewbdMUiEJlSMKzpA7zR1saWOr9OAXtv+EEawDZfZ22zX5ao4jjQcAvf/dzg0Pe
pKmFajVHad9Gi3HRHpMJsTAIimmuCGYmbaeT1Z9aA5hrOfxV4mLkQ7O5zv/CISD+/9hk1ywHxkVo
1URZo9uxlQHBB9p2Ac4RR4N7H111Fn+zxxx3BargwwaY2ojeQTNdRyRG/hI6V1ro+ZsGL36SQD1i
kI102iEY92SwuPWUZZVj97+ObBZhBZwnyuoqcwYHixKCqhlo/V/Yiloqkpw7q/XxDRK+b4FzLiUZ
Mo/PkMU6qhu4x3oLVdh1nQJyXtk7VosP8W9JCwSHkIyqUmkR92zRyjdp1f4MSh3/vLCLkkbv43Az
AAtvXDDgnvGCzXm0EVOWk8F8O8WwKil6BTHlhIP2E48GsF+DgsmMRLiK4rV/QiYRC6i3voGoZnAC
MO4mQoLFUfwgdlOHnaSExnrTJh1z3f4FFr4u5tJiPPFOlKPUbX7okkGBKW50F1wkfXrdgZrlLjtr
SyCzXFwrtNihgDqyU6xpyLg/fvy/TnMpaRM+iPV19xIGSkq9A11rwjhtLNGfx9x7mQjSG1wzKgD4
BpEueDaXcea7uEU9rowPZabQ7rAQjzO59B1p2RpaykAH49cso7BYWvGMcyUcUSsOWvTqyJgpFx0o
CoIoht+rTZz9x7E//EPHR1fQ99ZPl+inoVkDgL6mrd1y1pOaSdVDz2E75KvpAyDNXr+nM4jom90x
tjWvVdS7MRqwvPE+2m967t8nTujwm0o1kOd2KJeu/vmOLpTB0N96aILEcl/UWr1hfCD7Q9i41aa4
b40K9MLCkkIWjv9L5H8/IMUo/xnH929B+UT0k2ChbBZwiEcYwFEPKOLFuPfUSmQUSCCOrgv8FnXI
ZZy3ftfMdyUrbCJtYolOxV3pAmGWCDN0JGqCMjiIIHdUBraGRlSPJOBmBaZBGqcFoJ3NRXtfkBn7
nly7HzyM4mPcR1Y5i7S9DEru6rd+51XkknkyqiErRgK05dmaG+7J51gyVprGt72F5BqZhbkgDArZ
cY34TJLt2uVElWZ9/fxio0WfCGbcX6b+E1lOewCxdQwuRY8k63nlgAw+QMnPCllbf937lJ9nuXsB
H8CySJkqUwZKLW1GFwkAMW2hLRQgWWKsy6eqwNUSXH6/2ZeemjTyjVyjYs4ggnLXHqOfIGKSOzOX
S2DR9nAtigMw+uvSb77dcT3udZiuetoFfnCOLh90tcs+rrVADx9j8u+skOrGn9MVAat4zt9wBy8s
aZ8fGgKcZFhV5S0+Y6OjZsvbUT6J7fCd3oXFL4tWldGHSkshbLlOxGWTuMVAcCjr3zzrejDo8ZgU
/gIK5r0LZeQSHqLBNkPx2qjeJ7c4X1v+TO5ntpiTpBM4E5n2usPAZIIRbNIIjP4BuPbIOoCDEscl
j3934UL3bOdY63LoTNKFINyG9m0412eqZq7w7tZp4cas3fbi0Brnb5Zt07ebPuI9g8Xo9qT56KLk
RB3tonFGd6VGfx0V3wxysiUvSh5D8TsWymmxAFX2Sgdbv/palY5h90b3ONoY7kIrZWfg7Ipf3Iin
j7/802JsQa/GZMKVzs14Mnav+hKrd82nfinM80lhcP2PMbJby5uWu5FjbC6oqLkilzyHh7ZDh+fR
0y48bjI0pTcsx0c5mEUCaqvPi0cVmlvgU5mzqGh76VATQd6g5cuxJcX2lUEvRVcJ1BCs8nYqx+23
8Xx+Q+rFvmvkYquBv5f/XqvPl2PV/puY2WQU8FmK2L8Q6FgkDxBEdDaaEmogU5UE7lg/VQNYOi5N
wGA4LSLTg6taau5TPwr84qsxsXc5bCNPqtza1WTC/79lf/z2GMmP094XdNBDq1aYM1nLs0XzC/gP
ejGu7acDMW1bE+rPja237Bet3iSesp2Mz25KRFWGzNEJxTkP9x5z37+wcB7zZomC7M3DNk1wAVGb
piC+gyHGanr0cutwUMuqBm4JbCZlYj3JFEkBU9bmcnUonOzmy2ge6qgC99W2YjIumw3vRgoQ/i4j
9rEO/2Czh0AxDCk3y5UooyWxAYS7fkL3brbMfSToOucr4ohhu9mgIguGpnUPcmFbXMON11YL3deW
WXnV/8AX4+XZQZWfrNsVH/jwGHFukpunxgA6jwWMR1bJA7oZP0KPBDlWpOhmcgY8u9mlsl0UOZaz
aV7xbSY7CfXitlR3aaBz5jLSBlJ/IlrUziBH9tGkSVTududMRDaySxRNR/M31wkxpjOHEVvUwza/
8rUkJlYDNmitFkbN8hk9w6BbIdn/HHYM0JTS2Se1qpDVZJ//+S6Zp6ossDIaQ7726SA5SgaD7W8b
XWMJF8g314Znb/Liaspf+UcLhIm9sGUeWQgJXPxryWHpeBZAKeFRqpBlaD89zSJ5UWq/QJ4+m20A
aG8Y3JrKMiEjOaUOVFDxp4E8lsxtX2DXgYexfphUWrg1jU3BhURvrjR03BSslYKT03aWMHOpGcbQ
Ze+QcpVcNmgpKYeadZKRxW/b2oJ3WXMa3Qd/q6VE0BGA5jYt87fnuVX7/PCVQPEQX/k4Xm2EySBH
5T3dlI4aeZgXKVeSM24hHbGjwUFGJj9iFE+o6mm6ulSzn2D7RpAJDlgO+EV2oYKAuhWGljQCkFK9
U/gjE2gRQdrNVkzCkAWPbgum5l3744UP879s5UpR2/gBVZMAzDIc/guuhQP2UhO8VA+KoptLDD/Z
08BuC3h9sDOHP4p5hE3iGubcZO8Ln3Nh5Dit/o2dnTaVHVQV2wyO7sLJYpdtHVFvC5sjhTYsDJWp
mnkSg/cJhJ3s2snCnvG/Cr1C6MF8w0CdzBrMUgnFALEm3v90edf/MbJozcK0Z7Dd06YxO55Zxnzb
rrD+/r5bSpvP+/tv/2a/QHRvEGH4ExqZYXc95qM25+N/XbppoDklphkMCWF/JlSTHaSrb22jQ1Zq
MiIph5n30mUm1vZ+2dlr2wc5+tNJPnmqEqBBst92cFuX9SZjcIjFywj5F9KYCIJhnZ/Y7ZfA+yRF
dCM5s0gHzUzZ+MrT+roCenppSmWDs34EJANPGuAaQoKnjplywE/aHwy0meVaMorTTCz4Hn+bdIfw
sQgDNtVz0qkWWqE4Z+wo50wSasLmpxZFbrdrqM5/xuCU8eUOMzvWUHKIjiIDQIwxrnTjL5/2wW+0
X9mM+Gk8uwxX5YQQ0U0hLx0fWtcymTql63VpUmFW1UfVCaVWNDs1gbvYUhOHo0SsCv2HOgpM82CR
sJ13WOxPxF3yQRjMphjM1FTxPoDIcBz3drtOjx/qMtEx0qAVpG63uyQzQ/FMtp8M/n3sZLcfV1qm
ZRE477Nrp2KXC3cYcmeWOFNL1r0W5Yc+Flz+k3kuSXs6QbnXBNkos6oanrLKH26HgP2/MPK77Aa0
huPAZfITpEPWfg2y62kpvPhcx9E17BLGt3zsP9Y6HgORGJc0mOzkZEgnSuicuKUIfOqewmGFQiOF
dKvhLSpO2LpWo0so48L4MEsCf9o57XXX6bzbA6+ewfQLMljn/0BGqPYjM2Ho0DmcFPdTb92EDWc7
DrxaHHqN6DDYHIAUy+oGUn2oPCDOfs47O2FtRpHeBap4iby02qxjK7ag1+xKJi/F76ZCegtakdKy
pfCz8M3vC9fCq5vSgmJ9OWOS/LhwM0VEeIsTUKV8wc2ebNaicGoFZJ1ZL26FNlLOl8isdosrEMK6
u30DxwINCH5VRh0D8Rjry4Hfs7q63xP+50XL1o4NgVOsRxZMSgrgE/0ciFrUK1I20+k3n9uXj4zq
HpES3L+KfRzIhXJF1OAy0smwhuo0jwvc5990hJWIvGtlb++/WbRAi2Q8Cu8gBK5Y7ByNmfjhcsmJ
+h1dcLVJj61SnoUe3LG4df/fH1XG1etY54o9N2eULP1yrgBG0WXTye+qEdeZ/ZdBDdiSQW/+FJOj
Xu9rhTf1Cz4uaOUlaFdsAcleQxvyeHAYo8dIYuoc1CBZB0VXmSaSJ7Ti3uZL7v5gQ+QzIg52cRRb
SjtDrOrngFqslQEPMSBe7Q9EecA12GzTECMlWEIVBX6j2k7E+hvkYNHfFFm5AhyOBRloP3WbWk10
NRABJ/zCGW5tNUZxYNQYf+YdyxYwW7B5dHS2e2WpdAjt6EHRaJ8JsfGtDAyiGPRnnNQYFDJWvVBg
OnhNPRElJW6P9eUH5vYvOwqDRLdfU9fVmoyz8DcsnVIY07Sgc78RbdYm1bf0YxlrBnhY05jpArLZ
X91IvqYEbopxKFVJzqxSeDeUvCYyFe/G9omHgRxebe9X7yYNJlNRnwLx8ao6AJkCYOrLxMEFLZo2
kVm0o8vtC8sMyrc2Wwl4epwZpuDiGmLZIbx/Rt+2e9qHt9X+qDSK/TXvPz66+04L/K22QHeQojrA
1b8pgMoVxOjikUl13n0rNvnPM/9hkeNPdyexMPZxeEbrEML/pGIgNDLAWGVbK6hCdP3VacUnkHy8
Ma7EDBffUvyqPNXBYYAbdS7kaqqleFGmLZdqNbo2R5PWQJWYLOgibHaou66lzAQgMqXaCsIwRJvI
HHEPil8G4qPGtD7V/MTcwEwSIYJ8X61uhez+0jfGBP9dIDLmNGYXlI+0UitqD72nG/j/I5zbkL4p
tEoPfBppTOZwtxPjm06tKY/hxY9hyS1EroEfA3eD/zbs6kZsb0OIt0gYsHk+iON+p9CnBfj7M3oI
Y9tQCwZu7c/Uj2urEM2TlIxIfdHlqax8FFG2CPk1G62sDoO7ZguwrAuiXHJ2rLrXbMJUe5p7XbpX
JoieOgPwAYFxW5EPqNOJsZrCGvW072eMEySvwGzPgtnYgWLUFX73xqg4vEfQDA5uLQz+1pxz93C8
xQTNNcSl234Su8NNJX/xlm9mXV6HyByQb1rWcab1AXU32MVHjdCjPxR7OBjt5u7LmIn7dsMa9Wv6
QsnsXJNmO4uvSnRdSeoT+q4OjH+2cM7ZwSxbNO2l0e98wwpOO2gnNS+oTJGIzhPZYWumpfPPaqX/
A4+UTBtOO3Gq3ltIhIz1Sdk/D9DPkr1eew7T6OR3GwyRtSP0CUq7/yvRyE6gm60JFZe6nr03nt+l
Xt28rUOOL+Wp+TGNhMjqzyGznnngTTR+vgjPHjNcla6Q/JBlFemf6Go9bpyagPMjGh6efujH83bk
vhFOdt7dIyJSc3RXbYVf5oVvtnHm9hs6mUTyVrJrLJSzElcgZoNt3+lisvuR+6VMkGLw6Nzo6OXK
LYwRw2JJvbDpT58Fe+5SkbGtNv/3MqgSgLQzGHyNeKUvNyYazCkQdmYozUYZtN528zCJ70PckWUE
c8ougJUpxuEAazKtps2ZHnrCAGx+soSWwkH31MZe9j3Pq5OVPfJQltwOwvTNaY/SCHoRpx4rLhUW
WyhWXoXpmRXJzwslOSgCvP6w3bncebCp8HgyrWtdS/G0wRGrvTyqRgbQsbT09XGnWF2jHtd8MpJi
UhvHEM7j1pjxNT9JUvrHHiNksJFQa8mlDGQzZnwMLVjy9HhPyD5lMFpfphJo19u+Jx+JgSDsRv28
KEh3igFbwRlzFtbpBmhnpqN8eei1HyGe7ZwXcGihUpwKsBpsl4YxZyAL2X9aW4vQDjtwGqCRVETG
jmF4xSybY1t0Qj5+XUthjXqhWCnrUxndlQlWyBVSHoGYUu9QmQ9JTS/GRwEWo4/mM04LINlU1SrQ
sxTMHksNd07az1hP5F0VIndo5PsG24l0UfWUDa2PNsxmxtso7ICi6P9orQoC+oAf08J8guEyNn01
XYfT3AHhmoE7JfeQlky2dJxHTaeRm0IscVsR72Xz/MA17RA0Zv/f/HWCpy5k7KuBpbAQHTyL+CYn
86wzj/6y57Tqhyq4XlT9m7rIDP63lIvnjKCogMFA58ZkQMM1nOXd2ZWq6S0RMFfluohzdrDfZAS/
HRyr5iI0TCIA1gmTpPnLwcI/qSDHZYj3HRr2bb4XTS82esKl7dq4aOJmyOECGoHim+bF3xltWfpy
yDwf8rznlSAp7FytMUd5N66TVHSd0xhu5fJ/1YYeSUxyy8USu48UQ68uCCh2Q47jzFi7ddqqoEXx
J9n+wJxTfuK7YARkpAzoBrankpX0pd+lTkNuy2HRp78gRdGyAmy8yvhrmItgKuSchX/bszk2TJ/b
mjDJh0NAdWi9wBofMTeMUg0IeFaqwwhsC6A7pGVJxNGHyrdByh062/kOO9isEQGtgg69bj2UlZL6
c5IfBDmEoYt4l9//dNaifDcAxTYoSz2f0pyL3ZtDLhbDaCaFNsNHVN4/43vTGRm8t5gte/JMkDN5
usO+wjJKktfh8RP3IdIcvon1z1v/LUC0FGHx/VhJvzXK9AJFTmiMmdbklOOVFk/RNIzyjSWClNk1
mVgwcbAB34plV4Hndte6M/6iAWedgNfbSx10gViOkJ0KuYp2hKkBq+w/2S+MXSB+GAMo4pjwq+Gk
F+Q1fowBoM8aft5F+zBJgNYd+4D4XVlp+liUIZHFS7QXwHV9qoE5fHA9EtkVRhLFHM1rjjBtw2NU
2HwXXSGNKee0N/evXA0hR2Oam9oPvtULkfcVe2ZjrdngtHQnM+L2j9yO65QUYiGVU0nXVaxCghH6
Gwq7xbh4eh6/4s8+AT353ZjTPeLy4a7FYUaviozZw3JceQXsJ172SWNAzOB1LGNk/COri25qKE/4
5soAeHE7g2agb7eAp2R7QDCy0b36OiL25itzVYcbOIuFl8aaGs+9agXFAZZn5lS0p5RSbv4hWpqv
PpIgCsp3zzkPzO7yZXKHpb2F+quukwXrgR0AFsIWGFn1nzwrT9t3LqZTWMhKhqTtORpMtQKy9xR/
3w+xk6PyHK40vK6tEenaOqf63uG7rxbh55BbdYC7Rm5n8+AoyvzDg0c5krOl+vsN9sFL66EfNgh/
DVOqQbGtYTBtXeuO8GZK/uhqN+ydgS/1dTIBPZSS0mfrAZ1DSJbAbAIUo8o7tF9rN71zntVfK3tT
zMoHOl84Ql7WJeRB4zsADxLb1hS25Ru3P37siLaxM/AE83HzW0H8fqlUUpcUA8x0JQIqussJh6RP
tkkEsUTcpU5EsTKpmyFIm3QjCnsfA0nh2tefMqEJ0QpPs8d5YZs2JxNhO6tMXkY88voyF/L2enEJ
/p1uGNLrrlUanDUz4NGiPxWUPJ4HvohzDBKTFmY7C7v/idRzBxwKF0nSxBcgORZIP7SnvArYuUfB
LVzTiwlUDefrc5kcPZpLl4uAuy3J8ssG73QMiiR1vEVr5okYvZ7NGYaMfczS7THnCuplPn3Usknm
O6l+26WWDk4e9pi+fbQIVuwEptH/B8FMY5wW+dgQ1ilFRX1C/Y+Ca0DaW7+9H7SF6macmbg/aL74
SFHBOPltF1BJs+DQDt4BhsG+scERUauYHXbMbL1LLNALaFIH7A+NYRoAaXgeGrf8A0McQ8IeEdY2
wpaojin8BaQdQNVWE78VL40BZkP59ODV5mGve0U0oUOe8reLxGan8C9Kins7RpW6jRBAMI5tY7p/
K2Qw0X0oFtPjWRjx4A7AW8vJtjTLHLBoc7SDLc3xT4gCEyjK2p96DQ7+x+DJZwhnOWg3krpIeVsZ
8I1gn9MmeGTkFBC2a6eMwgJT9rtpE5sr+nLpOsMcxK5AtVbByh3jwW3UgjXgHyFTJT9TByiPxzxC
nAO95LEeTPEE7JCGTuTtpaq9Px25meveF9SfUlGhaZJSLK/xoVaO29YxvV3/xQoVKMfcVwjhk+Jr
ep9ITqaNzeEA1THKNaaCDxHQMHUNy2PX+y64OZp24z1CF9s90jREVpQxbka2iB/EzQHRTsFlJlkq
1ZDpiyIuHIrnae2yRW83oZFXav+oz+y1XgHOC0vTawyLAxxiHdzgsla/N5QZT10aGnTSth32tDX8
s0k9it3ZvuhnVmvqHKGlGauxaTnSQUyC/7lHxS74LgcRGI3XVq3EfLyKcFL1Sz58/quRAqrD9Zij
kw6hrrL/TmAUq+n4FnsfUPbRmyHrPpyJxUrjg3XJaqhadtZlTA5xiwfLVp96Qydgo+TeOQZDfhHe
mXLUv2JEnAFRYz7j92INjs/UhqD8yCGNhixuvoBXFACXit4ZOJ2MSMiwUWXTHIWMkXQd9eXYYbZF
2WIQV+5QP6P6O1FX2CNMBaEk7NRmnRWjWRoQJ8nFBqrM1D7q5Hq72Cji/AkqEXn0ZEJIAaNJN9i/
hRFezrJBA12wEQTR1i6AaDm1NMVycurPzoH036fW+ABc9WCaHhoCBUEc3ITo+nIuIgJntVTYqi8s
eU4jN8DTJmyucoO1b9ZMlhgbxPM4cVz6m35qtIL4aGh3w7Ei6KLHzaTKGn0ttig881qNlVNeFKyl
C5CP4fNIa/iWoeYvWL3t4NG6qognHvEKUODdLRAtkI1BShEwRt+jB2skjTEMZTbdXlMG4k2bcv3H
EcbW5KHhacw27/rCBFtootDyaPDYjWyMLGPTRX1R1Mnq9cZqK8R6sXvqn3YjyvfRMw5w8JZ2PYC+
0sygOEZy3q1u7iwUqvW12Os63/x4+PkyFZWNF2QPNHll2p2it3T4RBBlleU6LErJwlQ3oT5gp93K
QN6nNhMJvtA+cP8u1rbVEfjRlsbFdLE35YCk9gBcHvlID2ljp2on0TGH3i1IHrPNuM3BXqiBDgFo
iWEFThDcophy1ZYKCMwTp1aqyNJl64qAtSgkAjAAJ++dRw2G50VLGePmPhB6y1qVRGAd0cLm1X3M
kdV+QTKO0xzvyoOTHMANQA8UNYzH1v9DqND27HfO16f/2/fJeEzuxDVU6iVbef9dYcY6TTcbZI+l
XzfQ1XUS7RhhVXj0zCZSzmFekgvEVKjkq4LHcRcTe3Txail3X3srz32UlM2ovf6qWCd1vBdWomH6
7tRuNqCDWNYstxmWK2XBDrwMB346RydYhjns99rPFfyrL/yA/qQxE0WQxzUV+bdWQeKzmx2RwfWi
2ypLq+Do6oRGaiNf2PRMyTw95xvc3cmVD05ir+J6zuVIHxWbVtMWTn8N+a8YYAhhRnhJ9P0yClh2
zkpAq1ZGnRj/WotWbOG4suE6vRrxBLkfE46hz6VQKP+/ZuNd35uePsar6blWXjZiguHTCwCGgnn9
uIUELIqUewdcboXNJPrvzdcaD8HKWqKHeqoASPo+EFudNiWCmvwTFBpKbJDZ/TOPuSrRGWp7IqRi
gPpav7+d8odWbZVBh8OBYcKIgAqH6bZcdSS9qLmer8+jDAYQ7R8BulP7S9NjdwqxE7AfHZfCFt/P
sSVB/o4AswfhoES/FvJmDVmxlugVlkSHXV/JT3zrPMAceNNk1kmqSHahGO9dLzQG0cBpu2UW5u0I
g0w9IrPKFIDrk3BDqNNrigwlwKoXoQcXzTMkuhW/t93bv0sX4cC/0bruxwAnE5N2nZS4tABQDCcD
kP/K4UCqx1b8BgRTNm5J65AiTBCElGz1CJBYa4kTsdcmzfhZgfQeitZjqoSOcIpal6zSbY7+Z21O
Zyb/Qp05LkyX1liQZPiNm5Itz7eet+gKvRO8OcFCCvGN4QzgZY8AcGyotf3ENT6bLETb78NlIdoV
c3CKxpZ1CUxfrxANtQjbGEjx2uwN3mU7akxTUQn59lATiptJpFF2Krj6UZsxYbzG23Kq1OmCLZld
1RGPQEonR2sQLcYTorQ9Or/KhWXqErLxO+24ScrzBjZhkF5+UeZj8VLAy3SYUQpiFy1V74Lm4/LX
wBlw7nQ76D5KJarN19uWmryPv4s4W4ZM0nPssZUnd8bzV2ZiaQTh1O8itkB4RUzlxTd4mDPH8ji7
XUm34xjnn9oAGSj1u0+Y2PXGxdBi1a9rikO4O+m9I4PE6PRDLw7B+2sbLy3BHAYwMkmOP9nBMvD6
EEDfSkykb41CMkrgQoB2FnvfnqZWQ6J3XxLbfUgIQj/mN4hZorIAUqLrcLcCfAoc4ZVipGyDIhbF
qtvhmdk5bCamvqjhvkMcPcK3dt+mn9uA+q95iq7kucNHnO5n0PPgkXdGmy4Uuqi6g1cFm1a0ID5E
IKbcCKDb8BiCsUgoQFTOgCsdDYXVc3y1Ez3uwn2gNAAoXPQSIMLk3Zl5dMha2MOqTFGPJAtzUvYa
e/CCiLH2cD4bk9hog2hpn3aGekUwllX7a2nhz/r6tIXdcVfu67aEMZtp/6HywX8Khmt6sHM+kfe+
JHPjrwxHroFbBmRiGDgLtyZNUYAKFH0ogHk7jqL9na4NKublyxl32LmO5QxT3zzGffIWrs7xm937
xJlNG0whlz20zbb8MipSqJBvVVKr9JcgPVt/f3IoM4F3T1zYlcLnvoX00R654HMOWpSTdeixyqZP
QZhpxFo02zy3KVeLsXarQgOTrZR6HJWtVzny4YnIp60POPsEqvXA6gXDX+20W5tPe82IdAJ4hRWk
fKKMp2Cr4PSxM1fQPZARbM58kFse2lWREPFL8i/UONjOoOH64yFOThAEjLNUjQZE/AQVoqVNgW6X
9b+2pWHWRVTlOQ8V9SnZr9XU/LnQcE9vteMt7ZumHgbTrQrs8920iiZ+DSrjImF5wtkuwaZXxBRF
k/Q0/uQOf+BvV/mQ2UIVc+UF2jIDrJ/yawq4sxac2gVaUo1cMO1G+3RAuU3yioaLdrU8vJiWAQje
0xDACT5YX9zfpsscixznrDiLrVxjW6xij60ocuqMU/ywXu98ucug77k2rgHHk8sVLsJXh/i9JnE7
OVd/FBV7NVI9cqKr1vjBgePgX8eoHO2G+gWXb8CNfyxej7ilqcud8mmulQmLhGQ2M5ab6XNSWRLQ
YGTTk0uWu6mB1ug8iSGK0TWVrcouIGC7yX98wPwyOxSaI9A51oAKqt+sh3saPmQtLLE2aQR1Vwn0
jZwXBF4+5yxJxpnU7XMRWsqbNVEQkJ9DEGVzkFSqvgy5HknjgqBAGOOdr5l3v8hhPJLPkMj1r/6T
iXVYG+9paTkb1oFt5McBXF29CybUfxnNOITeHSzugkgKDYKX3MC1Zf757CkbpSMR2RFGWpTKTVEk
X/nGnStZNtuRdeXBMvrYlLkreAuqxzSaKLDPaeZBfHVRy331LbZrzmkt1ih0wkeI4QxgAmp8vs3O
gq1X7RtjeHzo+j3DuGjSLsvcQf5SR74Y3Fc7Wzno/weo64U+7vtDUWVvn2PF+VnA19Ge7kA2HG32
xix7PWxrEHjXvkzEaweiBaTzki6qu6YjAjNG6BHytjJXxFpiUR0HcDFwvG79Umw3RpeYNFme8fkQ
/K02EWKMLh4y+3Zh/uQFbzGVU7Bt+3wRIm1RQh/h1Gzxu1OA21Ulm1iDn2G6/F8ENoEAr5RfgcOj
3V6DnkqkrcRSyNzhxUtaRvKccsgKFs+whANXzLiOKhnMvQmZ3iJ0zb3jlyhqCdKhWgZhQ5nACE/N
xANoR14fioV10X7CsIPvCQhyPkdWZYMyhdbqE9DroF9ID9vAdITl816z64wBczs4/io5Lqh0YoUo
uTEx3aqJ7/L28SLtTNis2KLexMIJXprIebXiXpMc6Ny0T9N9s4XIGxQyo5eJHz1zPr572MUGDK2N
RtgHBjDBUsGlFGwMpyBOI3d1ihTUnRsiNwZpHKZyIb0u4zZW/8J2WXIr6AO7vpdHl7gacF8AvnnO
3D9OVO+Bpnr8gorObdcdwRLFHBhekP77M7g1pc9jiKglAQBqtMiUhXFMI7BqdItrzM5P4DNzcU3q
QUDDFQ/+q0Yu6Tl4ga0SP6mzAtNpbNbXvCkdaGbsxRYgSEl8vKlCCMW5YKb89ze2Nop4sJaEzO8W
ePdXcb76ioKkGLx5symq6S5hC5TrtuGYc/uxLxJ+3NDaJpUsWg1onAD3Visa0ic+0IhwBJi2k89P
mafiveW9YsQC4ohbGJGa9ZiIIJo7Ejhs3Pju0jYbARj4rJi8f93Icveax+PgvDslLkS05k5HCe9m
lgz6I1qlaLHXx3EzRRadNfYWWN+U/f4tZvRF5z/OoEUmFz975A1dyfK+RvOMAtwCHKF9rO4OdQqN
KBzofOmMHnx3j07OQF2MpskSH2CnVMDyFz65hOa8zVmGbJHMCuYjHrWAE14Cr8AO++3lmfUwIH4T
15ClbXxBHkmse7mOypqIaE+/Lk8wNWBBV3mbYZt8Tm6C86Bhj5UVBJInHMMC3BUVPKhAMZ7QIzKv
/fhzdf8laq8aobdB22qrMauRjv2RcQYRoVq/cMrPPYQoHQViN0Je338CjtsTjcZQu+VdZEubeSs8
wHvbBHu2EG+xQbFvOw1SGnfekOA11seNHDQw7ZA6swFCdZcNPLQH+s9xXET+BoF1Lqu+Bo1EwpRF
43Rmob1si8S+PTC235+zS+wbaEdlP1VKKZn15Mt8zbFwoVLhSK/Jz4Bl0/iIlsSn6WVsWNmG9vhS
2cD1PwviQdNvok9XKWaPYmc+BjBZPvEuYMEZcQJ0LfURxkV4OtYXY5jwqWD9fYy7Nc9k++/OJCh/
BzG9rVlrxr3/ydnceg7FhmwBj8ismWBmMGDuxvvM56x3MBxF9xoWaoYn9j/Z/rJMac1zqII0A3jN
jLtLChH8H0rmQnnjAED+JqoXcOma1LeODiqDhf/dz2GphzI+MX2DHgoLU1E9NxmV25FeoKVsr/Fq
gIX0XE81WxJEEmgzjeSs6RG+MqUbeVhA+R1GgrUnkpu9OSe7wwUKOf/D9qflecKZjva7NbiL0csc
SpL4jzGyEV4ZqdnEOr/GFFHggsG7Qr6q9lD8rDBO8pwwyZ5cGDz7zAPKMj9skDeyEhPEVOgcqSOH
C5LhfR4T3gqH1+JLkkVO1/Qt6K9N/+MYgPGUmPhUjQkZxY75qKM0w8egAg+0dbcdPrwQcP+0rP7A
bz8aduMIydS6q5ck6vqxvYO5dTzxHDcYptVm8w9jmATxLOiy2Rzae5O08dpzEO+Pj9SbM39hcdWY
WIoE/tT9xwL2vSLyalkcxkLEdRLJXaVHRoJg9ukohMkqD2jxaA6cXaQ6eemF/1aWLYxhUeL2W+YH
/IUKbL/e1K3pA9b7b15KvGC6T+ugZDvEzbQuBhrur8m8foEmL7TagkPw6f0I6ptjVJpQcR9Z/82D
vL9NAcwdTOjCXJ7dYRDo5E2dcoqrUlHKbOZ4KEFiyEeIAOVyOxDrIrQt+7FndGP8rsBplZXJq+mv
fS6O1AQx3jexXqliL9LRvoJQlEaFK7/qVKXTX4Qw6vP6l5njMT+4oxMIqa6fFRNL0ccUTw/0fQHi
lSh4ifwoMXVvespkJfbY3O3VkU/dwySRmKFLsLBaY/cb8jEQEJY6bg9aySHa1kg8gF16yRdnxONF
iUw98nS3UnaOhY4FtnMOuOHdG/moGtjzavFDbMsYG0rsMZiAEn60iG/UOL31AqLy+tnB8a+/Lv86
s7k1It5RQ1mf1LmM/ywpwp5yrDkpTA/ibtYAjVgp70qCehNpmg7sPbXngICxrTSj6OYkmHy0/+F4
pHnefNicRvjcAmUAGNk68rOMDsWLWe1D568HF+9BrJhAKZKhNPPT6C1gQhNr4Ye7Z/J/EIuHEPgF
AiyMmZEcNJfoisDsXs5pmjLabMQ/xhiA/Q0bRX9MbdJt6Gc4DHH21FdpApycvpHuxk9lHF6y6BQe
FvYI7W4fqDnF0YoxaMHFrcTAEUpQh1ne59bXDfrEQ/LLayCayv7F3glTs/mpI7FMPcxIU3nju7QQ
p2LVtvDoCSqhYFwHTTSShtLYDeSX9vCWz6FP9RPtIZf39PrEsGKSVPTkos0kyYtaoOefLdG0ijPN
Mh7poNKwtaSweAwwOBxsDcXmt9+93Nwa2NUG321tB/OLxN232BxQqsoofv1WvFuyzSvgJ74cY4xb
UQDGqlVkrMV98d7DXvtL3cXGtoWFdD9qZnDRS3zR3VR1r1v2r6bt2vU2ullsVc3VBLm1lk8bNp5C
9rFOw/fqf1wc7NZ62gL23BeeTiH8LGgysOuq1VRp8V9ol8kxg/ZjrXRQ9wipZrbSpO/2alBHSKJq
g/8Zodkp9VQgSGA3fJAEzqn/8IQo880LBR1Rz2XvRO0PuGMW0bO92pvvpvBBnfqOOhs7BGk1UoDr
mTZ+mFtOtTWsg7z4Yq/kiubSM+2Quc4H95xaTgENjRnyjHf3/q+3JDKlBnjvYWskL4qx28xWqC5y
Zuk12Eu2mUl4ZmyQ6u8r5+D0NPic6uouMwsbzORf1eYG+af0vPn8FWb0B5cP+sMQjJiuWcGjLhOJ
PcimG3phnqe3OrE5a3aELxjl8TJIKlUazHy/Jw1D/vc3mGtIxRWLZuhnrky3J+w+BindVBHSvVav
2qUg1ZEGaN/azyyDoV0EK2m/fDfA8Rf/+uf96FniFiM91uw02lY35eIFRZEO2AvDbr77eUqkWG9Z
XLX2UosyxiEB96JwzvKY4Lp4BLIacx1jX0aU452RF+Ch5WLrWbrlrvZty+tkqurdRp+WIYMG6lva
UHKXr2VgEpNn1yssLN8O1cerutqMff+eLxPVRIPqRNXxUxj/XSg+TsEYRAioraHFinaYuNIZfxdA
/OO6DMYIEM/Y90feL5qpFcnrYlp5FRB6oGwYsAb5VtnT9pf0p73jdN0hQkoMm3JqvoC0RjxtYWXx
qfmHIzVw2LkxKGticjbVeW1MmGiMWFoW8QSw391PiyOrq3EH7cOGDc85cwbP9jFoaY37CypuxgYI
14EXXbLt6vIwFSH5L4FS+twb73bdM+mFxgfxM3hXZZGQ/o3Boo5n5f3GMRh5tBw3V+VbFo7mv5s8
QeSyqPC+MFXXYdf0cdb9b06oDQLaAempwrHS9lQprhkEZesfQxvrF4540I25kDnZHIOFpyDV4orW
pJh18QS58ZvMWWH4UJTbQnlB7YNYbBMQzrJU1tgdOGW30EOySUF3OGxP/YCk4/MNFa+lytZVNLQP
FGYoHYhciuGmWxtpn3M+kXHAG632muKtCtex3DnP9KqUnO61sxvGqwZEJg7oV0JSA6ag8sHyKCpg
7QTXmqluCf5+rXAwnFaDLD7T2/vUpLjKNzn8GJCJu25HUKOzH0QoNxasri00iYiYqRWoTE0OYyEg
fOcyWPmIZO67C5HyczZ/bNgmar4d7YavEi/L/8OcBYAf49RmctSYAoAGwQAvtPOD2GqddsNYDmQn
IgsqGxCFiT4CYDq2yJWgzvVnleSEXisyf3TG5sYZe793ROeVWYy5vYop27pad7BdRBrEQqyQXNX+
yvUOiVrKYquulNPUj9NAE9ctYK1gUD3QmDEAgP5m2SYn5vXkeDFIK1N7y1NHjtzg2vu/FdAJiced
ZFWDpm5Q8RVgEuPqavTNpjckBAl0pKuwaisBH6HeNMvswAvkPo7nD3a7H4mSmnN+pW5+2FrS/v/1
C3AnCzLela1+VuofDtg5lB2jqVwp2FWusP6UcZy1zJmPOaCf3ilLjB8NdUlJ20Nq1jAYnNtJhclN
Xvol2x/ymMjcU4+JoaOgsrwBowaAcumxaiZGC/xugqGVr8A46SbQQkw82odhkaymDrw+lbH/cZ5y
2kQmC2aJOjkhKqAkFPIIDzEp4MO5lZuEb/fiTN7G5b++YLgvcM2cZjFK4iCJmLUWY9P/udO3VNDN
1w0D3fr6l/i+NLfQjY8aiU8a8DfqdLcIO08ypy5iclLc2x0m5OgQch2Hp4m1ysO4VnFMX7YbvPoN
fYF7KFiugyvUpiFo2bZxemxueUhkH6L1h0RK1u+G7OyPBHuQRgNu0nOHKKiUUfG1gl3b5Fnm6K3s
0aOanv9C+xAAxjBwYd5+ccn5gkQzCJ2JXIsJ7lapjqD2HIK9hjFJbWkbG6J+UiD6q19OpqJsYqe3
wIrE36lqf1vGvYMmkN0inUfR/XukuQH33RbVzjBYZOw3eGSsXlxb1ODrQMqT/HoMn6oqR4f8JLHi
m4QfgkMYtcomB9Pg3pvzLMO6yL0boz+f9jxSwsNvpxy04GqsQdBLZFQ7RXQ0j0q43rD8R2cVpPnh
YBlhtWPmnqvlJRwRDwmS1Cd++t9NnisVSY3CZ6yxqK2B8tN8nq2WJC0L+9YcMJsA9SELJDiiTmhu
Jaok6FoPMb3j62HKFvPVL0Kou/x1+QLhcz9tYxuAreROy/an4YEQ/F4uXNrwc6L4FtcbZiuJ9rS6
/QKEOOQ/cXtGG3fnstAFphh551azQcpKavkJUryfov5fvrH6uSYlvw8/meZvokodZQU4lB+GQXoP
cUCWjkSmJ8lIDcJDT5kWaP6ViVvdkPtAGrg9A2OeCtSwhMWWUM0u9LMBPEGRwNrNSeLRi9oZlMo0
q1N8ObHsNUedDdzNLXO4FqOsyhtYYCRoNtR65oy+GxKHBBzponWvASij+64YBRBxC0dmp1Q9VWIt
GAUnU+OUli+dWXQiiQ39XDY8uQaxKd6WxrVRX2wtWHfJGlWG/ecf+7gwk7MVBRiMGsuIsM0c7OTq
/fBlAhICQOG2nR4I2RzjCrU86f0DIDSmAOaMAS46IQFhH4R+xTqz5+H+v3EKiHQNVrm6yx+xh8NL
kU5UoF966qnhGNbKiDkUZ6l7rO6qf/7zJJnq5Iu/DKIeDn/zhpzTKg6BSqZ6lnE1YWZtzokmCveh
vFEV+bxVFQElvzq0KN2/Qm/SWsecZowAF27Dy0kO6Gz1eJdxM+8wcHJbtp4Nwjkj8Cx1j68Wp95s
i61P0GCjySgGCaVw5UFzsihAggmjXXPvONRtRXE4R6YLH0ePVG+/qbFiPhooI0gmNlQ7Ybp737bJ
WXSe4Vi3MvTYVNMriXG2K72TQnecCWlt3i7cC+RtCDceC6nVQa/c3nz3d4aN4JGPi9AJ4JASm1xj
mFqF6tiktdBlzLZ2ytlBftEdAFWk48m5lwxK4OecDLFEv8vrCG6olfUPfX9XOkddq6096Mxt53NF
pk7y48sq6bcihvfYOkJvLSUxCY0ln4Qprt78+H+uD9S7SCgA6TwZyli3Xh3sFtWGI0gF66MOx/UR
zScN8NLcy6mlf4wVbXU3ZIs68YKQudUNPz8by1S+q2XAoAy4tBNaCnTkYtt4um9q0Mg2ixfPIR/K
5w3xMQVuylSk+zCAjdrJxbElHQocnprNtoa+181jJTeNQQpU2WPe2Qw+dz8RSpDD77IaDwdZ2rH/
kIQSEVATYw/f7vBjmIgxIIJrsOqq0tVkmCk8LQeMQFMzRZFvZDXemIkV+HO72siq4u8gkV3MraVH
/LjDDGEEdPzEqPkr8LpjoCbQkbE776bJ5GPCp/R/9ACBHGHn9lT8dbYO7J8R2Ttgb2f1p9VN2ilW
Esi/00Cy949XxfIlwqKn4hy6Rv1EtMfT4sSu4cOlVSdo1TFaHUr308fy7m7TZh6qVF+uHtki9pi3
T2U9OyBHCezPyeRlW+g5UpadPfvaCGizKieD5WpOsiJE4SimfCHFkIb522FXfEh5NXJEPQExzwZ1
paxxHjg9Ixe4zlqQ95R8N+/xfq+Y/m0406eCF82TZfXVNuoEeTK/T3XLS+7DCRGSJFHfSFPTt0iE
7kUb/oG4PpMJmlD4ULyGGix63q4EXlhIDd8UQR00LEAEA31qqyJURUMxwXEy1MJjhGxwjhNWaLL6
eKcZS7FglzT2pnR+ftBgdrWKl9InM9wFfdmsfRDgvlPD8pBBzSSpT5As3/uOCUKBicMos99ybl5Z
lM0JfH/pFcfSyQp8G9MBlaN21GaGtlL8QahmLeb47/pNahtoHciNRrNmaFTMWT6ROuo8dWYafu8m
6WU+mygI7Q5GFvKyIWKvMytXvqz4VQSui15dH3inGP1DILndvG5fKZP1l8QgwbJap2K3GGcCYjnM
1Tk0JXI61aYghfs5I+G9AwlNM143V8QIpVyZjA5K4A86ITUOkBmlHtHd0m3o4+goT8e4X4J1GHTq
bE+gvYvtsZmG/A/ReAgB5lSJfqHRJGuAk2MSWTgaruIc8sdT+191Ltj2I3MKqFsXCSsWk0UwALmO
lLEGasFyh4Q8DHmRapKJwIY2a5a2ngOiIH07L8GqkAh1ZhtgyfKP04uCr8Mo0O0DvLmDgFCHx9eM
Bx9H6YlL+bv5yv1YZAGTNSGKTp32EJ79iGygCIhEciVXgg0TY3T9ZNfGIDO4HshI5mabHbDm9SLs
AwfB9Rk28bG0ylOjhneRsayLAAu+4vJvV7FQYu44JlEEL2dokReoFQiV0F9tNOxg/wFl4ca7m9TI
PDmw+Ij5GsYURHvJBb80N5PuHM0u0nim9LbufQyeF6fO3Nkq/aP1yabjqlPeVOYWCCEG7s/hIX18
yVZDgP/1v76X2NvE6vNkksmxNAHRWuEj3cgq299o4RJj7jfJUV7Nc661HQ6vXm+GW1gIyTgDVoLN
4xSzJ9n88LsLMAdlOpim46qIFiuXBDPyAJl4RJbDzYPNbu8X9x4c0HtSJmtVZkr00AxRdsyCpwft
2l6gTclBsFX5OAMWzGKRFwJeGlvF1sVVKclIijXfMgbPW66d+QrJI4JNzWUyZHMJc8GHpJyCKyc7
3CIHsgIMIHWgsZnh4Wj2Ua92gceyTDji1ebPOBK9ZwApgfnNxLDgiMFMtWq6D5tNOKYZKLflPg4B
/EUhPGFtcaOO6fGY9uFG9oasANw8QUobGqesQpOcP54CQgNj6bKkuJYclZUQG+93MBAaS1CPI60P
tN6xLJTaW7aPROdoGZWS+k1SKaYZkzUpvSTcIAMRcLd6t24t8N7g817rni/5FbMNrdNOYmPL4OC9
UQByAouJ5zwF8Y07MuZwey8eFb/99x57T1s+lhI7SOFFusiGSXvFPIwLUtDuYP3JAndMK95+uwoQ
g8g6TE4yKDvEC2YAFCVaWiOmsiFejh2/hTTe3vGXDgHTIStHVn4u3cR94OJlYBf6rBgmU6pqRkfV
sVbRYz6LXbBCrX9riXIyX4V2OayvC+4oE+IJnK8WAE94sjRNH9QFKCtaE1+B+tSq7Z06iZlhCncL
98uMjKY3Zp8XojU5U7UMKbzLZ+dRY7MvbKaamOWHbrv/VUNnLPKBDe7CjbEyQoZ08M9I7onIkFMI
96RTH5D4aWMXodiAkQ4fl4Fg/g6CiY+vzJbeCoK7xadVnht++tdcjO5lZteegeOntbABfcRnOjv7
pKe87OSicrlItH7+6/D/zxw+UayWOlt1tyKmWX8DS5gyTuQwObKqG5RiwNrCBRR2XDgJCzUCObu0
tEAcUKHphrapMTCJPux1KppiaXm1uMexXLJyNu0g15RqPX54ESvth/3gynA9OaCEF25CVywNMj7E
ufvnlU8loyNjecnYbR7dN8IUanOBZ3UGHHx6QVHQ2N6l75ht6ThzjApryL3fYbT2YfAllft8U8Uj
f2aa34pNUD3qaVoEyghllWOcnZSihD3yQPNvK/7RIy2mt4PJRVP7L2rYmZtQ9aCm/79a1VCqtcAY
CazBOBkaXUu911cUp94er6yfzJqzmq3JJk1BYkGSIfVeQQarMj3CVqV6tJ9RL4UBu4VOo8GkqdZG
m6q78mRHKg7nRkojIP3ZciYnu8ZlrOCbBihwpmzkHdLDaB95d1IPV7R67LTYrm80+uyr8/ZALcvc
4HYQMRkRd2HgLXBOYWYbZ6uO2OlP1HmDbe5IR0x/AZ9jlZx/8I8gLxYTev09pdCb3zx9XeGSt+ze
v9I5qEEOGAULxLZs303fm1cpxQDGVyKFYC0S9rXyoFnk+2QKbhtYPOzxdA5dBJ6Au4pXIJz27eSj
WimBl0dVAzhogvA12b9WBf8yjiOe4yU3h82R1S6RHojbGaHMfZydNJuweLztB9IBAhNJ7EfUlzlo
+A9/WsZtdOlYZf0nJUu5PdDFU3de0H9UShb7MO+Fdnds2QK1WdNPeY73vnvlAaxnX0c+1itdLN42
c5MK6qaV2EWJXGiepPELXQckhWhEziLcXDbwtCxsBRv3Yk55GrKyDDXPoYCk2mODfMYG9hU+Oo5A
6jR7qksrjK49UkoaHcmtLIqoy57BmiAwpI9BpClZPZ7Vjj7OO00yIU1THUtKNNIMFn0GWagsKm6c
I+zAs+UsSZoAltYFx7MBl7ZXcp4s4njvkdeOAalgfHcQGGqT4gBc6azgmLhbsuIROBtD0l5pI64H
vlRfhxJ3fKmcrxvGy47ABpUNlgKJQXY4D6oDr0+wniOV6crNnIT5cXsniOaAJlEjDxxgjBvksk+m
cntGYd6O71jnkI+4YaCC1Y23tT6NKA73+fI3odv8Z8JtLLRKCMVvbJgpxiMW8EHDLjk10eWcn8kQ
Y3SQR0S34ixwLj7PeGBs/5ErVBrBXHCSqfllxaZBotWiLukiWb5Pv7jrH4ByEK+PL++Lsudq6HG0
gNpFd2ZHxWypgudr08L7HTYpMicx1DYot6YfY14FQ3FVphe00ULpaBznVhqTnSDaO1sOeTO0dPEG
7B2+OyGnfNb1fL1lxXFF6W5VSPRnfgRiDUA2KwdTLulZhgmfdd7kROmbQY2fNq/OUOCUuAOJOp6O
P2wKHWOk4s9k3lbibhGm3CeC7uyATmMRs4lCkeunasGEzfE6TYm4wYy29BJsCSiOoLvXXv6Dd2uu
6pE7wPvAnqE6RfPj1QZgHWIXvuPrJ6ixr9Q8HcgIIVf5EBqlQTKa5pjrTEvGfGhHMA6N9tjFGBUm
3Dq+Np0tUp8otZhWHP3PGcsqE+rG1YpPDdpk6w2UHTIF65ZbWq6iXuLhUzbmp3gi2dTUMOCcwEkI
MRQ+h+my6qdhiKnJL3swlqXvubyw4AYFJJU4UWkb5xRAdm90SAZJ3e2ETNBE625xG84a0QbbkAXj
TKq21fjLa/ag3gBnQORsbDM+zt9D5ye6+Yp6C9+TdYINPW8uoFV6BX4NCA/njdh7Q8w2969Pf4Vl
pTphUvGatu6fwjCXfJaceCehFVcQBCMqdR1j2AEs0cdcG+aMVnJS1SbiBI93AB0NauMOYmzM9o4D
0DSpClguXF2s7WTUxMIbhCB59yCragHHxKi6Z4OCgNFMmmqUCFtodOtc16P0VJKKmPeotFXnFXr3
pkCaZ4/deRZlSUcoSdxNVuLcqqN5n++caCThVmZf8VYlRQW8W6qwXLfv86uyTlPKJfXwH0zPY0d1
lFuXllox2+qiURazctEj/dWQiXaAsT7Ylo8LQD0K+WQJ84pNeS09tMG7uk12xnh/EMYTWNEY/o1X
gNU+/spFpL9TnfhgPU7RJd1UqvSlq/qiSAo4l4cx2ioDLDVzEVs/31LEHbqsVSLL9Mhymyzc/rC+
EAJiOoO9ciabKvzkTZtGC4hkn8GeEbhDLcLduX7Q+CHCd90K3NsD/O+0L9I3lA/+y0kJP5xe5f7U
B8bWBMN/NdNUM88CGUu/+qe/iETxH4pXvFMyoB2AAgCm/Cr4JLH7Ay8cPi48qDsN17gqHm+BpATX
nvkRf6mqGVenyS+fbThUdF8kjqP0sCVQg3j6T6byDxiuvMyVJFthBDwM70SOJs/O6MNdTizdEZCX
AOXpAArEH2MJNwA3sEMhP6vMdzt50+p/EldkGDZGDbSkSvnltLWZzpqodgf6Ns1euFGht62dohTD
AOlnl8rTgwtdXonH/e75OYi011+CkzPcne3cpwm7d8WdD/HsqeyKJ9dnQd9onts8kDxd26+iofbj
pEOXJHxUsUfBOHOBQtqQO1qRipUL1Ft8acrgayJZR+HRHBJQSYO8X/wA9VjgKjWqDAq5KShTmekn
LVhkS+O4fogEHWeWVKI/PiGtgZTogT4+b0Fup0SN0KMJOnaw8dBwHDNotDHFXxZPrWD6pQiuD/xx
DUgTn/2fqQnV5XYQvKzLbCC1alE+qsIcYRqJlnn3J2ZTdLWpCDO0vxVcHxxtkEUUJCJ9NTvBDqOp
QnNqw1Tefc/i615enmWmxDgbR/z05JFJP75yhFXeHA7yOIFse8dHFk0vC4SWMQn3NZTpy7aRglKm
a6ZB5KAoq+50UfiwX8OLiqLynF/XsPQhM9Eu8KnQclzwNkokT7KKQPFqlzUm0aZ3fWLKkfgLsioM
uKeAH7kugYJRUOZtMMrrIWZc3CaTN+2Nit+Ir0cjv/K1AqrWFQyVYaBU45QhgnuqfdDj74V4e7oz
w4Q0h5+BwcpMZP0b4sanUM93D799gn8LIGD/QYjCWoGBNPWsSxEhSOR1jfq87D7Y9zgEtd7b6sAl
V0Bq/k4ib6gXDPO7PxUx/e5nUAcgGwwb3n0XMaPpZ2ZCzaBAIKUsOADiIsg8CPnJQB/MrEi1rsV9
PRf3oM3IBVgNGy+IOoQDsUslxsV0oU2SXbmI1lM+rj62DFP8aAR/xgeYGpdOEVwHOrOWRpBTAgSL
guHeBsjczJrjSuqA/YF7Y0DkEF+fnNAzcQCAZ7S8hWNB2+2Wu/8EpNvMX0pCnb7Qs6WWIlZOUD9u
a2KGOHf4CLp9N7qCb0b0Ltq3f+r1P3WAHMVTfPYWzfCRfryn57f/1C1aBw/e72VnbapgykC4hjXX
n4u7V0wjqgGJpWw5+zUkKT1L2A046s/Im2HgfFUVfD1pe0uecTr8ftHFSbNqjEN0g63Vw+LYDrWP
TlyVBlFSgwsWl6xoKjOai2rjwbEXc7WKxy9MlSpn8QskSgMTtP/vIPQ4ijBEi4rA/j4zwDA4xKm9
CNngvQD9Qc3wjVAkZ6cwcr8ll3YwkKURcq2cADUm2fWib6p+ntLWcoWdl3UNEQD9bGv3myvJAgam
nvQwZZFnjRzHsgflJ8NPZ/rO3oS1+C5ApEsA1SfXzia2Z/DaRK8ScmoymM23HH1pKbri5jAOtzQY
TPAocTV3AjznsSR7DABKk/Lw+b8SHOIJAi7JO05ysGouuWc4w7ofiPJ64iX5+hQIMjNohhMiTo5o
dv0SCsFXJhVxn6mQyoFcGq52sMgp48IXOfJnFU6HokExftSW+ic4qFzfRTLJl1XHBi1IOuA8iFOa
jfAVFrbxoXxi1261Vra+JpOulmX92xVFhuiWrMvKOfAme4ZqRwaaXtMT2RLiCYixhYepF7r0HiUO
pcPpN7VYo0GO1Drb0exRPKYsufhVb5ngXKHqc3JX4NzSwz1wiG6cjFO7JHkfy0qaoBGUQUXO/S+n
pPNysl54kIvhgW/BGLAM2OgYF0xG0SkUyXgk07aBEjKzXLh+M/L+li+wtXdUbfhhiJxOjA3QwHr1
H4lTUbdI4K1kYET6ZfQUeRPF72RF0MhMNfPKKY94OLZfRLgLl8qN8fBXtbSAxYUKbm89GzaqbHaa
6fB3Nu9cAm/6QgM/P5iGO6Z/7qp8Vt49etHl/cuZDzBnq1hSDtqhBs3XufVP9yqyMFAJh2DMB8Eq
fK7OkWkSBmdMG0CPp8vAcKwGktBNc8ueuGw666xgynjKnYPk12b9NLeh7mEtppwpU5ftdteF0rEV
sYa+JIKIUxM1P5o3h/ellTZQYGgJo48OoFNWVVvCHi8NkOrI7uzBmquxteSI0mYpH/ryR1e59U/j
0zfj4AhZjM8iJRjqtUPI6uC8esPt/FQkw1mk666bYyDk9Kh1gJbPISKxPUVCWvYMbxNvdvANR3Iq
n6KTu2BwbauapIa4+AINMYeJD8e3bfjka5nxzeY6NJ/rr9DHBbjiNrk5UJRKyRMCl5g+wMST3I9X
/aj27tAbgx/E9F66LSjaFTU3+Fr2Us1tCU+wDJASyEArQabbR6hy0DGX8S0Io+oiuaadexCF2TAm
lWBxMH2Wd0GFHEg+OePjdOZtvByRjhdZJlOiVO9EWyK/OqCKFGFrAdfN2s+OKnAW5BTDfsUVdhru
bsPhS81N8NSdSMvD/eyfNU5VE6+SAIbRfJA6NIj4rfMMgQKFnBFkEpSyEUT5dVgOkwqdrZM0IxrY
T8295HUsidpr3Nh/G/oOkfREx1XEYMHaxPweEt1ppTIYeUZA7BOZp2G2+i80wUZ/d6fZi5j2xTo7
pNYrAZu4BEUBrEqFhC7IUjlpCzffUqbjlq7f4WL3l+d1hlfS84EVbOsxQLVKVTmHwPHXcBHmnQ9v
3zFi9EJbatvG53P9u2cFei10CdrSXybxpk7WvanTG/V/8Hs+y6a9uDqaB9tSAU/juRkDWkEFiOG/
Ii7ubU8XgTYQXq/3mm+0KESQi6rQX2d5Fs61tSsusgEf75M1AkgXt1Y/J9sF5v64CJdHfQQWQptp
fggRFYTXJ7DL9c/AqxshqqRelQpJoAiEuGI7eYNVJugDAQAe46b0NyHKTx5kNbJWi2qcFeK9sgX6
G+DJ/xVjwZa00fee/c1qqiIdzMNIA0bXYnSKm4Ay6RJ74Kr021x53PkSTyPa4EoItzxgTmz3UOVs
mDgCnejg4CzKTTqDxJeb7JCDZWL2bxz/RHToNVZyPwLtbEqNlrDNOKhtXJZwliR5NEuujKAI4OCY
KVHQNqMVRyxrPvMu1PnE8XStQW19xe4m50FjMLjPNh2Aib/H0wENnWzDD1M5mpyiFjMUv0q6BztA
ozl64EiyPoWwnxFA3DO7srhq6l/735olt8mrfASCvVXMc64U3FwBYE0JM6PQz6qvvPSWqcQ+F+dU
mDAWAHGGq/kn7ghZqX41kTqWpUD+7bhwk6QgPoGgQTFsuzgc3G+BVQZR0qPUtkuIBIXYuhsxhG71
ysFBZQL0RWi/SCzHHw66IABFGR77beDfC0inDTNCnJI+opx4kq6Wsjr+BCMTdihZF+vwnCvu6ZQN
KFcs4x40D4ZQarNKhrC9Liq2v00mUSDOCwu4kvc5IwAr8FZnqRfpGvJ51cy5sln28AsfYgev2SCW
C7OPZOsVyv7aQ1GS3Kian7wiZFDHiuICbtGrWMu7NxPk0URysZRyp6AU44BsKeI51FCWfP0qqo28
Q3+ayizNu/L3KkI9cxj+ZTPReocuMH1QmLstrKPWazxLNysl7/Mz9hvGwHxEp1wB6p23JdFQ2XqU
RA90t+OvqxwKJqnsMrFUKQ+mztWcfsrM/aEu+611ZlbaycOjSPKSi0RnkCeqZ9ynXPWhK8eKIQWA
76D/VNLVaQOU/J5L5hqtkw8h2QXwOJ3lVDWRjOpSwTsSaSMh1IgXJheOODIvUX9OatExSayCcdN2
+OFAX0G4Xm53ik5VTuEQmhGiqmNE1OQbxDPUnJpmnnjMG3ThjaQNahOECS0JrAGjjYWK/gsmvZnM
CbLgveUlukeaSiqfIEU7Zs4GFi0UmfzTXEL2xabmDn78emWpD/4iLwjwaQPTeH4OEoVvqoKMzJXE
pCUXMcxs8yGoZZEOjEcY5q0z1k1UkMtaD4AWdurHcV2wjOUixvIR/kZrho7aHYTx2t+XqFxdfMWN
Q+/QU/WV9j/Fxh9C/tcdEh6ume3Uj3T5emQSqTKTYsN28xTK7vRn2BsgDIxme3/RD5+3+RvkSwLz
dTQBfy9U+BD/BjkFHUC84bShnEAGvxyB05XG9j6r4Ubp4PPqhzuiIcAO4IXgsKzZuetZdfgzDQ+B
7/bg1UtHDOfagB6SM8SGBrclLFqjlwca1HiVWW6E04wPFR/SNcxPrH/czNBkZlG7GX56HK6DLMks
uXbmcpkOYCj/Iwryctrf2LwvZXzIzESi+Ak+c89ejrZSNzke8SvoBpiuFysDQ9JqdtRCr4jveFlT
lON0KgNoRMUJyno1jgH0QMUEJppXHGk2u2MZBitWFtV/LKiK+FqwU4Jx/xOiYcLCqukiWDFdYb8c
Jk+i3msj8Gfk3tYzPerDcEbdoiACGY2uhrGHeb0FsBoZuUZ5Gs3wbcSoGSjatJHVA5RgSFBor8tj
F9Cjbl4U6+l3uG0iS3c048NsyTvDC7SOwSq8rXAnlE/CU997+qAeSEQiHkKS0PyZqpoDEGKGb2AM
iy731H6cH3gHOwBbKLXctZzIo43INbvtv1vw7vwp48EOSH94WJ7HlcYRwSMBZvnSqVlqHdxeEQlc
I5oPh97Pt/i/JkrtAyXIr4usitC9ube9Hb1g79V++cEU/AfHKEvBGL3Me4rjCM2lJkfLn10/ElM7
BbjqR5UmzUgng0TNXlFHJwdfitir7GOnqV+qAeX6LF9Hl0D751sUdOAVPbyGZvoGLIaVG+H+7jsp
EG1m7IIo/D8ecncfgpJvk0TyBL6buJQ6099Xb7tU0qXjIpDwSmeaPYa4JgSM+vR4sa01HeE7A74e
UIAwZvmJUO0nJpztnCdWfxHjf6jNTLqBE/wqpc4fIgFFB7NkmPsiw7CjE12v9Xucst23mRbM/sbv
e8/dwGE38P/ozRi1h3bmIrhg9JCV0+7RUusfwh720pfgV1Rkzeomf0zX9ZIkQVs2nF0D8Drn8WJC
n15bhRdSQy7TVwUikL1o037OEpfGljG9MGC0H0G9RZJpmOhCrdyWVsGJiZgibomPb5h1LM6BQILT
sQGZ4JWTIAeF9mFozCTE/1IrCXBSj++nlsRu9BHxUse+ZM9CENP2I1/w8AHjhCn43nCuDgIFAFdM
9NGqhMPJ0C/ZOmDRg8e7WULvVWCNkSlX8hNLbFV/UT9puuY1mfvuLLkUuZAt60lQW7QJDCxGk23O
aNkrYXj8SSnE6hnxSrHMBe//8S3hknTPzP1+1B3OkoLu61ZBm+Uw+ofYJvQONNwO1L14t6d4p4rP
WKc/EZoySRB8yPkrYbQwsTAp2vyOXv3RhPpz5yA01KqjQhaZqheL45pze6aMuZ+uqPn87kNSgGQM
ntqVwTsTtk+kPsn9CMZ++60VgaUho6Y5tgHFZTps5DDnpvuREjwIi3DC8lmCeJ8lDmzjG4brGnGb
E1FvZ6F+voUESSws4jhVKUBQhBwOIYjO1YlSLUGQ3ZTq7j+yN/0E1EnoniKQnAWpLAN+YE5EMoX6
ZByLA5fSCbdG0eRAmkevE6FJLGsUd/3IBurURM0PEK39xsGcoz/+cE375ODOTN9dBbYcESqThJtu
oN8c6XzzR79LDk1LXBW3/Jrc5Tyz+wfbxu713R9qP7jBzhz2Nfw2tccE4ErxlRVzseJ5OXHetZQQ
dcJaaeDDQCZEreNY1SULIZWubS8/NhB6MmRAhG532qoNfPMb4YjQIkxnOFJ5PYP3FIpO0eve4Flq
mg+gIWEvoknPfZAWDzjhJM6JGdgvTLt1koQ/6Usoek4f9Ap/uhUL8AJ1leVs3TDPxMPOy3FJSsee
xnudOE/TCfou1JylmkrFp71VZMNaQAlXPO7WFGRkbGcxJfeMf9vKPaQKuWqs6NUkapuT3ZjB2Qfj
qIhvAj3Ma9TZ3nigedMjvC5jSB5XKJnPYh4pwUbcK4VLdBTBEHlcaCsBrAv+TyyBYdU+YZyeQifP
QKQ7XxFqWtst66cvPo+EZ7wNhrtcnRGES0VyCrCMlOrTrkwWdsuvmDvrhnbHHLKy1GfYcNvhkrj1
ul6uviI/M2aXl+xfV9dX0mL6E1t8Q4Un6m87gzbccrjrGX9pp5dNHp0YOImPB5n/FPsN1HtU3aCg
YCiQFilegYo2C656/zBFciB3D2hH1BkEOXcSXVJV26CJhsvCwMU2Sl6bTPL5lJG+5ridpCXjUTxg
2NpGn49J+ySZJgrnVmgiXh1ty8CB0et1L4qcWCFzQtgnEpdJvWwEMN5ZBpMTcbqB32T6HPT2U7U2
J0ug4iiKTFHsOErlWMeVMaQp+InU22NwUxckoZcAUOa4c84yJZEjE0B0krgy6zhOy/+aqohHX6S4
MfDuUXXgKMNvBffyd1SQK13M4XNo7pA58/4EKGmqFQirSTfNk/GPhlkhlBDuMX5GipGrU3ylo+jb
+urmyXUmlQ8vK0AxfhujyeUcmNYyduVdhivIaqp9H2yaGWfM1NK1LXX7md4QGYQFETwgh+oauG6V
1y4bVJQHhqYHWh15t/aOSOv/kFqaeAUzJzD06ODtMfag8LBujI8yRO0GUDRWixCZRQfl2qa582dg
YFNOU6/2tmWw//0U9ZDfgsw5W3Q0Br2QLo9Qi+sbeAYVKf+VeU+EP+Fi0KWTEsZxfB6HLzqSvuAQ
of+aZ8pFvDrGvzWVjGeuMMglaKLc4tjIAUrcdr4sSlkt4FUOFgxCJUXDHFpVWBYptuTbXNK2Oz8a
ILcAgez+YET7w0p+q6f+lVSYvWzO8E5v8MYDG6AFfcV8Zn9LgXejPsFRL1cVojPfk7ZM5Qf2DKI4
06LtctO+OJ2giga3U/LVOkLY8/Wkf9ZE3ctzAJQcZ0ybIOfy50dlM6hMmfLRo4nmy83la3LWEMHg
iduFRd2GeN7sOMqP8Bkb6oQhEa7eMIZ4ctPQpv33hgMiFuwXgYxZLGj57vPVVZgOZogNMITyJLVQ
NdAzYS8HrcXKCSD41KT+4CJyxzkuI+ZG5AuThdiUA+9z32JEx/B4XRSWMRcfUZIYJDpVpkEWlcNj
ELMNnbngzoSG4ihh5SP85ciBQooLQx2FFY7b+VJqke/hdHoJn5f1YDqCVtfd+BKlfk/WblEZtT4M
ksa3FK2FJbjToDeYJaWczN42j5sTOpShmmupeUcWP0+SNH5ZEWFhIX1FpGfKc1ZBr0ShSwv9mo5v
kJqOWNC0YOVS1o2K+mLI2edNZFx/sxV8R8kDNadBrZ3Vej9jVABm1RUSBlr8T+V+BU9PkulgOclc
5r2LUcEohh60e7qV+e8znO8c8k1PZuGc6DRZ1q3IBOFuONDdBGS9RPPMj964P2FaQCMjhGW5+MLF
0xy0Swu69SfmnbKjc4lWamnWbs3J6lOWE7Ua6HWRRYUqlo17gBRUv9zPaoDogkLNIPNopjSXPJF9
7n+oCREaZnC71UEvZ6h6g0PhTYF7O2OjgzDBSZ6Nn0rkYKmyyxP7iwu+n6XThJVpwO0EN1jwMC56
EjnZqhjLhy/xJBJz+zHyOa40xayzgGa2AhRB5mfCsfxdeMuzsdattvg5KpQ7e7szXDa04bdCb9WN
mHqkAl8782h4MBe6OICHFuwe6duKCb8a7mns6pKz2vO95zszWQugx9g5nlmObtKrfN8WD7kXzGPZ
bksTJhPEA06u3ySFzWZzICtfsjI2QcmrOLxZo7mIrbInckldOTmDspQP8Rw9o3QoWX+PQUiFJA/Y
PB515MUCXqZktf5CJehrSM/tkBYMP37qhib5FrSFxNDyUvqnvKhaLLjs92gTf43PJY2CZQOynT8q
UsobmxWkad6LxEqRBgSRabCbCytEIPxcRTGd9qiFZOnLMb3r1vBPUFPa63sI1cNdZhmrS4TgGYWQ
3BI4HrT4lLgKpn18WELQ9mr4EU4umIyTbiyPlKqbGmwdP/nbO2f5/wFWswMsNzIzYF6/8qUoohrI
LC/vQpkFNNR6lAKjJaMcqmcQpsHiuJIBBJH22KlTQn7KuO9IBjnjRyKTbIGB11Lev7WTUZcPcj+t
fWeaEl4yILc9lHooHBruErmIa/BcpikarOiD4SErMKSOsioV8TkP0WhhA7a3Z9HblDDTnZeGBXxB
ul5CWCgS5uBXkmB7ic2OuMr5rIbiUpLh31ggnYBy2eeHF01ZcCY+BIPm1ZQDBNsiOXNaCgB3aOuZ
oCcJkehPmTmZGpuEk+XMglLpN4z9lFMXl22TXfZg0F0rKmB5BMVgVC/g01OnKOs/lx25FoLjRXun
2cLWAm7SUTXRo5k5rXZhg5a/lMIT1c2HeYIzV6WooluARRxQRgNy5m4cFUPA4W9Cul29PUpRMw3s
HvIqWHw9ntg3dsfTLeOuYeOcSz3GT2Y3iVlJiEl9xQ/IO15jWxqK1kfSkbJ4AhF6uK5xc2se1+gx
9exR5qRaGmJRUK65h2/98687j3KXyYXOiXECH2IvC3dIxzIb9TuhlkvkwpX17GSQd1zfsLWA+WzD
UWf9aHqezLRYqhVYSMQpdcstKsOA0ZJx+l862XHgqVV8lo/ZyLbFJb2SNJGV1dJC3urGAFuwUe3u
Lx5Hme6rJe5Wbu8oVyJ/BF5R/gZU8/bK0sBP9UoG84HJZWdz/1iIfbOX4EpG7+PtY6bs8ReY56ql
uageRIlTnmIyVaN+pVw2Qidk90w+522YIAfJpbsE7KYWWcgEa4OFzHeGIi0GtufvVgIpjD7ArpXC
yxnJwaTy0j3Mrxsb5nLzkLJ7Dryr2g/Av2+KUERtEtUl6pmNFNJba+aTsWGNYVDV85fbl8DMJPQ9
mCrFFI4fCLMWnuKRjLOedtyn69UHuiaT+3eGH5Rdwc2ipw9SC2w2VXnCa38QJun9uH3w379SFHqk
JvixUr3KR9QppdSTzIQEQrMK8Xyq4dH24PcYle8pMd/0/qn3U78tyl6gAV2nGV1c2hXEQR2w/ezG
fg0stCg7pS1a1SyEJ5Gc03V3Z1VqHNBhkVUP/W6UkVplWhmQTDB9XZd9sSnI4W2JO8TJ5hN0G9oj
yiw5wT16w0FfjIcP+itBcZ3ZqCX4JdLHa+TRU6Fcs2dYvASYTkx0A7PJoAYe9ri/dr97yZ2jRZNC
vLAHq24COSRUPWa3spnjSVwGrZOa81dTMHFyrfKTVNoxRPliXCXkgY9TT4ydIp1Lqsp4d4dFq+4T
ckUsgwLjY120tdBtm/aK4A9CJOWAXPw79HS7ptdHNVfzWLYNlNi5apU6ok4mLR/poQvbuefSfUpn
seZe6+Zz3OkfbCqirKN430ewBsZOq2/Qpv0d70uTCcfDczS70iDvCZgieKS6nuM+/CwoT0vRjqDr
T4UkEDb5IQ4JQHza0+3DukFNtG4az5Y6EmGeDtS4MwJ12b1d7Pa7p7Ehz4lQMbaR+aT9qdztORDG
TCqYTIcvlkScz/R6vYCLy6y9SqqgiLWt2uvdtS6RyTf0Kx3fv7vrZuHabLeT771vhW+vumDQfOhT
YfXwi4G3BD6NIyLk72v4AJ5Ynh5jsWI2Ymhum+Q0pXSYiJ/qySZKVlFQEH3Js3rjs9YAvJ5Kj7+d
zOwV2gCK0421JN61QypMwK7cOjeAnpS5Hz3vkinehK/E86S2xSehKO8spacsAg5TljPohWhpJNRU
QEgsJ4Dyj/1BkwmqXVSbap0nWkRafL81shuZaUtXzm9KpIhnjBrNJDYPK1vO456nqK5x4nsTxt8v
63g/zwZp9/hizYu4j42JjrDLvqKvRng2x4yjBf9SoepR2tv1abUvBzSRH4Cp2zG0lyELE3ttCJOb
6AOMsB9ap78P6S/gG7LvcfB34TjrMITYYIjN4gzHT7AgZLuSaM4KHlY9Swr50IvdhMRnJSwqRQZf
+68ksZGUlzgmWVtadFR6zKs940LdRC27YEs7oSUizfqTZj3bFZNJEEpdLz/HRFJgeEa4iPgL7gqX
KyAOGxzY0EO9YAFngVqinrgGDrlf20iwu+u5JakBGRJk0dQGJqpEBlLME9O22/w/fm1t+dr/7QWv
U4E6YtZY7Pb3wKCtt01byNUOa8qjGyiYLoxbYux0/XzLDUWA4NSSES7w2nE3Izl15gTp6sqW514I
rZEXQQiIAvrpN620hiWGX7tsxcuYv4/EUHZtiTb4YTVVhb2mtSOBMHXZi8NcHAQsI4S9KdufbJ1f
nAf9LezQIqaL1dJM0MMb5d+RRhXHe2ymXfAMNjLu0Io2L5vihBITqkFLzkJ2rurHF2WPrGU51x7+
SHMT8RyZ0iaZOHixzsWFi7BD+nz9yPN3bqNiFZpycH8tB6G/4R9Fp7bpmUpr2FYoqq2e7wqPnBUn
VV+2tSsi8TstuTqE+W6nWPr7sE29bMwFkj9R6sdqHBgjMYz+rKG7QP/Rr0RIq/c03F9LDSKfrK63
Aih8g6sN6nWRgHWJP4mT1QUlM3kt2PFA39RRtawx4G87oN3XGxwsNOzXIVN30KQTUI5j84Dag8kV
nbDyAUjU4UsGegWEvRPOEEYLaACBUuPiUH4nFZdC4Oay+Trz9VvbawLSHazYyJxWVOuhxewu90Ri
p2v1DuJDqAXkWsLvX1tif13GtfrIqAEdDbqXi43ZkU+kftqQWYrlzkow0SK3USwt6Wiun0m2zW0C
rHq25nDuWpV/Gr1RYcuwNXqdcUn/H7LrHWIXNs2d/Ss/gycO+KFlfvpULs47ZC7xWzTBn/x3Q9+n
yiC1FisSw0vYIS1GlqMeqYSkYnIJCrO6F10XQwgjYYCKZLWco4S26fMxx1k3ECbmsAnWWxY9bicO
PPlJt+4hFXVSTWjZKEjNUHQzRqrB28VNk0RnmaJ0iBN/++8rfSPD4++wd7+o9QGaxz7p74rlTllh
KprdIQxxiDB+vBDRVb+C4/uLnMvdQ+8M1F2stR7tw6MwojQZ9fbkMxnZtvFTY86HHBknOSGcWzBt
zVDwajCTgA9h6PVvY8/yiCjZnqPrJs4fa33w35JFaIze+8Ka5X6aZWNyPRxsteRHTxuE10mIj1Qy
hBmVRT/xfoOoAJmBDygkHrg/J25RI2Y9Ig3cOqb9bWsjv/wqwhWI5kGw+cR+sXKj5JYmM8ySowjh
PSJ9RenuSznjcKmwL2UW8lcy3Su+5c/FUessIja6i+AtxVZkZofMojc5S/wJ5mC/Sf9bioYl1YAw
xfX3OJ7y1F07OdM6LDxN/wMxK8F15idSC4/wxsIGcOkrlP2VjR1mbJ3fPBRwKbO13UK1VKw+Sn5K
Fc3xAPERrlJuMeszKNyw7Ym5w62uPk7hxoaCsTqOxQIYoVgUEkZ7JcTgQ4PYtOjW+OYT7nMUi++y
l+zm5jIROAq8t9pvFR+oZvCm91jw+ndVrVTyRKCsN4jnmEqXO9bhbRvS7EtTXu5uG2ZuQ8TysiaV
nF6GDMJKLsOqDuqmd1cuKxkiVAl+gT53CDKxMpOQhKxtTHtCI6eZR17URzz7NmF5Qfd6EaejthSy
1d9J6P64Q+vbmbc0+a0NxBeERhktIJHBzWE/lTWvvBGwEp8snLOahw76XunvHZTVrYyz31gxrN0W
BNr9UMJOu2Nr+4CfpYRUa8GZ/yHg3sr+b/7DjhWJRHNQv9gCvVHLBSTj0eMstF6iwwxZBux/5u4G
ryzZPNSuuDH+KaDzD/Q6lB2teBHJDDO0MEdirhpQAtcezd8fRFI77R0ClPJQTrtnfTzw7HvTye+s
dFbFjlY8pjgAbfCHYRAyzvpixX2cNwc6VLrc2OQWiwQBAw01C7EDAcHZyZf8LFST3UON1XXR9HUy
4tvTUgK2AghCjA7J6606BO30LMQ+mYXxkECFXVrnVT/zoig3q3xtPoWC/8FcLHO7t296WSM9F19W
wwEfAgi84zCZ9R3qF29NBav8vxECFcdaKVkFh0a4nnOtndSxchY2m9g6/NLMTxwpunZIVRrkrXjR
EN1sFsZaLpuS0/LBD+Ls2vv6+YbnnBFG8KJvk3j6zmYXgq23MAnfYksg7WoevD+/CKnpMgX8yFxa
eIsBOnx6//T+ZW+bsqvantWLqwCc4SlkTpd7x8H48yMZtvbZp0XgK43cJnciWLKYxte9vI8Mi6RR
QoyqAvSqy00msc5d6v5q6mlQcVGotykY5j9dcVyrACB8JVFenKzJQeTE8a9V7PfFaMbGQB4izh1I
ya5FPOfbBqhqI793YF3YR3dqFd7scm3FpEnl4o0itJn5OFs1unm4MwPqcQLwbpmFhXb3z7AWFjV8
UG0EDmcVWPChUZ2U/3eRqW/hhNtDN69iz9gC1C5Q6R5DW+OIaGBL5ryeA5jNR8bBmxSkcwUZxJj+
Mc/yxv985EYViTcwcHUbdEVAyGj+BwxSUMuX0OCy+AOulSoHANsceuVuLjHhNxT4vGQiCyQT07wY
fbdRJrUpK+5WoY5jyoX3Q7EKDplm/VpFSR9AM8Q1Cf8lvOqhn3iswElGfjdaf7+qDGiX915YR0Ub
W4gFUhsGSuoV3FDzQty+mUHAJGMlpoShjhUCXYrKX4K2L/F1qfX7rpjV6iP6m6K1rJw0GbAp9xQz
XMR/5Vz5tJ4mr+0I02lsH11foo/2W5VvBs4siRwdLdOwwoIffdaS6dcIaX3e3+/nbnwjDD3q2G4P
Twz4OPWCWsH6Nhu1KhPGx6d+/uAhhxFEok83cjMjOuIitFZgDtzKjtGhVx9iz3hB+sy5qEOyljkb
bHKlt4empjpcUEe7OClmTGKnrzGXgcR33P9MB3vt2+wZ4q3CQCigP0lUADzJXGltjFylljbONjLg
HpGRl+MJqIl9LjtF4KpGZjHqIJBJDhZvLC+vFJNdqy56aAANk2/T+bB0eQEf1g1QtUDfuv1O8ewh
oli0mTUD2Fs+TOFLb1KAuGCxTxZ1TNxv9F6unh+K8MEk36eprtWIRnAb16wrW9O6N6nqpabbT4Vs
EfRCJ2b9aPwd1p7lFy4W8q8oAfFqXsLpNV1SKZ8uWi9Ikzfmyt9y1xse68sNo225CqiLiFaMmIR3
zCIS9K5VMb8KP4Uu2vdsB8ElqfMHC5DcTgyO8CseHYE1l9+sJoDXgFQvYPVST3hRAXak3SGZnLFG
k2jKvKZ9UW4GmdHiZrTmxaCwtbkdVHcGCm9hrPWkTvyjm9J2rZ3Q0WyD8v+nZlIVLESnPbU0YOtS
i6GZXa9QsIk16jMEAdk3N/1V9/R74WZcAJg44rgs/8DMpppwKiu0oBGu2HC5EzpmGArAJWEJUfgl
sO/2vhWMmruf3WaTGg6aI1PXoSvPJn3/ZJBBSEZPMwFXvubCJ7XXOZgwdoNCFfva/yEkVMigblxM
VaEifXbmq34u7Y36yD4YKg5d1u5RBmKh7KYDUAbOpcaynrtz+2lBJooVZS3obhmUkM6CejtbbKST
Yq+aFlmamBjj2pXZby+6MXqlVKe8AgCtq4923BbGbXIL+mm8MU9fPNvQ6EbG9jdxOA1Knmlf7T75
RnfqJVqNu/67neYkCvz9H6OlIiRmQ2Zd8V6pnhnLaqwHWGBXosjEaD0HbtZk/XBcfQWsArKxuQJm
nSDmyE7F+Gk0Mt5cYtZ391g3Yh9CVuCVCBeD0yOpRvOsQfrPHwvlAyQ7WzrUJWTCLaF+Wqaty2YA
oPI9GtxSGGSx9x+bxv9GYU4Dzax+aff1FVwpJS2csWx/Kb+FdZpFHeVgqgpR6JdIOobgtCajBKce
QS9iJx2lZZZLp4clcVht+izTr3iW431mG0WgalYar02eNSNnL8mJLPcx5iwgE4AviPajCe8+/SJN
PBdm1C0rLzL8c3L3CIwOkLisCwfJxRZCkV12xAjhsBmqXEcFX3c5JeXtoaAn1/x55+upJ+ABD+mj
u0orIjzGrVtV9SmXL+xuGo+Brm8+M0BJKbnPJ9D3YlabxKuxOXU48RpnNCdKUexEXRFr156+HOp7
tisN2LC8z11V5TMBMlSH2UluFdQncYWmzxwbfNUBf7upZj4/V7PbYIDXdD36OqLu2oSXKpU3J0Fq
sxdzh1ppkjh4Q+h6narW5KotLzfm5dU/Qc7BEoBPBuiyRw1n/Ik8ZR514gaI8YJq0qvaq/c3Xah6
35b55fyvY5EBSzJjNkqemAd7vk9L/UC7ONiuetnhzyrBWWtFzmXS0uKLfgJxxMTClgYKpaQEI9Tk
kM4qPkYGoQeez2xMvY589IeX6OdMAqMtqYhT3hk7urKHnB3XpnESAaWRZqtVcU/3mkbj3IyA/7j5
0WZ3B9MwB/V7r8mZdpT1o7f0KTKQ8RSoVv3Sc24EpGAvbXvdpk3asoNQyoznJVZoHkr8cYqrfuJt
QXh1AH/lAJU5yhNwS2y6stYRMOYeAHLOpV7DpKf5jGe9xAk9Iz0PqV454CuYxR2FBpwtwhDt5Frj
i7NiUTosF5mJeWUYzPkERCwHtjxBQ0a2uiqcgvH5oH3Dd5iXMoyD0HNZLsSWyIcMriS2jgCxvqX+
RY7HzgT5/GvMcT2iPVJvT/HB0WyQGOCq/sFBvlvqsbNlqovfmuW3otVu5YMMMUAIs8EbQmGA0DMk
8GPW4Y2gK+EvBSHoDa3l1P2Fs6x6NebbfXm6KEtTs5KRjvuEkayOuDuroQDayn6YbEy8AyAqfDER
/sxraf2hiUOM0NcJD9tkBD4WQuNOnxS6OEnnXPMB3IwVw1PqB5kNFkwfqbDvzQIzOT5s7Dc59F5O
AN8yf97JxaBs11p7DmYsFpsQ1MeuZXkRvS+Md3OZsOzIc/oL2d37QYp4BPJt5qqN2nUXxmNs/RIa
yN1SrHpmE+Ymk2FEPJcP/zwJOFtywowQKM7vaMbCxYBgBPFm7dHUA1eus9CwmjFjA1yhWwMNYUhK
I3iO1D6m7SpznJiPoSGPT+CTpm1yzyFX7RM4nWgPhcrwPnTxpgzO5XixuSDcAmpyus+dRQAc7daj
wIGhzsFcVzyFf1OluUSuuqdgSbPBYnpy7xhkTNZSXRPAfkwBN5w6/BM6VJg7gzuMUJ5r7CqTtnHj
0uGyMzdT0BI5cXUIJD2mJ6FfBpmS8i/4lIkvWibaAhXZEADs99Q04s6FBALOXm4qINn/+8hHtwq5
zMUQTf2sGgnORU3cwM7Eh3N8mHqvWOBLrYmyaFL17gVwoKkdmOfLndNv30qqgDT6ExACqTGowF3k
Oyhtfer4EXl1RcbFpmEYqedscoiOHBeq1ttaUOWUFwO5WwXHreVBxdmVNzD9SA7n2L9z0fydYnP+
nmDXGORJE9kKLyI8zbxK10r9SViF+f85/h3uSbVotkw/0Ewl4V0FiOK9p6jZPlXfqW3o05rVZ0vi
4p2Y6XRVt/tgJg/V32bxAuVWMbaJ3qds2gkSyLneJ3PYQmDh0vYwgx9apSeaFhdfr3lOwCQUi0hG
9+8nJaxTRiQ1TmnI+cRXHINmTOWaoSRF3Oc38eSa4kNVN1rJ9Vji7rGkgpLjyPNieyub5Sl8EeOq
Z0VuwFH6qNT88uyhA+RqKAYtUNaaNzZt83u5/cE3u38A9dD2sW5Bkvy+JkdGw5VUbKZDUBGnpa/+
hdjUUVHkxSNL4XC3xQpdj7BdqBCSqZfqG+RWAmYm5MhP4MT2FqM5H7q9NxJHHgGHPX+XXR+E9fD2
WSbXlpiMmr2oXbwLYGBuaGeg8Ze3FaMeYIae3qzOrM86JVgCMCv3B6XVPhEqtZ7tRzzUp08NE7YT
mTC+9MPioToMI46ZqlmfUlof/IXcNzRdbQ8NRobFECJODGxKR3wnW1pnzcV0rsJYDf81Ngkaaga5
bXUUTYH+vuARlAwjQDoOjKS+PpTF4MeP9Ab/moaqJZsOQdbYHXBKKBsFQaZJbJz35g0+AT13Q+j1
ZiD2wXGJGJIp5wW3KIox+WT6t6eJT+yLfuTw5d+tUvqLFQkoAXZFuovv0KQnmpBK1A1sHNSasQCp
1f9nigWBGHRHcZHf5Olo2t+WGSfw9SfNnHNaZ2pe+MtRD9hn0yO26WXAjUtHSrtMEJr++fATG9zH
c6dM4sSug+5X5kEmhl5at70xT2TVsPqldmaAPRABtljw4wh4aeKHx8KQyuChujrh5tA4z+AFnDu5
rb20JYsjKn3T8NJgx6Y5h/5+Oy4Uj5F0IP2HxX+SUDqqcDN8mUeOz2DFf4bZahizBq+kUEfX5f8h
Y3GdHYF+fZuQGwNFx+kwTmyDRnPFdapYt7BLBoBTcmcJ6q2CLcX3PZUmsoIqLU5EziyhdJNnRsdS
GsgQIKamnOxMik788RtXga8OAE4m5y9zC5pYNyJC6wr3pTvqDc2kZsZmYsXCBsqtLGxa7XHrizP3
oJ2rd54zPMVBMAPuU0HOWXie3fIL2mP689nhDDs61gZHKmSFnNQNORX2Kzwm03rKYyP3gK3ZbZyK
06lsAayNm0l4Q5JuJ8VIskE+RD8AAAYXfzUzm7AKgIiya+/mqxitlcgfvFylwpEtjQW75jNmEvDU
LT1IPmcompBkCCx2y+kPmTYtpK4xqtkuapPAdTQuuHpEZTus65vJtFUqnGmwj6WcBRxGSP7EBP7Q
7jC3zaXlbowVqEK2XOnqwnBEGpXIb34yJdbA75uKy18dv+hbfYMaG4JixwtW+kTaINsUxCKMO5xs
zCpIHFWT3PU78qhtrhhP2bMMFrY/Jy9beZerZ4eLX4xrbREqfK2KEdy9UFQshgn2vT0xcVWsGVQX
/1GI6WR0hDrbGgIlK4P217AN/nJesGRPb8N+PLCSgtnlbAPyydtJMoHbhrq2im/V/bY0Uc4ifyU3
C2Xrq4FXh+0EfY6qmtrFGYOXhQTosLsQZ9SFUXJN8raC4cYtl94Kh+j8wpm8JttkFs0+9j8KPgeM
3W2zfupFECKkFRn0W/jYSFi+bUyxH0sgbQoIMDwLu38tPySpggNw24HnuGRHPTWeYtJJKGq92RYS
gmHADmRz8M/zgVZUHoBXR9NnsaHlxUGpC/HpgNfFbAaIAW+W6VznJrIQZFoaM1WTc52ZTOQma04l
30tKy9Yg/IyDD2OM5kHap1LND6dymXfCHxaVZv3K2y8+WY8UclFIL8iCv7upEGxwtSik7QsOaKqm
VY2E3Xa7ykRZW26FAH4JPyNwvDWeXvqsDjauCEf9055jb3j3ghr6FxORV66fM3/Po5GY/NMmVg+J
/v4VPKElHTLr61q+mdmujtRol85+x1BZjuuhchRVdiOwv0p0KvZfSJxP6vhcdxJVDqAVVqLu6yfG
E+Bn4Y0dZfg1uGbK7lvKiZegI/hrCShqQiHesMDSgIoFTQXcVGa7+AUYzDgB8A8g1farnY85azCo
y/Wfv9PSFzJKcovL2qmeROdBEGh3+fK597h9feZp37wP+i4THNHUqYkRbAD9a19pDwJXYYF8gduw
KjeBOrcdUBN9fExc/rGLElO0y6vfCpEXCTHsWe1oQ1PVL0ch/x5Jr1WHMohKSwHj7D/ODa2BgY+k
GIqnI8YamIoghTp2nMad83XXNbXGD2PIlWcspxLJjQKTcvNsrxaOH1yDqPYvIli1tzVUAIeZEU/5
WgpjtGn4kuGty1iLdFYCa2Mkce8GugWJVeCvkkmIFAfHyd/N6aeEGxeoL0KFoBki9VoaSMTsg5MS
0kc4CiSocOlRKj83B7zk4Pl/u+5unzSF3QRtWci/dADJPdwYRJByFJIuVIBUAFyTFi4bUmYD2ZvE
ayEC6vglS5qUQCQb7fiPlaiTgR3ldxibSM/LrlcULETku5zDvbr9M47lGDe5GasMOPPMZc1YWY8p
9BkNIveZbioo6vYrDxiZ6tylQSoJv1yhEAwRPjumaZceLjQgpE82y+QUgg42nLK4LgU//HbyYDYP
mkUW2gJYAucVe8eBWbbSzPM5tN7R+QeQB3xXqSfhND7K/6oz7TFbbDKmZbazM/Gxx6+AFjb0vYZp
lH3eg1cCnCHO0MoD4+oCSDuuaOwXdlj10NwR8H5OLgfui5nQxuy4KTi3zRmNitBfF/UrXFyEOyjr
PZAaneSWVMLq2n6zZn2LknE097NbGLSOvjFr+fd+GYsuowpZiYa5krURcZPpJCYdK1K5W8j1tNuP
6tOtVB5YAHwcT3DJkQvGCg15Pjvdyj1zlrgXKeWWZLGUrp7aw4wXeAU9Leqb2FraU73j8P+AzqLW
fxgb2izpbbNiMKxl2stXZFruerEfDamn5SK94jX8owmkDGbjErvsxtuNUoP8di7RFTWqPlnIQsPq
+UH8bZl/tfSiAtLYDdHb7JKUuVkyBUu5to1EjF5NViWBuToAlxbTPanQB1RQU7ryUZzdBFJe35s2
C/wXZDxUyZi5++Oh1KA2eDujPSOzYBFE2fYx/Wrvoo4g2FOeO7BZyF5WZVAnqUPMcU4wTcpvLZMS
ltFghoJ81i0oL7CWcXJiHdijGw644iQmkwFGfGUwX4E2/RVgMn1LXd/TcraaB5X14xNoqiDpoiCO
jvLIxALz/R4b3qGlxG/OxN8S7D17PoDI3enwW3jQGhvSdu7pZL1a8y9wlVDBtCWzoNWCNpFyyVdE
wLlFwzsafaBIM95q5GTtLMtjHN7AhMSt26Y/znfQ7Qak4wUVPuav9k2Y7HeJ24g+oS2Ott1DtwQo
BntWr4a9OMnBW/Sglq2Y36q4xzDlTfmjYPkGhgxCgzt5eOm/ozMrK00tpkgvS2BnDmFa1maKosj2
d0OT/1trp721RM5dNr9qlhgkpbRrNOiYgwIzEQXhnybeph4rwmPjRh8Zynmfc6lazkFbOFnwL6Ht
wwRTgmPUEYbCiAO+jwxWqRI5m3/WrP1L7cvUJG9kcVFfu5zRT0QZH6yJHrIp0MM3z5G5hij+C5xS
b5aK3P+To1fnP7+oGRbWPVrhRAmlQO2G3nqk6kji5vdDuieZ8OZMiYOjgLnSRuehSYFP7KLgIjn2
FRmaoaUFzxnRK7Nvi6M3Mc79XKBOXtrtk11r1OJnmVjZ8WqU+8LjupVa7v/YL0WRIb9tlxe7YbAt
T6w9vO+OWlpFIhJJa5gojbLbzEN1PrhSg92wyHZk9jyTx2z3zdDplIY2ud7UO1WRwEAEC0oSAEoj
XmpN96vyT5JrFbfjoT0yl0OQvqFf0B6sSNBqUVsNGSodDpmUvB3Upy0E6SgOK5tOkKDRN+srjZcV
4HvlJJkHRVsDoWa70WRvuHJ2PxTwd45C4aD9c6/zF022TyBw7YMQSxvcy7KaFvtlEl2rf8z2Wpno
+vXyyrpQeR1Ltg/6+uiTh0syzbFmHYbYqk6s3zpyOH/P3A20dgIoxvCADZpRZrnGBwMc7646Gl88
EckDindr9SqO6nalD9fBTfxapp7jMTQSSRmrL7tsj+CApVqdornFfl31trqM4flbrLSK8o903Cbc
oMVnHKR3ybNnFF56bZgupT4dGUq+0ZcUvac/0LLc4R0bdMy9sLvOCRhDGQCCef+EVfbQnKIOVLrR
WsuwmuuUbbyIJUmdNNghLOnF3GLSVTsWJYM3V+u0UCaKRYWKIf2vGxHXAKWOBs7kEhzMygk0dHH3
mjv8D5uy+EyRc3u/naQ7GgeeBjZV/f522EBpma/Tkmi84RB0XaKAtKUS5JmLDnO2qF5UjiY312kc
yZENtpNkSurOncqoyXMtLWGhSmRsDDqkEA1z7zpRJ5Phq6lH7qgo7ArXFkkiXhxgTbeaQvlqd1Cm
Wcy/V/REU/PQn8y7GouumQKgmC1jv8g00UsndOhWDR82rFYCIIC2boeKPEsrhEiB6C1BEganh8Ky
2SjR3fcV9xzVQ1c84O1AnNDHmHVWHZldTGDUJ07QNZIUfb6A3tu4eGBFrCm8cj4L/ustjC1XiXyH
kc9LTgPznrwZgs1wXxXipZfWOcZBVPtw56AyrsDRG2KeEIwG3g3j4MGFCgDi6RHPj4n62ltV1WYt
WZ75DvX9tNeba6oPIWkf8ntDUQcKqZF34DmOkDKlxbeq/Xgm21B4Rvcp3GMmtMmUaypHf0A1FGpt
xuBig96Q2VJO1U6TSQXoXCDHXHMt1ep3NVow3wNhztAOE15sw3MAWcEH4xRMS3Rtkujxo1p9Yeij
WaLiLioYVvtbg5LeP5qmwq9qw8mTjgGSuW351SzUN4GTdo2EjxqdvCYgGrf+afUZ1DbLW7w1Xp/B
Ox4Tq5nDc+iZIZXFz5e1AvnxvSARDPQi3SIqwIKbpmfiRFhZyv1H4TEBYUp+bH0PyNMK0p0Wphj6
q+3P89ZasfzocilLM2bKzhWV7ThkxNUAj0P/JmZVLhdvX/SmuGczqEGOclaGuLdRusO47XZgPiF4
qZRn+Tt4hD4nhiZA/ATKvnbWUGIRNgA6K1z2JqGx5aCb7HBvHi4dIPemMa6Y/V376ocelWiJmVl4
r1VVVPNkC4g2r1GoOkSGjgjBz3JCdup1oSDpjTxrWVEVQOHAHU1xv2rq8VAA6IKsyhmYihXI4xtp
zMndIPYoAalnBk8ht6R4FjGWry0WI8XTGnjEfIE/4BQyNOkynFATldZOJVubjBkbhj6SJvHwIE+G
zll9H9OAwaz/wLJymuqqSwSO43HnzNiAocgEtLgTrSB6PvP0roqL9pIm4dpzoxY322cP+6Pq+l10
14ktoinaEP34TNCyHGersyOKPZTrkcdzSDsCxuIDbxH7HKGkvmX5hWyuCgvBu6kf9CvL2D4+ZkRN
IAGqt0dlJ5uHnJukqp67Er+MBprPgAyl/WY2XsQzbcI1uimOdB9eByWK+hfbpN3hztuFASKiY1QJ
g4VuNehtx8Fd+E6dCP0U++PbCKeps7s4EIMMjQbFUZwkjGKrm2ESvHkzFMpWBWghX7FunkDSriZZ
ocFnuYnKA4a0fHMuHal1AuetzZQXid5mbI+mTN+UyppmBYHcYZpexB2M85nwbnUxvVDsvnSuZsvH
DYJ33o5RXo8VRsUepl8gu2E9fb68c3Iu8PFJMw/+esgjI7TR4UuPlwc383eKppoBoijpivchP8Jv
7z14HkTsSHIFQELMHEKAZounsJv/omOP3qTO7MXs6v/RHVvslkNUGKTgdbNxcywJ8RZtiM7Vku2r
aCRvEQ6dxXbSMgRw0UGvH8wMaEK85Nl2dSG2DM1oHoLQF0imexv2zf2Ej5Sfx/mKnQnbjjOppmqm
OtCfs+xelRmsuWCExd+Y06ZuLdgImDynar0KpCSA9gkTaDdA+NCCTjmbFbrvz/7e/SA2LoSyd8pg
px7322UIp0kGflIJRl0Rl0z6RTAj2PG7JxrB+2HAPt2QMqIiWEXW+6b3WWA/qrSQi8eFzgivv1Me
FHmZYFtASapwcXUo2hUjDiHD8b8GT/pC3dT6OJYkxcRBrU6uJz3JxLSyfBhY2eLOB7gsYNsIE8tp
JSEPZ1ev9MyP/6SPu2XDFXd2og85vgaEFkar9nc7fzgjRZOcQS7ikbbEp/NmT54zCcKVfBno0KXs
nOz2oBKp4RiR+t4xDBJ2wfIp99WPyZ4yN4t/UoBfGhPcnsBQpxuj+l1AdR+ts3D9dCxqhVNMBGew
T3Zues6nRdRp8UViY3DH8mlWabb1YFIfbWXxuB+0yGQKFFOF/e8TC+xuDvCtgPU2VJT9+GmxVLD7
022dzb+OatsglkuRQiQDpZ5i63umxJQqlcPNr5IFECr2huuKIF5COURBdF26ktVCmXAYIPq9aujv
Fd1TjMsnvEb83iOcZ5mdS9UrLgjY2AnOEKUGmjjHUm72uHQWY1LfUtVELBf+FHPfYRVVwuGb6Ipz
W26dZgPLvK8EJjzqLyP2tJ740e+oVAKzq93Dm//8gCkKxUesahs7xhFQZVEP6UGXL6FeR3fA7EcR
8vFxIQW4qRpcqtnNYxNGDtqG2XSIylx7NccPVocf4y0kdnjjIvaeDGqeieq0FVt4L0emzhHe3nxQ
ATgIyleo4n9zxWTyagimNb3iKbSMSeg98rSucagJpyibTxn02QViVNO6Bh5luUpmSHa8//KlgDmn
CS3kV2MQoLzx0mt5s6cvxNATHRlep6WXIuR4jgeQq0BEEbkzDGPuhFkH5KJn7tBIG2oE7G1AIbBC
PeqUFVEaaAuU2xm1bSD5aC0GNlPF7+hDvOFQdibzzST+25LLm3/nPsnqNanq+EYduWrNGdPYOXEB
moMBxwD+uWcESHDyVHf9rKf8r13sZoUJ/AazJysf1b5CYUK8ykakg3hohoZsOwp0LVVZWX09N+8M
ELQzasl3g7xHrcCv5rk1Uj3q4kjHZSBUKMyG+XxqAIggupOHZEcVSzeuj3L4m/5AxhG0sEp6WrU7
tGOBo43Fep/ZEhPsxRJ064voKLqWcGvat2ustktqmrJf/UjGJ+0XDPvIgvyF6Rxr2U6HdIQPr2Gv
dgS37puD5W97RQylMGRz7AShm/RXoTMMTTjSYzopuZwQ1Ot6L4p3Yqecsg7UqOS1KxRqV51Ty7v0
rO+e261fF1eECbk9i4yKGS0h+7khj01ptVuGG1PMWvAwfXqIL3phCkNaKhPLjLJrt6mckMP4R6m3
aA/sOWTpGxlABGyNaW6rv6Jeve/NpVd56h3pjblT1/gO8oVR6Z67xp07KIqnfAfRlUGqqaDtzdEi
I92kOB/b17554V9IYbP1fCpslKk/XzoNP6nMs1lToPzjdZOMl3kAigxUoKURzqSZoTHyAJuXxfCc
WJe0JlMhp0J4sSi5HnPvvfreiYDM94gr5874Nrom6+I+Aa+Y7rWTU2+qUo5puTYVCbnsz1cY8fsl
kouipYiNoDl3gQDlGjqmlY761Dc/nMVE75lW5tx+4dRqoYh0TVv9tkMRbY6SCu95REPUc1xZu519
VDjA+/cvNr+wVe8IiJsgJoY0K1p9nBsDlUeKwBTa2Rg0+/fiXpEPcFeEN+pKo+otfC8oK8VtJ1JT
/ECNWUc4lhEnrfVs6hjKKZB4uSBYUSbMcNROinTIn0B8XYrTCBUyumQCSPEM3tbYUWLlXRxyQyPx
8G6vgmMTCbXGom/TKQKI1sIOzGealRaJl1C0ddOKHUFpnVosoqD2c/2iwRktg1jF/FIODpZ5iP/p
siKX6XbVeZyPJZxyIJoNdXE7aKziASR3kDbTejlgOMaCiwwNct7dON8Bo/P+pG5BgQjyy1ij/qje
XA869h1hXdnTZN52oFlfKtJSh/1ZPYeRsop5r4yqxJ5GmNDyACR+8VfKSLVQ7Y/ZEyzfF15xDNzM
RB502BHGADvfjKIclSRChNuNwezHj+gOjqGAkAtwquMZYttrO4sb4vguyQpp74p+8A7vi3hsix8Q
1edRD/75+FdGdwRbGEX04buNOojX5HruiAoeZWbwreVIBemsFCSIc8x0eP7B6r9j47Cco+s1oTvp
TZ5aHIf5EfIYFx01somvzIlDr/BlpNRiSj3VXEq/xgEKsSVo9Wm2LAFy38DV4nyv4yTLdGF3KKX+
jM/gjIiLlDAuLABDLFLmKextXRnQF8S4BOFIY6lfYNIruzYAh1p+WhPYEYlOi3WA+d6+nU00QDHc
cRzIgEFJ4N3edvAVP5WwUj8ocoFvbfjdOjCIR9og2EiyVjsoOiCC+ZgS+CZfyeh96nh5jSmqqXD6
TH6r9mwve1EmpxpDXzr9Ce3YeO3PbQ0TevpBmmqmhblOcWnrSznqARZeZJRJNso2SrxXgX3ViDon
GhY0+k6IVCHkciewPhiJDzBW+GaFtq5fWYtWnBX4VpVE52dXSIVG1unBjyPix1FKO+pYaTe3ogaD
3S7o3aZtnLCSMg3fxRysotRV54fKYYbregJspo/F6k/uAF+LtXiA2uLpY6ENbjKQUbcRQrCTTPhD
b+krcBkkxxrRxTSDRMukfxqHxFAvAp4QhAZm7LnrrLaDcJsDrSvK5c9W6XeOZkm0BK3qZ1/JRH6c
KqEw01UIEQnEXopfDPxssSbFBrtAoaQMVg2KCu4Qse58yhc60kMkWXL1SmU122u/ZnDPaBGeXLMZ
GJeeY2xhcWvvs4C23IGOAfMtbETsOy6vMx0VHJ7cFzmqKaMlSpNqYbbVESzNJfwX+lPkcAw+ktKt
FOOFnE+39tdOD1dZnvrIiqF0vqjttkyE4opzz4zQUlG+9ixWzgYfRKEZZqoLdkfjosUrqi+GI65o
WDqGmdo8eno8r0cMqSeqh/YKG/27E7zuO0LWqOym3uegNthpZdvS5nxODFIL5yJl2Oj1hXwGWJWy
FeUu07JKiQWzOtHm/ZVbr9Foy94cnXL4lEHtobkLiufX1fS2hzlItwp2xFsHc9N5s7gJTW/Y1bky
kmUjvQMnQwI38chJnYx0kum8SkwKkxILq6qqraIJmpfKON3ngqARLPLdybIpbJJbg4zdd2p2lT6a
7f8UTleyqP7Ftnh3IF0ADKLSLAkdDRJwdw/0k49kMNQ5s4GAe6oLwZ6tZyWUlxKataxD/JkRd92w
rQLcSWU05acpFE6p98/8lVtN+Ugb9BE8TqdSatZ8yR131MPP0ppsK63/pztmueEQUmt+ixso0g+q
18Bdiwxk4meOY3t11duRUAGtksWafqEnClQJ3D41ouvsmHIxR8wwe10D+Kgn66P64DMV8UJX93Q5
dXi3nZ7LYEyuGsFKpd/i/R3OZmWCRr6dWD5AvOAaqgjiDwbMr0Uhb1yji4q/HAksZ1nz3Isk5Hep
/kg1ckRjPLYkzTsBqb5fu2qcAVkWi8hFm9G8EzyH1crBj7v8J4tGWODIxpY+MayE3Ahqk1arS6Kp
OkkNBnp1UHtuQH1ReGxarNaIGInshLEL7WQ6q06APwp7wmaksgqbcKUYKy1GiQcDc9Q/QR1JoIyt
VYymnKmVzUSxoqw8IT8203jDtBmUOJgufVR2egCl2/zK3Mu3V2YRlSKJ5ISQhgG4MQLTl42/12nD
94NW7hV9ucdINb3YrXcX40fD3wo20VtjhEQmTksL720+eV+2pKSzcC3Ohhh58KoD7udwEi5O78EA
6qpXM/A8xvYOxci8tM6NP6/ugTiKfP/BpI4zbXhuykd7rNwGFHXs/Ks+zNi+JFJEYTvAe+5YQpdF
nL9qcnrwNsuXN0S3TW7fXRzBQ8EHFf5N/sMxwv0QPuGRLALSALv1ZaNGLhvhfsmlmGmfuSglY7w+
59rYScevdHdTLi1Kbmvn+rTKxVEb7ACGqJRLGLg0/D81fQrAgWu3JWn0i0bojirYm1uWrpjMQCJF
OL7+QLWkJ30RMMg08yM8n8sOdU+I8i8QNQewwZwMPZ7xmRZdnq3mX8jttes9mdQ8QqBp9x/1PTUF
Jqi3VgpqGdsUq2Zt3PULjzkvSov54eyQz5pzStYZZ2l0ntw8hv87O2H3APT6cmTy9NVIQtyVMDoV
gyP4Q/TzzJO8OuvILTwyhytDOXkirjIL1NB6T05FdKnw1fFxUfSthaZ9il41/M+y02bIqIvxQwX3
VHUBzTh0yZfcdElwacKKmlOpao0PEIMIPZteAcdzNLWrpngGih/bf9sdaSWWdudMZjfMDCcAu1l+
Y2GyEq6QTl/rk6Oq5trs6xBA3naKCow8Q3Aai1DcY5y10WLdLmixtKz4NxnhhMljMIL3TrCYcKJD
L0CEBWs7K+xKo9oNndPPt5UHjT4gmrodUCu1I16qTiP8yFl8C6xY64fjENLIPi5MNbg/sazBB0n2
bd3EK0RyzmotWL54Gald25/Pm+OVz0WzTIUbmC2wHOZF60BFiZifqHQjpjdVf7yATbaIyvh0mTUA
U71u0TunRNeFhfv3SiFLssP2VzTp2iDgMk2OzpcMpk8NHOmMDLH78ImfEAbDB2IXbMyqP1oIjbfO
5BW+SJFGhCJ2UNVj5edNzptTaX9idfo0ngWJStsJGYQ3ZCpLMSXIkF4f9HDsb3O6g8RNjYoARsrb
dKMbFLMT8lzgICtgkhBSLzW587rnXVDsuQ7FZ0XmDg8tcWQPQAkImdBi7Ni7kCJ4qGMk9LBmbnBL
EF4R7UKnDs9Wpx9AAs9ZXv34I4+cLWTQM7QsyOKWEZqLBVq+mf+XrLkzHaXrIVFXcQBFn4dqIChb
FCwZxZzwqBzN7uYEkhuvzrxNf6lI3JSIo+YK0wgWbxCrMvTNYbuJfSVtujXMxtjVWDMC+H2dE4lw
dweZi7yYZtJZS84zx5yKNgK/9rANfFJU4nAuiWXCjmAOSzM7NNxFdrdBEDhh97DFNJVIzAHSP+Ar
jAOGMglsS631ncEZ0YTwyf8mQtvtww3C4JQHpbrDFFH5RmeNoZ7L4mUZtDrJYdOh2pbYKEhVAXsi
Z+3emgUzPUPiy4La2sm0OD5OtvuNEz6Pi4hhqeQXpM79HMlOhf7r5gUtvSZFJFVZhLRNfRoubdjz
1t6CSyz5Ixh9mXOvJ4aq9v+U4AX1I8cuDef+/R2NHNFShmIYbgolozJLPv8/uk6vVg5IasrTsqP2
yLgQUJriX6TxKt2JkxnPpbPJlBxEyUiLE2aX2IpRuo8DStp9hi+dCqKx07XW9aIJ9sP1SCo0rhFD
4KIftJQdOsySAu7EW6zPJ3XkEQDgJ8kWnol78T++MClJ86GO2LdLN8Vxd7+NCrxKU0Euqgf6Z7Ox
XGuHW8YUxy9woP81xcbbKbZkv44Ic1axRH7hA4Eq/R5AQevJk5hHEm8pc/8BcKu0K6M4T3OX9m/t
4BHbqYnrwk8KZiTTZ4poy6cyx9pKKq+He0D/TFV8M5s7OOhl9wV3lFJ4AS889cLGb64tMFLgaBi7
1xxD8n8nuf2GANKcoS+TXMtKfeo8oAFsZk6s0yCXtCCCf5ycY3khye4Z8qV6yIKd2k2k/imjjnB0
4d4jHCC2v8gdCsabqAKfhHO4Gr1BcbO3GasC5wItPXXmvnV8nj3REAZQ1waylhK0K00//PcVZgp0
UmQSJO5iqPeB84Sb2Q6Vf7zSiFyExjVXeuakaZWLt+qh4v6lR0+k8dOnWWl5qaiRdzE+oe7bEhb+
PANQqpn3CXyYDFsQDA57M/f8idHMJt2qwpCN+sBKtM2GfN1MaVyaqzrvfBBGuicod+MiJv05Rv5H
3sNx1GYNW1U2D1xpeLxq8CjPeUSF8ni3M2ZsDgssEPGroqSaheKwxTDeWP0CQNm5a25IVbIWJOvH
GjToGqC1OJyXnLDdeIyNuEfIbUGrpxKKZsiB9vbio+3Tp6OmTLTUjRsMqtnyS/9uHSmqW8TOlUii
wP7QjDpI9cMzGcx5bm/KAw4y6dEmD3x5F2AOeH6nG/LJozcfTj1wX12buQIBJIy5LvyugHcAlaq6
6P32CTRCvrbRqk+eVVYl6UxZvvIRqwnmFZ7g8tjm0W705cvpwfP2A3gM1a+2IcN2pVPGB/8311uw
gIrN2/S7e29IVthPDbNbD4k4XgrQCbYN5TbgD/FWvf6yluypOopybwIoQvMy5Y3OrfAR4uZV77fo
132H4i8jknONAcGEAw6DsJWdSpJTcZbG1/q5Fa66dUlLSoGdbrLB1PfVy2DNK5n8JWHi8W+7ZuSI
Uo0pb31g/iDkJ1AMXAc9cW0dO3erieQQxmWwYpGE8T9ZVLUA7KkneHQheKP5m/HkSNUHiZYX4s4t
Q+i5jDe//lgpZvVo1RtaA1yYhaWJ9XWMXBOGtkOOG3BlE5bRE0bwelLnj1NRAN2lwGk8ppHhiekH
FFxocqO2cke0n+/1OoVzczNV305WaXMDdU4e6zkaHNebM/qRKaBuZHinD127zHNn8N5tfP2BRG/j
qTaVu5fDkuFudtbvaIJmyDU1R3xQH9ZRX0/6TddWZbW9nC41Ndf0XvFhz2VeG1tbigCgrHtohNDe
8sTUwx1lWtpld8fcupkCCJ9WEPXQyjjpRGnsLIFUiSv9XxY7MvlXAkHaX9JZyGKgq+xi5t9SP0Ec
USZF69pjTZQHRfadq4EYnEriP3UeE3ukKQeSeqJ9bPw44y2h0kiGg6GeLkojsQpckSCzZM9n3w1N
KIb9XZjCfvXBZoFi3u33M+S41upJean+Bm5+MCr3oYA97/vl46gERf3Mjt/edeCAbRhBNWbwvS8b
WXEwuIc/v1SFi9uu/RK1b2O0fxo5RXU/7JuFxAz/gfnQ7HTI+sE5eoiv4MCXQzReLcMwd2jFHKQB
lFlRJH/6MOLeFgiSdw07ydteCU/l0EcWONdEWj/3xKcnxWK0jbOCx6GvT6IwppQO28ONuRzI3fP3
gfIT4eSIA1RU6GCeBw9zM+RL4gKnB1H5vu5cvPT0J2vkcydL6aaRppb6MrgmlTxNRGKxJFSDQZt7
KEN40D/nE930i76HFjux52j8m8zz6K8qe1j/7MGSCuPj5a+VCm/f8ooXQ58RUKNK3BMbsR6T+MJ2
zQ3BXGJgjFLrjSiWc2WLf36ufdP/6rpyw/8UmsVWVSxwtyHi4UsiwL8ZaPLw7TtYbqa2v3G76yme
L3oENp0MZQybrO6PBk6u5d++FTpPwHlfJJfb1wGhmg9XHcHYEofb8M8zm3KurJkRJ+UROL6gCq83
28H62aA5hcK8pTPN+g3qPlF/Ym+GWfVvcxmz1/CGXJaZXJhgFlesdCcBiA4pYgcHM4Qq46zVkaLl
zsrA1aTDC0nmbTehTNaYwGH9zKYVrS/+Ee8AfFRvKGlxp+jquufzSY3MW3kjoWPDXtXRwU7jOMSz
0HAF0+caofAtu//qcT5+3/DL2BcQoNGIrH6Uz33c2zgNNzxM74qC4gCgIeMTBfefvriYpqjocOQN
BpEJIJ2nzl5HH95fYED/dqvaY9M2ubhUfg1LnSnQvb3Y0E8rwazI0UdavD5Z73RT7qw+6JnoEgnx
v81MdwK+nIOrxF3fggxSb/dCyrLL2FfPYXvzhrSxbrt4KFWOONiSoZCIsb9wKbV5O/y/wMuLVZ7Y
12j9/4DUGzzvMT+ktt6b/py1n601G8N7A0SoWnwPqT2hgL43qLd+ygMPVYoOPUqppOKGeqFrRee5
TOpQvWnmTOwRH1ywMyWlZUIuYO2YjJx5areRFvPtcVQ+LX9jLesjuZgn8XxzjzJcLkOSYgClhXJM
HK6FbHWHfNdxq3ZeeqCIHD8cXanMEAJjsT9lEiU5fFM90zEzOP2IuqxoK73haq01ykaiwef9zFZG
9/KK64EikkAv3vKHRx29rPJaMV1CbXlBkltsAgaMXbaJLfcsAHL6EIQWUR+TQzZkVfLaOFU1JexO
neUBJVbFwxdzNyDSrVTZHeiSJMIRlkLPzmkStnT/swHQGr+t2oy5KbmXIV65vChgvPLAD3Uidn2d
Y0YVd61VlY09f/n5wuSW5/SHnFQIWfLtZ/InW6OQ3a62aUToo2/rABVRVJwJ7nraasun7LbmpN4K
Qp6ijI8AjOQx0i7FCt3f37ALxusEV3nW/nJPOlTaJvVhNVXGkbhVDJf1qONXs7JIYr2VC8Z00Tc8
n1ZRdJ4WJ0wGR7SZtudoec0EPlTNnB2JwICO+7f6rCzh5XTZ7rsavFjiTP44z2y1dKUHUSZBQrRP
aYJlkBGk/o1SyijA4X9i0ql60LHKyAC3kwVogOaAOwGCtyxXEXN9b73qLQ+QPzQKhejf8Zc91Yr4
uIRFqsWjlGxp4UVNI1sbRvdKSlZAFlbdGy5+YOwTm5DcBjKoiA3bB2Z7OWIRh00979tmc5JH0Bf9
nYdRt4AJxmNNNP+RoaZ/5PsaBElBbfPnk38cgR0UZk1ilqaZW84WTeYM28PU0dql5sNLLA7xxUUe
kM9iLS9V4EHmTQZDtPNlemDQ5y14RyWQ95wGA9zY3Lfize6/5oBsxTu9NtFYiXXT+WDCkjynTiom
WZ5/STaZwHKV5X1wYAOkqcfQckrDtc7BY4jd5q90S6qD6cazIBZRmLMRWocTqT/DeGmWAyLZsGwK
GTbpD+nrm4dnEf9PhDKjbNkPt/QrikRxJTWG+GX7KNaCMWYzBh78GdVHFWM1ZJ0S2+4k1oXJknxi
KHRi82sc7hfFRTzPHCIcd9RVCwoVUrnTY4EwD9ZLeKxca8MQHjZ0YiPRqf5RH8lqsV7KTd5qdG/u
ZpzNq9Z9CxNfFTRbMi98hFOZrYwG1BU7qPSIIt3nFbsgZQ/D6OZwXKc/dLgbcrRZ3HAypMESChSO
sJBA96/mQ2+Qu+bgsMDq4+EQelNqtepIqn3MA7Fa0JCeTd4fhwLvYBs/xw6Zlu/ANcVgikIvYScx
DKO7lq8t9mpdjkMu/M6g9GdZFg5QoigVf1Vv/kpxuT6vga+ZchtKilaB0xaazob745xOR70DqHGO
YPIw9C3HjikIOMsU0o9LY+uz9k7G+ErCfjk6OjLv6qxxXjoxdOqgOrWg03Ycft3aD8HNHeROqF6t
aOYO4bBXO3YGCVjZKCsiVfI5lNuodPcG3M4lrX5tOimUObeNwjGibELsgpDbVDqoKPJgacetcnA1
VuDqcptvkRZOuisvD++4b3JUSioA/acZ6qOu6mHKEa+ZB7uuvJT4gn0BPxT4cMSKrCFtB/2suTVw
qATUnh7X16Gps7qVZuGW1y+Hm0sQUuPQUuu6a6gQs8Ti60wvGJIAFTlSPh5e4PlgwevNTkTeaD8B
XYrG9CkRW90aWAVXn+u3EU2PePkxgA1GCW0F052H/KXhLlkY50A28X8sfTRYXSeXzMW/vJgH7TcI
c27iHEilJQaS4AHikg9AFLJ1S39C/u4cG3ZhoOUZKjQI0EHSxzMqW1oRXY3hY2MCtiwvkN89Oxv1
5Kxe3vYkLCokBaY1Fu4dT0bqRT3z9t42NGOtT3h5LPcASywanT3pXvb+CbBGjA9vO6F7YsC3IpWW
oMju4EywG5apugEgOYTbE7dKzqveI31AoaWHxpmprv08QnIfgeFT5cen+nHtN10OjaHwcYyERPNQ
ihqCKXUe6vQS3/ve4CLnGbCAkevCaQKRwbQw8H5dXcI5VJ5JNbduQtTCsKdMu5i38/bD8hq3Wnki
5ZzDo2QkO3QZ7WGwlqUX1DBUkFiJ9+nKXoyd152jnbgPVtLpgQ4hQ7hr8p7DnA7eMSb3HB3UQs+U
QllJNksdlgDXrfkyjdqhO5sZ5CyWcwreOI35cqO1EQiKz2VyyjY06BnupCKOO3AopNVRB21lEvii
G8Rph6SqyB9ErU9Oz7CxvBiGU7fo79bEQYwcaFXYKSWKvjSwLp7SaqXdA31AVUbY304Y6ur+7Gpx
A1AmWNbI1J5ZcaHo23Hd4oq7Lqpgy3hPjesXZ7utDey7L5iBZBtztpowWg9OMGMkvq/wop1EzYDZ
2H8O6kA3PkewbIPRMENZwg247muNxic2erL/ZPmUmn4+E+rA7qE3xqlmLqqolvM4c8GDk9fe6odB
2qm2EgeReuOYLYCsrGoZeKD8kpys4IAhSfALCJj0zMNLSDKvOzbfixeiL1+qyapFGhI+aYbAQ628
zL1dMTAHhar+FcoUi1XlnomMdin6tdApOv/sbMtbBbCTCFaXxBlnD+y0+u4GzClTu7dUxZ4zqIu/
usCsUyjYPaR5NOM89Ejsip697kba6gqSei+Zfo6wMNd66clZdNW+ZjlEa/P2EV9UpjN5KSKyyHv+
IeNKW4cubMr53MplGaPUOS0B7uj2fP67DRkv0gdRl6dx8LkrfvBKkz13H3TFiTH4il0JEChwdXtX
A6EGNl56llt5CNBUpJ0GvUU1ogbsyLlPxikXfJd/4rmG0bi8JjRgleZHooEgk/jjpSAjJjRolqu0
cQ7AWQ7nrp6fa5tUSF8OD6VFVwbG7J5fpkqy6k11bNw6iDRQUkiv6YWAs4nVscovucrHEEWvdMMB
10ST1CEWFd31E1ajl5yhiQhgKAyDO4sQ61QOPQhwLUpcAFxWL2oIBNxik082Bsnb2Wt9zu2C0eXH
ftJpDCNCF3zj7XpF3LKK/MxGET1K7/Jc1YQsfsmeU0YUNkfo1QOIqqij3L041b/Xv2Y+OCaARzK0
5hn/HL53GqMmOuH29gHfaY9EzzMzE226bXG9xervOGwpqEH/l0lL6kTEP80LOyfTkt5sX8omCWWu
OxHJ6Bn0u6frFMKPl7nFGBCk0KilRMNfbj6VgS3+VHgAI+wQyB4POh6vUau1tBdRF0Py8nScR9R3
Ax23KVxb8TBqi+3cmYmx4sEqXcwnUqXfLRbZd4lddMXegu0ZWsg8nTb8BTuSSKK7fsHHHvW0lPNT
UJnO0zBFCW1MuB/dbcHp53i8MUipjXVx22uus764G3YXBJiaM4jSfhmPc3sVQnQQ/6dgM9ro16d4
oHm36QgayTYwL657CXwqZwjh3S4Y59PV2mfYFw5HjZLicZpru1ZF3pOtvX1YfwGpXDXrx4CL3Bt8
9hAdArvkXNoorU2VE7XWbT9KTtN7fyVhLaA0uWgTYQ79jOgcZsjS55XFEC9JGs2gEs05FBC5w7Sa
KhGlN2KRHKNcQlYSR3ApNjRc8PNtL7fGm2d6WbqdhRmSOKLc7RYGHbSj9o1Rrs4jDgr3F9qZZQDQ
/DoaDfTDanDdOEZ5JnQ18Uf7iQEB1e6lG8RRiOtJfqYKat9G7Rj0NVcIi9SiVtrGsDV0qkOe/47Z
KydPqJbf0eKCJ4hEDRj4sIDvCtCu7/SLI7TuLf4RGw+BxWii/riF/tqZHMMM+K0PTGjVJXw7f9u8
aRhXM7NcE9cwwzoXqna7ZTWot/ax8Mu1GQCDbdNwltqcHyDKf2EZqGdXgygsyZvkNIuHm07O7oQx
0weKNrUUePqo7IaAsfqXFB1IS3DW/6xQyElsFBAfmi9IhUU6vqy2JNlEvQ9RA0ehjCMao9RvMvWx
xigVYESCiDsos0Tth3q5f7H2CMXzpYpmj+bKwlbezcu/+vJKonU8hwd5xKALdN705CX8GP5Bqsty
5/xlEswlESBGaEKIX00bzD8R8CmX7NRBK4F1VMBXunYpG18i1T9dhy91koKJGHNlywp30sLYVGce
r/pUXWNsNBihaL4Wz7gHxdSC5mb5/WeM1hgMANXtZeGONmXRHtxHt4x0sZUJ5P1zj1TVvIbyLMcG
G6pDdP1xWGjxXxvpHmbObxXLmdmFDW6e+xhHozlfhdEdoJ/TELI7VaOv5tjzDoWsJpujZ3ESMIV3
v+DHxdAritXgneqljkZXiykMr2uoENv2O2SrenouvUgALSNv6zDp8Hwct/3CrbhILZSKqZdjdlT8
Prkf3l/O5mi92YwTI8dKE2i7k/r1sxIhat45J9pVqfpKo3xZVuYgQvPeb26zD3Q+3RUaC7yGVWn8
8FB7hKJE9FG5nawisnltEj0k4Htb7BPiiP28R+pAryot/tQt5rA75Z4VQR7mvuGeGahtsphOzO32
rnb5y5dZXaWRTe7t05IE0R6ggQJv//wz5+hH17UlNWYGzLKce1PrTgerFVP0lvSBkpz5K9hIloA2
Ox0FOoCcaGL9ABcDkQ6os2tlgzrQXTI+OViT1nwYdToePiHORjq6p0Zvcsqyn0FCghmLQj1aR70s
5vbdper2m5HnTsv5jx3kXiwFIWnDm0EtYy8Uv6O6Iyq+QmBTJlsHV/uW/uzhZ+iKRNo5vCrIN3vP
1P0HvtUf8TnArbkPBumftlDufiXf6CCqTYaDZKYh5FnetypdPqn2tY4vhdhnsOnk76Xo58dU2QaH
lS/q39mLhx7SXBP9VKswv70XkRQfYeYdEa/nBqHfpWpOEFm3ur+TIZ609aXxgb6G6V3l9BKnGGRW
dnQc7yThOeclD+FFSSt+gzN1yKjaMzU0xG4mZPqicl6ew+BM1UZ6aSf+Mqlb5DH51mZqRU6kszgU
mKVHUOgeUJ0iHSkCXlWDnSHYT7v+PrHOe5pqhwtGLNLu0wnJbpX0BCbkLn/gOYknAJLu/QagEkIC
dRsoPt1S66im9M+AaW89Jj7miKDk7PDq56J/ezZdcJbB+yb2EEVXCeoYw7YV94Ue9bB9fUa1PTjz
ECMQGS9PfQDu+HlFFmnLx3pYN4SwH7cdovAtAhPoYzobrfuAZg0yIBIfbjmymr/mpvr+P8agchyx
Cg+mLTj9wm5utfJ2rhBryfZaSzAzMLtdvU6W0PSvjTGXUyjNe8x0fLe8hh6oBNRpbcleXxPmrRsY
9i5AOs1rW/Dpm4U7wR9sXngCLS0qZZWa/9KRDH58hHTMH0Az2kEeTTMPrBzVGzJQQQMbF/PJXxWs
/6yeQB931Peva1INJeXx3bkB7BocKvU2u3nN+ChgrMf4KrekjA4XxKRaT8jL7MQ0fL+VCdtx1fpO
a+mminIaDoqHhbD0rGsJ/85dl+qkAqqLUzp2BFeNfFLAbfYHRdg+oRvRB5T4wc9FR0eXlamCmzeL
DT9+bkZc6CbeeWwz+XXvOwfkSn07nxztxUJIigfxZhnL2+zPy3MlmPM/tjBJP4KrLUZPRgDDJQkn
pqfs11vaUZf53zv839uYjmbQGJKlL2bI/gyY3cNFE1RDcmmX8PjC9eRzAlE9f5di9N2g5iEAxVHx
aS3SVIVaByAbbvZE4Gh4DxdaJUWKHfHtOSpAOhkQi+y41sZpi6d/tfYaFSNAVtLXQ+PaRA7YSSIE
yGRFDAOJsDMfeYx6YE7lo3lYgAizmfkRxBOu/01X1GOFABvNoIEhljt+RgBK5REsHnz51Juus5Xm
jb7T5CvRiwxKO7r9Ofgl43kEDCr6hsV4kC1R4jd3lF2zUecMZqkN+2yKrS64+PPQ+AyV1WBYbeL5
KtbJNS1vnw8B+et/IafriaHtxH3pJs18nS/7wV1NuMy5KUOCKEMyGKl0thakH9WxMQ+mJnCt9wbE
IGsKw4J3Ga2ayuwrtIewm6rYuZ7qfXsDssYT3hRU04gZZvsAk1A01FAhn5NcZZLT9xyI42BDrOIe
s2Poel89u2hSlUsbbGyHx4RyOGaCYqQyLoAOAzNsnu6BKw1f1PmHjTF/em+640+DS2wiH+vDI/RX
dJ+AwY+OIgEucMg1VGuz3blnrU0YY3kgo9ynMbOxlRD0KFwacgtCsfbI3b5LBDDFwSGpGhzlcIyP
AZjycQlHxNH1jwD4/qh92zSyUyDT9bD40kfvpBr3TvxLvG+zGeYeENdOt/V/9haa+wmN5XiXt9U2
pJv6m5u4TP2JjNmbZpPrJS/pCY/qaURTrBPGYUWUi9MrNmQwkZ/kZHbvUwZ3ZlBmhe7SMXHC0wvo
mc4JSKTONF0igdUyOMDJVMHe5+p5S8MIR7NpEiVx7BrBQAj185Gs1kvaf52TCeyM1CgGNy74Ccbs
URzoi2Cg1UNMJ3k2Dzyz7UlMN+XoR2hBvIjopLXk+dWcSeBuD6+P9QvvX3xUVEpKCbKQZrkGwBLo
n04ESVore10wE0x0ZiEGGVIDu4knXGXtt9G5vVXST/iteH50ta5fhdOQ9Le+WVXp0kfTW3hjXFg6
QGwH5X6ii+hOz6yxL6QfbrTVnNWn6UPSDEv1nMe3ROWm7RZmGFgGv1zaDXDiRx5gRxJCqJ0Y8lam
TDyNgVVwUH+iyjqiMrmO8NioVWLmSCcfgsuO2Iw6TciXe4/rblysz6tBBJz9ZAPLLAlMu0Se4YAB
1HQjfSejZqg7xAkToZh8HMtkuYbWtm0gvArP0R3+B4r0gSt4+C9/51zJtimRnRsbbRmORrp+gYLe
nwZOSqZxLPysKzn3vyaoiZxTzM6l2IEgnDNqVtnRalZbHyjXGTVdkI9LnRVkNwTzL6MlvarKKeEA
bb0MKjFLR6a25BBMJHp9DLLGi9lrxjnHKrg0pnbqhOJ6ef2SfwXgzem2e7qafbYWzycCSMwrKboE
muezW7TbceGjlxZAxMd3KesQsRwSQVRJjn/8atDFBOi5OeWXoBNTwmt7pFVW/ChhQQG7GPU2m7b5
IYA63TO5aXKkAn/HYuR4vT4XccCndjgpYh0bsQldWYmEjITIg9CotyzZ+/54sMoqzH4vccMA2ULX
CRO7OtVMkJICkXww8f6MqfvcPYe5IuWvXRQg6q/S9yL9GuA1PHJeJPOnsa9EB/aaGc7zAkOKbS7d
gxky5vpdPwN3fKvxgUuKD1lX8/Ao4rtph5vGdCDFm5u7N7ssF+p9f72m50F87gkGzlC7GZsb6WjZ
C9xzIZV16w2KiVkaSJf/jy7xmMg9PMS+Exl7ZKD7Xo8XNr9BXNviw+yJpLjm8f2jt77GyBhMBxCy
ig2VRyHVTrisqWC1GbW/0N62TJ4BREAirXANWo8ugasS21MubqJj+rG54lTxrYzpUF4q2OgcWbcy
sGPuYFUtyno+Y0c6QbWWE4pP8I6qQVQk26yMoxfInfvnSP45IqstnyZBMFb6L1CwoVcmJnhYf6hA
9A0Qcyg/Wt3FdQFAsQN2/u/1kEuHaZO5hKEc0TBem7JrXsn5B1Wc9W+G3496ud5HOBT4MN0ukDnm
du9RZMEH8ccPrs/yJwoVa0LdeI9vhobEFzb965BJak6k3e05XemaK+ybcN9yT+hXhVGBetjB65ZW
DzSl1Vhof0SqgLwrTDfOWb5tCmHKDyKI9zrbPMBmbsugtZIjmmyf17zncodI258anL7Zqxg9N+fn
RajfFFDlfgb1QLgqWpwzqI+z0fB/4bb0WczljIFXu6d87H4GYXl4ESWjConQNwO0jbG8vijyTivS
wKcyB+Ie3EF+287eDOSnGvj+RzPZ1Rp4FWFFoWpFwHJHClxAY/twepGB/vLlYXALkqwTa66fP8hh
C48Wfi+DtNZyRIV9K8GOZ4NzG45e7pZDwFwEwvBz6cm9sNREPGnf+b1TNi30nHTnlJew6afn7QAW
/Q2GDXvkHSOXjyrrqpnMMlDrbKibfMLyIRiXOqz+r2URQzMsbB1bprYAvYtxKDmivVPd1a5u7U1P
LpgKUlgz0w1Sa9BN3xzk2FIKR3iF78f2eqARBdwgWKzpp+ScLtRB39Lpuux5pRO5MBdELurVecDB
ewuhTm39dJB8hvTj7/eGF4BSSOc+stCkJ6suhCLHZS3rf4U1+SAEmk2Qco2+D3IpjIcQphrMSiZe
dZe+R4+xN3iQ76m2UzqY6QFv9E6t1Xw8wY5N8Ij1ZfE0Jt+iPmVXAwJhUPhTW6Eay9XeX7QWxjXA
SRHwDOAbZJWeKKc6j4oPmEkybZtjpyiznj90f05NLwgwq8I1JgJgrxEkYQnRv14eAIGH5vajJlfS
AzHxACHXKJjx3g/zwJX7Lh1sop0U3WK/Gjn5Pw5UVwa1qfVg0RIfUEswPGEMgh4Tvx9toK7lHTPp
zt1Uij8AXJ4/rSS6gQr0SMxfyzAftctugMfNc5rZkaHdMGMfS95X8tTlYkWUSuPsN03nMCs1r7qo
EWwpwFIx3g9lE/FQ1EAGHs306wo0DgvwfxQ5g/4loOfOXkUkBPT+xqmROzTAy2V+RF/hwr7sSfk9
EXKRF8HnPHHbG0RtiegsM6DculCH5I1LhrjKQuOrQY2PNZWP1tUliC1j3MWk5hCNreisHeCQW8gO
ZTTG1x3swZhDmiXwhQHSJCOzP1tFfSmFv59NmahOnuQ/W4fOYn9Fnw8I/wXDtHpVjBAp+1/DIyF4
j6P1GYur64WdW0K9V0cr0pZIOh/TRA4Rn/8wa8lBlWchKldj+uYphfMpp0CIJPz8K8TA3f1FoKPq
YrpmejFD5ODrlQGXkP8Wg3arqWjRhHGPzpIexOpL5q2qW13fz5uDquJbtr+X2i67OwLGd1Bzu1Td
zrewxGxMIlU4SeAL62aM3m9yHbb+QSskFPYP9rvvP+wzSBC8QwQeklGVTkX/jsEedKel0J6bFrFa
pugFqXPGFjDAVQ0shgLt5D/twbHYYRpd+KvYE3/QNNbMO4H+J+z3uZ3hvKNlLwqIqxfldsv2yfdX
gz2yw/M8/83kgRB80ifuhlPS3r6DXTn8kxeRJjF6d334gT7fuRoT2LGgEo0BrywYC6oJaL5idiak
93dIwRQ2JPQYWUF4IcnwnsfmcKTMS8hsgBhh2PuZQJUEloI5gcCe+CNFmy1lYFgjgXTFVB9t+cx6
KXCCFCeRtYiOMzBvkf1jACx5jV/WVEDvZmC0/NE2FnORSFdxJNGGbf4HrsQQ1mgnqZXRr7IW0+qt
t3RVndRyfKndg6u8sxUm4vyiI18MdrLGeVy3mhxEy5hAj5rrkJfkyCYvRJzDfWaFJ+ttlJbPyzbw
58i4LJZpYdoX/JhNLIeJux8c+eb/GJ1xf/CfGZctZYijyLqh9wVriaUBT/BJcfxrTgMY4iOHUfSh
L3R4sUzqPFLNEdSAdcVttcU+66YdsUeARKdbFa9Ds4EqaSDfkwpEA+XPaO8eStBzHlkNVT0t+dB3
3XbPzo/QZ14XUsw8zZhK7eqrG4bm3KXcxtDEnAkogCJ3xOHlVbCBWTxw8E7K9Fcys2Nb6+PqvSUV
y3+Z3orIrFH7vuwmzI7DpfwS0P8NVrEijZC07ZXWDzbsR/UTf444sruA6BGpZ3As8YpZoLvyeIWE
rLMm+1TwYKMJxjLPbal+9uZJvvweuT+WsuOT807PYMUTlbvxNeotoZoRh47nyeVkVslxWjOlHUJQ
q+KDNcxBgnpKoOLJjOsFBmq7v4N5wirXm8espKS6MfLs9gRuB+SsS1MIxqkB2JsBNfj/pbJY7XVB
S3VNk06gDOjFeVArfhqG28VJ/fnSq9fhwMiP1LI6DfylEIqAiORa1ZfmkWR2iB5Uv7TDHt4Uemw4
ag/dwFjdYRler2ICKTgcFGr8FeiQyC8sg6W9KbYrxCUshy08Nq2rPys/FNsNcpvMSC9KYKOycQHg
8Xs5wzfUCKkZeuXJd4JCvm2yrv1lMG/0/gUqsjx8vye4b+6sphkG1sTMulxMHyJnxBqL5BDlOnT6
f2fXS/LnsY2t7a47i9Zb6ECiSGUouwgmVJQW1Z8VWWOGZ+x8tEKD5sty9mm0xKHvfHjgTn2yqFmH
Qfkfsp5iooeWkihU2nK1Nsynj0S4MZFrES2NYlzEGHXBhHXjZbUq8zVOZdum2pl3UtypP6zm7QOF
WNT+5LL/cZNph388Zj2yHPTiTns7F9igevAso8KQuCwP34PUu7nkCrsRMfIveQyENG2T7eWi2YYh
00r04J2icjlJssNO+w/iMOUJTBUO8l/O3tblu2CtrdnkpZPIFwLIIqvPCm1BXbSFQ0TiwJVlYqcF
Fgf0da4aI580OAb82LK73UM0qhQVcxq0hTZO6oGTF8FT7UHIOg0SGYLzTScsdnnsFxJF5E3EezHG
KT/t49hyBGdJgyUyxXrsC5SAmoI72j+7aRhdbocdXOH6vukRonWasETR9VaQwy2BzV4rP2zFvFyf
wTYMpXkH/zLCRYEQbpCutKC5V3/vvehK0qSiJaAxStWH2Z2PJuaP/mRiRo7ZxtC1hzql07G/aFgr
zDQyKAu7brppM7LlZeHeW6McytCq6n/o1AfM+BSCcFR6frQrLpwuB5D65VeV3TBDbh2/8qxkn+zh
h/KwPZoIWCKSgdLgQQ5FigufDjoian4RsMsEiVIh+L53XPidQWEokVFbm0QGMHytVQKa0UHh8L22
yH0fdyrcw4zwk14zgk/iplL0/M7MvmGiMhSO/jmrmt96SY7gIgzaU+IaKHu+kb/Hrb4tF9U3e8DD
VtzPL2EtpRcu3qBabkHTVMEjJnpQqZd2v+Z1bqXS1Vf8BTC5hyL3BeWqyqtMJ5yTCYEXsMc5JEJT
5uq1R2mzbyLqV1HEHIVh7yRBMma6Li/eHJK1q+CSf18PmDoTGSkpRzVybSvtbIDPgAOhs+IKtw7d
H//H68+zAOzf97UiGJ7iVysh47RruwqnpmUQMUXyhXsJBoSM2OQEZlA/M4F5bH6jar25nPt5LDX8
tB+hYiHWNRFX4y8Ee2bj6FiOKLnFob2kGGiHpSI1HXvXd1mbt1xU5CLTojA0E3VglTqnWV3Yo/xD
yx+tkazwTCeZqlGk8p9KerTA8Dk3ub/EG2HfUe4afX34vBrEFwti5GmuquifvFPTpleaA2fh+n7H
h3Efw+IgqmNYFlAcImfTTWfofaNYpWFU6vFlX4hRuY+dlDJZ83UrB9vOhA70EuIfuMcEoYTteLqb
YV35ZlM6C1IA5QQfjCIRkK+kwLu0TDEim6Wtfmoi1v3vu5s9YLcjUGwZf9BkWX8+in0r4GKnayt7
AxZ3UlbUU75tJ7Gzdxc3lBhI05dhz89NLy11IWsbMZmOmQiYuoQeGsIww/Mj7qMW8j1CT3MPUht2
PlHfiVIESokkdU3Gzz+TwcdlgNgdzuVMvA5eoTZwzTuMyKPd5x9+PBcZfzqEtHW987Fyp7z5nrrq
9hXjaxrnALUn45/WmzXQc7dNvnJi8dT036p+DlbhKmKGwwa4fApuYq4OA45gYPMDlojrOZQC08DX
UogF5FqvFFHd4AYysDLmcppXZc6JYK6buoaYmZBPvEJkcFri/5R5sJjbej/rjGufVhTp/jvSFFF8
G5CWNgtB41oqIxS8gh309y3BoaDu3tHzEL/Su8XoLuYp4uquSRrhhKTRCN7hxAs4Hqf5izYSQZRi
byL9wVv7PUu16Sa9uETw/mYnpWQMxVcUS5F4PY3PB81yxvuJwEbU2UBmgcuk1CeJqGezUtCrerkq
UTG3znRUvY5Q7a5TqsMefYqbgQ3ge1weqvX9VfqjLGn/ShW4F4SIFE1ljXjMXXYlsrMhqOQz9Ywn
qCIoF2dPjyT/4a12He8BpTCZ0cwdF0vJXaOsEDY0pK3Mtx7J4ZjQMz1IxYPFICQwmnsMtRGmeNes
JG3Ubt6+nERNL9BQtSD1kF8iUr4jhfsGo7yFRKB0Yo2gLZG0+1WRJmz7oeGBlHaITvSCHreeWtfY
RZRBOxxHoG3zak1/2FULNizVKLRU7QbYzrn4gDgKGahvp1LddNe2EOJILYoAwrGs7MReX3Nj2g3Y
dQ68EpJv2v7wx6NpzQEOnNKunPmHqOIuSr556cnjyEv1UsHkaD17dBiMnXXDPpwdcOt2uVSyR2Mo
gfKUAZJFYMJjGOv3ws9n789VscwqNaZPS6njpHdyIL2PhVrhf8qBryOMKYtZ7wGQGekjoTc5Phky
rICUgXHY5fmb0BRC6FRRKX3/OWYOuEGVhRGPaofzAe11UM43hCSm8wN+WTJ3VE3CZbPQb2pb6Gdu
DcLLVMZg3XWTZWzDE2BLq6eiVfmp7GjuBm3uHDbzysjbIbfPZsKEbiBzV+h4KOzM7Wvt1Pk6D7Lz
e/b2cLrAPxdNSUFgCqobEBJODnc2e4iuMWHwFutcKBxvPf3FfBhr0Axi2r/Dn98rx2dV0N/yekK9
FJVxBkA7bTSNCp+n/1CYsDlmQkdbu5BcsZXJLf0zKeD7t0MailGNrC1ztyvOXqHo237VX01927GV
DoYpsRftMxcVY4sLqDcnwnlNJ8sTwpwuBT3cq5ofYE8zH6xh5/6KyazHwsCPKbT5U6hmxYAli7Ei
l0FBASXvrhQTrV5/pQyXm3Qge2AtAPFcFmTFHJ6h+XPoGwJN68vHkqL6Jg0IXoUb12XtCKUvbQGA
z3WALtEcZE7gme71ox97rjfrPQkq4KwoLDT4JM/pcWqAmSqI3OSt6FVkR9BAFxKrduPLZZj2EcFe
5k+Oy94UcRBWZCo8BMCNygVyiNnYAeljcUUNU75NsJYvvOO2qTwAUjZV4Qm56uk0ckGiTaZf7ZTh
EDTHwdrIiavFr13BcQydunj10+vH0ArF2wUHKy3W7GfaylTCRSukKC4fEjdeQ8z1/4z4krbvtGTS
l9yC95wo/Ly9TFLuZ+MdJkCJ4bflEUE6dNT7zN42iNJ27Z+Wk3ZWmwX24edu+m/N/D4TDwIe72Eb
06K3Q4gEOUwt98qIBQqBzR+Jgm9+ZRYBwoH/cR19ES3oMRgTi4yBcBjG3iSRNmtL37ev+GY2Ne8r
rVpDK2jkJ53OEmp8G3bDO8sVl1p/j0OoxwbJoX9qLzjR/y4jnbhEguUSssGNZMPa6o5t+Fhv14EN
pwCfXHUE345Pw996vjFnZQ7VZwm+NDE1la1AboYLr3wh5wAgl2PogL+6yV+zL7hYvMa0s5ujicMj
oLD6hVPze7Tyv/OVvievoUMBLsIP6ahZ7yJ6wXvznnNnrV+syhVSGpcK/YrRoSBsxjctyl69Lx3t
UvP63JxoFCM9Er9bWRIX6X+Pu2nNVYx1hAlhTY780HOwziBhvML0JyGvfgARRjo6UM5u/d+1KgtV
AQ/jgetCAC1IqrvHaFvVlg09zTd2bx1J9Ambm+qoi/S0M7+nv8C6m/0Bxx+p7iIaoTjKgkBQHKjT
osgDKsOGc+NWEWm9sZ+sXSU6kmX3IOKEWn/lHhG6PL35bkBVGMe+45+2N51J7cJbbGHZYhp88C6H
XAGQ+XHyGZIM7Htcr91ZCIXPyOdR3lwYIpZToA6AgCkHM+pup8d2QB07ALFFyG3n7mexuQjDn+kZ
S7W0VCZFF+k4W+m22PWrsVBmYEXNfR9jGIYikP5ojL+earQnqnBep67JqRmwt0bBuQ7ZD1qYx/8w
8vujJeUZGFgAKsV9ig4SqULa6YG38RCYd1mwMuttdgVSRmDdjb4aY054Xmn+RceZziruuMtwduRV
ALq4XF85dCv+I45s6NWn0eZMna5F2aLCgtOi+Xed0z9X8v77RE831g4ptLXCPBotfnHy+CLrb+Qw
H7Gwe16bdpj9EOwDcxMNlpkChtVnRYEH64r76/4lLMezhRqmURNqbw0yKgk06WaM0dPP1wOazIyq
/cWrcwidN8T3KTkJ0cxHmswVtd0I2WThlYMqFZCZeC2MbvTTHIpZysZZuGCHshqc0JApDi2KNdDd
nqgplBTxCnbzRwh02qbJJkMdvJNJJQYMCCvuTsJDpKFA09JfakBXjIliDbex5tD1XnYkxHbW0JQw
fHIX74lAsK/GWpwbosUlUypv6G93dGsAoMgiYAJF0K50i9eWve8HszLKdlbXewtpndq8GXy0zaOp
yOH0lbvb5hwo/UBANv7aJhtCjOf2zQDfXfvg1Dova9accDf/gDnGldg2Rgps5wXfdLiDZMxg0ArR
Vg5VHzdT0TuTMpfhStjxFKHHNjxDGq7nc72+FX6gWe62dQZQTgID6WSpfpqRUrllQzYmcHAABMil
JveJR4FcE3wFnbtbgDdCuHQhpPKR/Xslmk15t3V0noXxGWjVlBgsATcyJ5PX5pSdlbXBYEQiw6W/
jw0xaiI563b8NcUMtJGPJfw/AdzmgfqxXlsRLwLo+mQsKS2nSCMKcVYoajPpzIYdvyFdOil0l+Im
VtPl+kYAOIgaR5SsVH5Mv7HX66kKavewcUu0W48GuSVbOcN1MZaDJvFHi3x7aoh7YluPnbvOpMkF
AmAQiBRbnn+3ZTCB17CzcXWhQOPEN+EIA095DOfQ3woJj9v/e80s0RD08Flm8Of/q+88LS0Yp9IX
H8cpIzEmaVUNchiqZ/LoWa9KP1N6nXc7VJdeo7yUfJ3Z3irq6ReXNnhJCOCUFSNIGyWvNRhxMvVX
tyNdcT8GnK+wif+5P7nLcqcKTbFtZaQdGOXNp+IR6CPwZRIpPkabMdc9JvY+myZFB7QeOb9KT92c
aUBmrncfvs9T9Be7yWUCv/M54X6NmjPADjJ6vJZZqwDP1oKt4ty5juY9hREfVBH1aRvsm6OxiiRZ
Kr9/V7MBzb/k2TeV6qydYVyVmq3q2ZlAJJ6+TNtwqqPrX2taGwAAfE5m+f4ukMS9dgiN+mDnfDvS
GeNnwccYoK05os8MS+5aZLtxP598mHK2BKHK4ClZKaktSHzmtTrJIyfQ3MFZVUBCJ/wFQTuSN3DF
QeTnRy632zG2rbu1iC6GvXx1ElDMRQ7jF0NOfyyWUVWydBJWUSyGi5fnq9WTXt+vhY5v4orIWtke
8Gu+bA5MA2ymnRQQbTNMt8lMM77ejAMsXfKijf/QxrUWS8jpX9LyuPcM7rOW7a0rhfqsmd4gKR4i
VWUI/ZDtRo2NNJHV6ELyWmb4D3DITRONQ+9+V9RwJ0U4ePh5fIYHyqTuOcGGRM/UxU4jKrq1bwUu
0uEiAZML/LFThAkLDYws2d0L0YUkMhg7rs3GI/PkY31LddMO9TAJMN2suwi8DsUVWXU23J3NlPV6
cdf3cSa+bjfz7rV+qUT1TpQuT7aMIWWGOrTVa/Vnk9sZqPgoevX7bLBViAGQaKJddX/t5hzTYPqh
E4Ay3VAMFsuQI5GhiXyyx2JB1nT0JzTe0wOfSuqRRoGfNDmCBtXh+vVq7EMbyXABOvFIV0HHIJJy
GQhnU3DxKtOZL+0pJbpvKSG46UwFMK/+5FKEydF9+7LF48AUmlsD7wsPMNrWHUuTYUtOwtT0gLh7
uZHNLYxJHCSiGDFHs4Y9PGgub6C0vz2a9QovL/MxKsjsi0bQjXCNbSjikJVp5fEtY7+dUBf9dq/E
8diMCY6x4zUFE0cvaFhobGbd38Y4DvtlCXsBWzsikOkTPRAI2lRYEywoMw84oF2P6/5vH9R1mpN8
8O7ZZCb+VCb2MCPWCZxaOmrfgicTz24UupKmjLZgzIWaaAS+JUNkDvoWVwG4PJDa3iiZjdV0OPXa
jm4dOaice+vrj0qMdgilq5/IZENMSxICS2/7Fj9pDNlBYEQkmlZYkBotHwlWP1Bw8R1RklZD8a/C
oAohm7C8oFdBX7BRoxxptB5VjHkunCt4FuZCZvSPrCkZGItwk3VaA8TE7GqM/IiZV6sqpf0h8HED
Gx4gJvzjqDzHEqDuokwJYviEJm4CSc0hKhxeT/6eO1HU60h1+oFA3ov9RqtIyc+fbXsoIyj4v5V4
3lAVfAnVDLNDaE3irarWlfH1KUiipdQaDD5HKtKY2OPSrbgIP3iUH/2HneyopxViTJasP9I4zEeS
pCaglarUEng+tkWQBPVe7IUDpnVBmYShp2vNub3LwvaIY80W/DeFCOjA1PlwIjN/0NzxDPctxdxj
DTu3GDZzGcmkMz0AITrcftTHdEBZGoT0oa0LHZvFBT/iKxRxC0JY3o0e6wixdm+W5PVrW8v4bP89
6frVeslevOihacvWtHZGAFJS9drsWPajB8MQU1I39GxcqsAj/Cn3HyGqATbo8kcpY+QahVqdyR9R
UrZlxGUXFcQ61N9oPilkOIvS+L6C2+G+LWHGAKqKjUuywMgqkGC8FosMvQ4iygkiV7Saegf6rz0F
B4Q49a6BjGrbkrbNr5p5l8DRFqG4c8WBaH58+DmQ4OV/IusmzSKwkrJtBEg+JnytVpXe5A3ez6EP
iywDIa/tckhR2rmbiKpLwKzqup4+CB7QTtDqloPzsMqlsSz3NA5lKUtilzdTla6YaJlXw2aqKZBB
b5kkw7KYXRYySkN1tqzCwG5yZ7FWbRyO+eXkHj8G/j8DcZ9hYcyLx4CBIVC5eNgVaOWk6ZtCj8Wa
3neotaKEJ2Hk7HiO44cH3SKfK3U6W2Je2tu64Iw2B0Ie16ynNxDfuvMPP/yfNWfWhtNvSK1fXFSl
sy46WnwFoGYPFQhhS/bzAvkziGz8wg7O+Gq0a456fm0EPjZ1+ZL286gGhUOsvMEu9buWo8nmKzY1
SY+h2AD8t9w1PdHqQCWz5yEUuFTJ2Xo/xOl/H4c/6C6lvSexS9on57sARIz1awlWHSExHrySx2NW
FEH4InT2g83l/GOXwjkXSEbnRb3KqMbz28lBTRW+jpvSCRezlkOCybEuHEqZTbWeGQcLTGmymxBs
Bfg0WrSE4FyE/HZyWITwKgptC9/WRfjubFnaC21E56gAA50KR2mgT19NoBfKzeAHw2csW9cfMS/t
vVuB58SwVAEKSMB0qoP/rJ9a6zbgazoYsS/gVdK8E4LxvrRRgUpa9+tQxCdo3/H4Jm3wsqYodwiX
0KvfnQyrIVKhUTCfsqAMfKGeijk21PxaV98KxvrloISM8frWKiv2rknyglxtXAWXpijSfAALWzRH
V1SQIVJcvLIeJ/9W4h0dZTcx7SWcXJSnRZyr9BXAo9ohW8+l+s5T8lQCNTNLhVZ900h1dwDJs+7K
gfRLH8+WAW6DaqC5aVtyO4iAr/edc9Eu1naJk+BICKkqNARuDQq1lveXjfTCyhWI6k7o24JMDpBK
4nLNX8wT1Xyammc4SYYokVWC7j0hX2pkN3zG1EfgV1n62btvxwaNzCNA9+wU9w+BoVW6E+WF6jCW
dLhMkhzpeyNFI54nelFAB0iEVLIO9YGG26GiL/htbcx+/FwN1lLjw69xYfXPl9cWem4kQnqW8irT
C+M/Gwej9LtYgdUy5oHS5BVYX4T1EUPjllEbVlBmlmO6jU863LgkP+cop2ipFFOnvRHPP/7Zdo1a
80nJHvFcuVlN2quSzw34SuEgbQaeXuzjRUDnAdKX2KMLAXBFicWJAgf+Wwr8GFDnYmr047f3wI45
wrvyyVS4q5YQvU4SASNkcExO84B0A79Su8zfqWCmplk5BYqvQQ1QZFFvIqENq5Q19WRnID7PF1Ox
HdQD+HNllabEJ9HWsi7uO/caZnL+RcvKULv/KSqlcH3TGDL6ifiGx9KVaQ439zoX8e50vqtgjnPM
Nx/xW8lsXeOeV5Um2FoZ6YWvQrU9vzMMUhYDdt5wchzwu1RbSaE0IcWgmgkmZO5PU3ZJlJcTO7AV
yaMUgy2AxSXTT1+qTqG1vjx1Rhq/KmNvEzueJEXRMiLDTSxR4i5Qn9dH1Qcz4U5KtV2VQ3VremKL
xCSE+vYfx15S7sqWCxOvcwCrJO3vBsAiU0WlcZfQdV4H+qu9e5DNpwGf5BhsvbmgBL4ovw63XqKO
AT1tW0Dt3a9qx0HlT7cjawpb5/nifM0eHj0yR/G+hccW6Bfvdd8174qs0X2Qv5W3Yi3f3tGnQM8K
vDLgHyz/1u8r/nkK/MedP385OhSBfgoAMGkLD+fmfDoXbtV5uEuSIi80UMQm+EOiTNV3lo/1GAAy
450KUKLz8FKaFqDOOQ5ud4kDnX+zFtIMTKcAmZ8Usgd+K8L8snd58YQPL+sb82AUB7PuHDc6XIKv
F9488tOU8GNtouJ1ECBsGUBs6N8z6c/J8LWlqYrnc/+aqEoEjYkLXS2GpwYGp4jFOsAsB19b1UfB
AQeTUv/Ph+uIDteM8O6J6YP91srh1higHP3+ZqXEJM5WY16SxC6Y0z1/ZzMTh21PWxV0WCTafepp
sn4rSFuTQZ1gyxB4/PfWQuvgcRcepKkoKTwvPxHw3xXbsDSpw/nYBOpwP6n+rSNqMPy4dFSrKjdh
hvQNZYD5K9UfdKMkBw/fis+GKrd1oNIY0r/wCNghYgRMq+GPLkxUT/raRrg0nWVPOHyIRj2AOgmU
HHXAWYeM7+MeyoBxL8LO16bo7eTPUItj7+qxXF+wdhF5bW6xYFH1xMKnyf4tDF7dANCHAsd1ww4g
dM8LhnZuwPsGTpToMF3835x9ePdhII+lbTyuRrhRLXuDSoZLUkMIkRHEt27A32R/KaeVW7tZ9Vh3
PTVnvuwnPUjPy9UyKH2YkpiPBa9Ri24CKHoeH0jAtUcgdjogXpNnDPMCn/GKoEzlvr5a9WLYVrJi
LOEb7eh0rOeGOPkl4m67O8nyx06qCnYFCOZDGIB2lJJX9ERPs9nHwd/2yfQsXp25NlS3O4Ifb9ir
CJTv9tNWcNCeNgPBkJ1ujuN6YtaOIVcYNwrX1oTgCl2ZvEgMwndD4VZqUrFe3gCU38WodZRoEudj
Cne1uNwkdYLsfbfu4uvgotA1Fp4PGHrSpBZDEZvcP7f5Qq4FekFGgENrJxb4VhzgmlP5NWDmJQr7
yX5oooSZsbxAvbcB7EbT5ElDMWL8+BR8qLIZnn5lyaO1mq1I9Qhdy5QQ86M2KMtpTCqNOFbz4FnV
+od+nXrESDPIicS4I1Riw86y8xylJ7YQyc14UsiWBuJ5gKB+O7yFO/SY9r3o9S4uJFvxBoN/XzZZ
MaIltRQruOMKrf5vo+gnHglj1BaUt+0LZuEHONPDC04zwR3YCOLy8S6kPpiWfbCazYbkl012AKVt
NcYeBs9LmZmjeVSR+TQS9U+vlJvWFL6cRL8Cfv5RcnT8M2txiCDYcaSESMip+YP7edIYvqtDc4Ns
XokM4qQStKxTIbjbYaCULQdc9eXImmS3pgTncvFphSL9/HOtm80Vu06Y+6pLQW0uJcWHAQDUHD8r
fAPFnMkUziX2PGL1CDn5Oenv1b6R2Bbw/Y3rBe6PXLN8CieaGIoCjOxazkix5lWM3eFGNsWTLHEa
oyLT5BWLvinvnHSZZ2x3lbbERtJh/aUjD0jnjSgn+H6JQJAoASpQJUnMbkeKfyKMIwftePSGAFyN
mYGg+/iNLCR4FIRBHPw9zh4gq2PDC60WKNq1hIl17PbAwPNULBs2JrgUwrDXOYx32fd6W2PEM4vS
ykkrh7is5IeePNrnyTIWJ0bbQI2pY8bgPl9ve3Bz6LH2Gdn/4PHJq6YXx8QMYP0wGg5fTNA3SgF3
Z5/ydX2uwdpP6R14l1UpTDF4ppO5iRmkee57gYzuVDHISHE8Km/hE2XxTboAPMw+PFSlM6lfUeS4
H2Yvnie/XQ27bmd11YZwK444w46OQFlD1akh0Uk66lkLzrC1Ufx1Bgfqsi7L53usgNC/E8A6al04
PKcpug+5CSkIYiuefMD3qy7MCiVxQcWjI+w+WeaoTRf+8jMYKmTJEsV7gE8l7umz28RbeLR1OL/h
bbR4FwMxYwMPKF3LXgUsrnYY/jYfl3fAfnkj0Tp4GHMbn181BVxB/uMMFEfSmSM4cGBkRxcx1Whq
trKm/0rhy7qOxhcPINB67/U3m3lsF3JClAduZiAfKjdbbUEo6NvB12s6y3dD16aHseNnyDwvakUH
WjMLF6oS/hLltniXYMh2xYk4foMp9I/vkUddnzy0FH1T6g+Q9q/3zOIGYla4ZfOCO6HthA5mhRYM
wFl5IAKJqDApHOtdx2UWH+ozPz8Dho+uuHVymjtt5Z2troO5uXuw3AAhIslgnn396eLBuxoc+IUv
UXNk4GiUlLU1cqLPmx0HFkRzWWZbd/ngOpz63JnaLCOucMJlxn566tMK/DFCRGI9VQ0owGN3JNDb
egAifvwHeXg5+KfHeDk/N9BMD1NljGTN+G9e+M0eygFNxxO+rQYjMS9F0EHwBXSX8wXJ7Dh/HPmW
J0ZfSIWg7fDPlSXqPSV2vErAm8QQ91ijPFEyvgu+pMCzbTO9MitD6dBvk7tmLMKOnvWOFHBb63P9
za1OPTH0luucN7QynBqxRp287SLLLgJenKuIRKfK9ixYvwVLOHLB+mOON9NR7xK94O10VJQ+extN
kbm8d2zuRFKgcD4gvjTK3jqTGlWF+rFX5pI9wInoIBFfG7q2qWjvC1hYUcnhNpSsjCbJ5NT6jkeA
UmQS/+RMeR392b9h0sftYLCEsSXDq9U+v/p7nXUyhRtRfc2MEeZREb8UI2UwDnex3fU8SWo2M6Dj
foNKynlXvKHR7KRqMEUDoH4ch8IAw9jS92ebpShiTsf9SBwNv+ovWJClEREFfc5EdhJodogmpDzt
TpUX+kK72E9G9Vdb4el0CL8cji35m2YezHi5znO/7QIPWTLrHygiPxRgxEE01LtczPRTIhb0LYTj
4ihjcqaZzc9yYZHM2jtZgmkEVETTGT7nnDzfe8lOnQMM2n3vlaUvQV4XBsnMt+kp/IaHrDzHyeeI
Ku5RalzAErEguCoc+Kn0D4MAzKFMqPIN7BiAZdTY4EuTeF2fZrPoSSciB53rUcO9tohq3OOy0Kzf
A0amkdBeQKuTjBerb1CUM7Wuc7kcN0c7yuDwVPrlLQZ7w9XeOGgpQBunYumeV8pUdXNa270XynYb
zD2wtMk/GFNGGfpA7tuY7tXIK/ryP5zSKREXpTL7K3eJYBvp7S3p4EsY4N0CdUlQeFukT0Hl8cnu
6k0yphbVxoSWSS8uhGPnzCnjp/NMG+JytkABnVRlYGMTzIFIvFX8lrasy4DalPlXkxFRVDa1wrFN
Xa+fMy9+zAHLtjBMCTVmXupK8IZcNB5l3kb8TQ6jm87LOsfwc+qqIEfk9V+4XVzNjwpDJ4WdzcJB
e+3PYMwoqOjVNjp5Ldln36iP33XXEiiiV1QhGOX+9zyFSkxw7WMZFYXxe69QrSn9ywgTIllVlM8r
DGgB9IC/udrclKckHGo5CORtEN5dhpzylZSQ47ogteh1e0vVWWiXpJNbdgfqJSEZbLzqQFbhdvmP
V0QFDhpgXx+Cy4lQ3SsVgtmZPBS3tSTu00k17fwra3iUXGx3asdERy9Cw07dIjhdCV9tVUCkWtZU
ikAGblsnedBk64tOYGND/GzatKdhCsUIwSgBgkDR4mMMlufDpnKhoC1aX1u3Nean92l8VzJJEO1l
hS0C5Ch/Arwchyz79Wcf4Grv/xXl7TCM6XPNaraORsIY5Kf0ORMtZDiMQ0pQM71ONZPO7G1rCcSC
/DnJQ9nZ7PiV9F70natNSbZ8MnA8zpjf6r6s0H5epcwsEjtTZedfSqGb97Nf4gcvkeoyzHsi2Ye3
ijMWwCTVySxVA65KdjgJuQoJnP31MajqDN/+a9aiJLrw3qxAnOm81WCqSALIrS2egXXS37MYaXIz
YiGppPGVILn4utEQvRw+gkR9/Q/RNncwPLjek71ECnKXNlpUiODZC1CuhDiYywQY0TsVp5UelHp/
6i95MvxgeEudYZqtaL+ZKpLOkegmaCAakfS8xEWITguZe5O6YKM+7nd4+QDobKutuXwZeF0SvZ5P
6zF2GUMJ9+TSwXfyZU7IyPE7VnoZWMQJyGQ3bl/1tp66gz4LjzJ9R1pdDVRr0L3ytUU6SzyL9N6Y
tu9svQdIxr9E+zNzbeuufyqKLcc7Cf8Y18obtI+8w9aF2tnayQY3wppNkcEdYZK82Vcv3xKrsY7B
gRmfQap3jJ7FSFBXHwyj9cf0Muuoxe30DKgu2+OkEI3c4fxULS005kg4Pndoir5C3WGe/HzyNn9W
n4LBP8JMdokt6poppyBOEK4ow+ISNBWV8hUmLPiirjwCctOKMJtRev1kdSY5TEW0NevtXAQBtQ52
nt/iUUOU1dGbMHhBash0OLhXDmJFoTNy1JyvAMA+Fyl39AJmz7QeO3mHmgAj4H0RpiHrUZCaVS2R
OfF50XaZ48uPR0pOwTERprMgrCjwtxriaQ+Wxwhjxq5NYQO2DlTlcdiO0zXkIImugtLG8svwykSb
WGqCq7supRW8bAxUoGxXufYz6TPWMrbH9cDxIkRa/IpAgrVHjUjMpn2JHnG3MfuSyM4xbvJEi2XX
nKreP2lVtajLD9jGL9riInjo8P0w8dlA0F8Q6ih8AusdC2uqAb4Fim/lTCsr91Hv5bQyy/bwArLw
ZOTx0wP/L3+7y/aHhcT6jXjIIn9JP9dHB2xhBc8Pgh/rWSU7QHsXMf67xJr0IsPQVpwPJK3o2BVX
6fIixqmhJ0a70sWQt4nCYkr1DdzffGwNZfgWd6V/LcgkzAZzXXMz5Iu3TTLWfyzdJG/aQBmyN3P+
9/uQSc5u+u+Pk5D+cxdZS/imTDqupKITBfqHkfUPQKJ3O3Ns0ZUo33sRJ+555nJTMOKAx/YlewQ9
QSUCJr6nJ0DstwAKmRDtK+6V038orrAhKEs5FBzZdbDBS09jlURMjsqw25LzVKofeitv0dMkmtu0
ZlJUVaq/9omjcNPZxia96T8R8hsUzRjYyV7kMelumxIR1YlatrtKArZFAgo8uRpt5J8N4cHAzaev
+ZU/l0KAz6Z6SijHGOO4UMR/RG5iOKTJeJGEd1XE7RAJPoIh8y/WnfWxHpI0U35Ptvp+sxQEFhrZ
24wvvt9PTubn2o00vDch/DMnSBra5jo/8nEOziNt82D3eL2N5gv1K2HOYY3HyS4uf+v7BDs3hfNK
lapfF5OR2MVACMgI0vUvtpDhN5IqQnX4QiB62zgBxblUk5Jbqs1nBU24qPA/Pw0T8XSJS5Ek2Zgd
+Ly9grhHD9O3wwQAR57W+fPniWou970Owvl8ules8t/KIkvyUNAuIq4+w0T1fRBRVo56Y5CS/IJ0
+MpXgjMzhjnum+ms9PYiKXNkBeqMeJwOq6m1GXp31BdeZdCtXqcFaS+XqBpgbZ3m36hPr83niDk6
SAc+8an9NE/nzRW8MJB+J3RHGjLcXTzhjBPibAak/8MVzZDNfvqEGR+NToYQAYAH78R95Rxcex94
NNWlMUkaTdKlMjpeH0kTMSBrx1YuEY/hwQOUorgGWmaIZBtduXhYTAOAPm4zQx1Rp0n4IeqgPQg4
MQ0o5EoR3ZKKy5ByzOKtBGXTCxmbeIlEiuRgF8yyDz5nQbjIVyJB3zlvm8AUzEN/GcWlxyAl92JT
BcCMGC7tfgSAiCnp7L7GvLYNB0ZJWnl80TgAXaPuGyZGZKz1PU85X3d7xdcx8dpC/WWWNHwPiyR8
PBHc4mUQFt6eHuVYcKz2uGOSuzrzjjUr8Arv5BhqF1JzzS6MT0aI100Jda0Q3iY2h7Rr5uBDgs5N
ENMiZFGgxhID/OaV0RQlri6CB0C18WXEQ5Wk5jrv3/a0QjexEYyS+bPaX6dZYDboB9YT5qO2ehM4
iRbRmbA2QiPoOjerGls3dKv65/WouVmXuZNdCfU1fLkz+bKn8hcP/v2ebFRS9p9ZBITHTAWDpras
RyQgNnZJ5gis+YjNGQuVexTcHtqRmGrYESjDIJjWorl0m8rn0IO/8VB6ThdveSzHZgZDxOcd0IFy
IwmnMvgh4qJqBChhWYgtdHCeSxcK7Jyvhbbki4Q7z+XGWbLncNJ4wrI8vWdYsng4q1K7DQ5KxrLi
UWh4JpnPo3msX7B1J7vyLHs08aNJwlk51AMYG7mu/VZwlTYxZxh8Xq0527ZDkH0j2IEwhb68RIu3
9fnamfeX69SoRBzYz4B0QyNfqPNu2pJV8re+kNuC1zkyzFDeHxQRNB6MHXqAQYCxsUB1WWohlEzd
VTYKcW3I1qdf9nN0V9raayxB2dO5TdcU6zaoixbTfK2wUntSrdoOsrRSybZhrE0gJJBRNuwgYs2h
6+aEQSZteVrJYcZQPy7bpQdioKhoiLr7oPgTkS1vCz0X84PxVZag91BbJYjxxJOiQCLLjkU5ulsn
8FQsF6J7hZHAxBurZtxG+X63trC6gL8GxVPtXWrFvq8zeXVwEd+duv2vnYgz8URMHnDyW/gpePwL
GyFL2nGMFIaOwfy9b0w7N5T0rZ5I2tTNpbxGRtEWb5YpT/PxwvCwvndxJldA/J1YayonGo70v8vJ
M4GtvlK7sSSpUR4WiMcK6IL/GabVU9EV/NHhdqXTW1OdNRuVa6w847YdXf0QBUTKErwrcETNPjeo
HBIy0IV5vjvaXJj0CnCmvyFo63+ZbRCENHKlZLoJhzQ9vLK4M5Ut6wAr9nKCCYS+c9h6/ovvbR9y
cCxM4qMA7tIQWj6oCEtosLDHT9ECWaFrBcrInc57uxinZ66cPVtAtZzD3jb6yD+dfFbKs/t1/ncN
ydjtfMvDbMNZUZsFPOjXuwyhY4Oww7rBI3b/axInDDxljtz9IBxiyMEjW+elV4Wd9nlg+nGjw8VW
xPQSBW9G4nYPNv4PQZ6WYiaQU11I5swhrwK+oFBI6n3ZGgpsP83jzicxpbA8rkxrupqKaHEQbe3z
lHJrW7GkLZJ6eEoJh/buewPIYyE1bxAWNnxdChOBgWp1a/RcSKyhRtuT0O/OelAmzmn0Bp6q8GS3
IjECkb+zcZMAsri8x+wmT4W94LtKWrpLpPayvi92ioSsOFWxxVY8o4nB1711PrxXIPVUP6k0Blsf
HnG8DXJnP/l13ORLBWJbuTOml4Ojbsn+nzSCebKSJ3Hx5hssP+okDPZRn05vWuTnb4TwM2ij160O
LgKomzJ5CM2jOrE9sn0w4ezKuVbK6F/Bo3EVXcRI+iwcZ6MszPSR/s4wMwTZc3y+y4agN6H4rHLq
BTUvwR8HHRkLx44jMWg8b8AugB3e9TjKlpGTsIwdDB5psCNjKHLeIsf+lzocbECET5YzrAnlLQwU
MRBPd6KP0NhjL4wsx/1kqHzDYh2p20I88y6Kzg6TFtjquunYmq70ZGIkynTrSEJlvgTDWBqpuDMt
OTT3dTxNp/711stGrunXjzzruCJRhDD5noSg3pW+SnEJ2CNRgj/o9qdJ1QRj92wa7IcU5Lv2L4H1
VtVTuwIm2O6lSElevFkdA3qszhyoWOcxB7mpTYJz5su0PYugZmzZx3H5uvNiqDDytKFcvJhxCHt+
q4M3PPSg5ze7TCqS0jDXmmlhN0h959DPQEvQPP11tpjJJ+4c7FO3GgULnpxoC53zKLpO+mtmuu9o
j4wvNGPXufTEWGI/LGv0/L/EPdw82f8L+z2OiEpPqYffVYliuovcJ7UAVmbUayzrPwzDuL/VsnKN
MZ924+BhRhzngU0OzTsf5bujo5dvvkYvCNUEUVCbvLY+Pb6mE2zH/lJv+6vTWSuugXeBQpQF+fhx
lBjhKo7jvVOJxw8wEBmUAfudIPssfz+Vcj5YSyxZ34L4XK5Vr84KiUNH1QKPBZ9sh1+WrOoNTIvn
/uapVvRy608y0at5mApNvdvf/QNBh8V3707Q4Uazm34qsoIDVvRmv1tPxR9ELcUof2nT3rxloLOR
YL5J6qSGmojfciJNSTrSincoPUMAvRmAfJ2pOIxhxwnMF7OI6LtzRk3jmhS4MVGOr9rkPVQ6HRzQ
yXAge9mYhGB8lU2tdIqnGnLsEUnzv4dBDF9O2bB48s36uSFFZunD47y/Hry5PSUOvc/VS39OrhdB
ZWLteI0gykDKJzjrEZ8My5xKHTUVdsD7x9PrCSqAy87tEorlTO53mIDmi4MyUwL/5sFALPe7mUvE
G94ogOP2Q/Hf4GGhsRLTioXz4jl8eu0qE4GowmE668zGjSW4K/JRvSYGgWeQ4ZrnilwdoS538kO4
KkKAb9bnqy0+Vp57YGSn6jB7jpqwOyIkeRZ4mmj77C1R4CYsrSkuC5gTnSS5JYaRFjjzCeZocA9K
Kr5tEj6InVbaQs+G7Zf7X4HDaJTKkbexaoMsKspKSxoyw+oU1P3q9PfNNqVFTIU4V4uH5EweZO3W
OTnC7uOAqDbL4xooBythZQTOd9c0z3bR5lY2v5BxWh6gafbjnyMSGa202Cms03tq1alhpSumYPcK
+AnDXRiPMk9tn9VT4jEsYcKOBT+8eJFsxLvkiRzZ9gjqffyXC1NF1bDhfzUcHe3uM3Y96oOir7ov
m4wh9bvB64zks4VxOg29nPfLd7yoGjIkt1rlibNjeEkYJSKDE3UdrYGE468bEiUuj2cO9CPk8aqA
R4RQev28GcZMJtoM2Aq0BKuNso5Fx2cX+/Wma7I6Lu3n/vLeivyWc1U5PLAsEPz13mYRgBzIpIL/
XX58/n+RQjP2c0wfF52kp7kVl5wWv6aobQddU0wVA6xXVX+qxi/NmFMAQa1rOwSvYuDDHWV8J5v6
OJ0jFNiCnUyEhbbXoRldpR2Wau3SygbAbKS/KDV3ex3ff9gt/9XuMctvrfDyyFW832P7pgLphfKE
DisTfIoBhtTNbkghW7z5sLMQofrrf0HflMgEBLEXV41XA7w7Zh1EEz/1G2wcdPZabkgvbESTNMlv
apMOR9sYlEKJ25vhoNwfGQIUSze4a1oBlrxl2kJ6NjYRqUggTHtjqxM91ZDwO80+Q0aTR7YJpeHE
GFtOdej3YFKqpMV0gLj/9BCdzbQNYYzBf6lSQTNAZFpV64oI82Vcd7dbpkUmi2pJkDOQA3CtRET2
wJ27Muernmib0MxxMQsmtDDJ5EoVCcTVzmVOAYRRpMtnxtTvFZml4i75gZ9U4MDOfFJ7fcgkf5NO
gFAXpoqXyR5jGKZeR0sjyHimzAY10Eea2xsjSm53j/BlPmtQldxYwQN9E0G5Kd/WxsWWCeF7YL/4
2K0hmU1503dWZIboYWVOVQR+7KEmc5GkJTOo4C4P8RFcmRAbo/6mch0JfgUjnSYcPWYgQJDt37+n
nV8akI1kIu0U+RaEKLuE5Zv3zqkJH9ppmAclGlPUyAuTy0piQFcAOM0Tp7I6TbgFXno3ZUouMzPf
v1DWoEwfM9WwERJctwcqXpKO0xx4pYNEnrf+6EmXIUlRx64sERUDdp77micBpryrxFUj0U3WXN0y
Lr1PLY5x1vbSCe4+4MNUlATFvYZ5klQgV3/dtEkPE/appeSFOybveEOZ5jY/D8aW4zKoBYvKtcNx
o7Xvjk1k40wNX+To/FEEiuE6GWZYiuRi+LQalyX+BjnzCp/DDn1jrcHWOb9Xkofw3OPENeA0/MRI
gMqE4lh5hYRkUAttghSVxiV8EFXfP0FRs1vvQwNlyLHRME2Yg4cLObuLOoJG+9eCp/qgp9UQNVm9
4Bjx2oGFwlFOGCCN1b9HVo+3q3uV/yRoisjk0JWvFTxfnsfUVKfzWCZooTIdxqRuItN5SiZvLOGt
+0EHZPajQBnRMmn4PFoC6JXbMJzyrY2tHqXd25PYf06mle18OD95+03eRvoZA0hhXqOS/FLj095R
jGsvikjY9UiGi9zhGaF38xv/svxMqJ4n/9qj5XgKrBxbbQFhRKny3ZRN15pckScIcwiR/0HrZ9zf
bWCzYUPU+xnsjrHARVPs+QcgprKy7wdmWaJIm1R+oApxlerb/7ZIsPEqvyU4wLcSJ1gQHxCU2ezi
2Wq6gXH+xgeVQ1XWB3xggN03kSTvy2Se50GsjeHj5ePXUIgb0knAgTvYxp9XbMTyNGG3EdZOcQxo
M52mixYLJf7pf/j3sg2sWLeywZCfIDsMWIUK1PAyW7aG0vovMdMk0KpaSidR0/Ma7YC66iSCFBIk
ciJXfwT7Jk8raKFjMkLVE8m3m09dy9G8w5mueC4GE75TJzaCqmHhN9yEF0Je3Z4aINb4+XlecUXo
f9vhDbI4Z6WJZPE7LAkCMKs0x9KgeA+k6U2GOYJBNxn1YaxMCmvFoM14laTQ56/cDjQa3+9I4sPU
o7Hgbw/RKECr1Xi3EuighcKH3l9/ERAudJh5qHWHwBuHJYqSiICPsot2EiGu/SilVfz9laBG1KkD
TusIhgcG3cGwHR7cJ1jp1FsbCgruhwwajw//3b0yV7cShlqbaS0pJLU3oZPtM6m5UMzYm8NYbYXX
DU1Y+SZS1ktICj9sUrr5sXcFFMcqLQcUr+MOB0S+c9DarMOPovqPOOMDsK0ZrC0Wd9Z5bFMnK4AR
InYh5HhOjCjDxvT7F4w4DUq/JD4jc21cxBQhuydTN6kl+XKg3RgtrsUZRm9uJIPVoGRTHVUJTUTB
Oz9N94QTR0Vv9FsT0IaC25dRbZHyMgk9TK54P+6SR5TM2TCA6vosPy69T13qm/NsQv3tCRI2BT7a
1bJGcJJFvea6lTrcg1Qz4vHoWE68EiGwKEET9olcr0He/u5KsHTpCqfxX0auYOp5XwlBKW6o71wx
G4VaQ9SJwY0f+0qEZ+pKcgzGK6PkJQAyv4UpY8c9cLL4TcAWgULKXGBYUoFTl/QGkzPBH/8H9qJF
/s0ewnO6a0RW4JXTdOvhbtN2rmwMCYzrPGe+sngzQqaWOBqJQRMvbGhgSEs1vFBxa9I8ZPaACPN9
+OpNKPyogLcCEP11FjyZOXcrENfL+GJaiQSlBUZSDi7hzmhTsqhhPq68SllWGj3jVJgdJabqP+eG
lXZS2ItIszrK4rIUj+uyf6ns6D6f7H3OiVTolcIvLmaJTe0jFKkJwMBYGuhCnwof4VTFWppOoRLd
o2EbhMaBIRNkeVLo2YVJ0uif3X0uEvTaNDsoykbEL6p9FPPHJyITAkqTnbtpUksRP+T+hNkGiNDB
gAiwaiNX/vxJlZi+gwHtClw3RspsnxEDfYYwq1ixpT02J+ZVYw0aAtapGcz20eGKKJ+9BBRbsmSO
TxQbQ838FdDmxRunB/nBaaGpYxLTomhptTUdPutEIdZZNIz4ghg9J2aIeZvSC4IfTjJ2GHYgjxRp
m7ItNwqJoj3pHGsWQ1xeaaGEtw87cpEQkMKtTqgSSMHtoyVrIm0VbEXvMC4mQetq411l/mcc/vNe
uze1XwSJSBV8XZjpg82gfsiDSltPpVosUJUKBOvHLJaiWNanH3rIPbmu2LhIkz39NzHyhHK03w+5
4KrCoPAZ2FPfAZF3wy8XrIFSjPfZrmLRSnj1o6wKgVWbJfgpU32EKuyzri0LIaOPWY+KZTvf01Tp
OzDjmbHglq5zlVZssBSRok9KnBVkkT4W/JdklBLUftOI2C0gu68RviGP87si17lJz8UIXlvkb9sR
0BOSUwdr0bityqlpA66gPbog92bR+lL0nezLTvWj0YezS0SMu/DsOUT6Q0EBPT2o/1j4jkRxE3Yc
xBTl5ghMZHHEwNM4d0f9Y8VBLZzZli4h1lfCmYuWpWcmxFREM3Gym49QMJKKbyj9kexmYUi6Ckuj
oLZxAfANMX5jUDJu2lGJSBhAfTiSRh4u/Txj+4H1CZX51s0WyEr18ayUAe7DQ9gdyD3cslMgISle
1vHk2D5RNtKtcgyRgZPf9UgtpRYdRKoUVFXm+/akswxmwShxsvCJ/1sfehHwDLaIJckdsVQWMIIr
FnlZIrMtT1jo6bEjZwjBpPWEjH95nFizNEQ0no4osE1L0HCFz7NnmFQGZYn1HdwVVRtwSL28cmcc
FkXObIfNrCEThYukYOLPAkbp5A9ZAFRaEF6rfIukl7/aNUqSGXSONV+ST95kuMnclNnCtAznJX0F
2Eqt5xiBRosU95SfJzTsmArP/BZZxHbvRqboQIyHlDvlaI0Celm6MwxDzVSAYuokOMpbHYCbO5w9
8SrAcV+4xt61xIs1zHdlru0x86i5gAk6O2oCJv40OpStB8eZsbrIWatCrUUVfYxzntXZ7lQBZMzH
+XWulQXVT9kaVlzn9/hOncEZATaPM3W9T+bW1g2PMGEvAeXMymNmTvSRfzkmQHAhnT5cKcVR7AWK
5rSD6gco9vit9uD43g1tVQ4jc5pAzl6rOjSyebHv2lzJEA5+u9l8eep6Kxti5dLxYwLfqLTh+8f0
m88n+TUwYIeOuJ/JAQbTAxO/HyN/6CoHP0iW8iTsNxqcBhYKFxxyO2Q9p15SQ5ar52M2D0Tby7xO
5kfqvsoFJailRAx08szB6ZSDbJrTI+G3qdK4Ujf7rXfOKZrZt24psHI20gJoJLTva4NVmivaviz/
aqxFtFog7n8Fp35yKIOovohXp+FomNT24GNXp2wzRzMkdPY6AbNsPSjFzLg9DVXrz6JpRFp1dfIZ
VBepOg3WZaF5GzvkdCynhZOMnbFblvfmsy9mlKteF91hu60A5xKZGlD1YjggmTzieHmPHxLUqFKE
g2DKIejKAe9WiNMMlNb6rq8d28jfaDRbLbmvhUj5GpknxfH8Q18mVGrw7eR7fPIwsyMGDCCrxwlJ
wSA3VMWhD6cm1ulemmpJvbQU8Q0VM1o0sF+phU1rS5S32cGkrigUAfoncOzilJ+Vd8rUJe0jEXNu
aSFm0Nd3KrRaU0py7LJbiqgyB+ws78Fs3I2qgKijITxx2BkG0konyTcjECxBIYi+iNOEkW63pP18
b0sypLaXvnAICgvxTcECI7JZ8b/n03vrUS60uDvf5L/wnUdNevBJ6nB+Qonq2i096qoC+bdc9pTM
Ag+avfqyX/G+2+1MSFDAV4p5jHraK+gYl6fNDwHXhksZSfygwPq32edS6pOTVKNCuIwNiRF+99+q
04MV1fX3z5w2tqEjqELqC+yIWbLVTmvx6TiZeUeUaeqd++3wqdNb1wpO7chAZSpYRJy2n+vBXhqS
63JPWsArM/UPrBv/EOs2n8l0aEkRKLXlE1rjYj8OEQB/dX+mV5emGRlvmkft3dh4JVDv2JloKOPP
sjeFT5xxy9/r49p0tIRs91GEBqUbYeuzyzLtcdhkUA4iHyVxNiWc51tVCzZqYVYMQASd23B8Ze4f
JBUuXlr+cW6zCJFy2U/Ypa9JeLRNmrBCMD/hPnxmDaNH1lCbQA57pb7Cx550S2wfYdRfCyRZaxxx
VWWCOGQ6DNSsiy7sHvMcG9gdpyoCjleHi0uCEl9o7X9HeLbsTkCcyEnVUUBtRgapZEPODK6Wk8B6
GndueBQbKu1zA63V8hszcArucS5gCz0wjo1Iir35FqK8m6phVvBgt7rXmD4pHZl+ODQKsPauA0XQ
VveiayTrefPcsbVqGj3rDi1uhXkL/iHAHQi+hC5jexj2Ei9Kxwr1kxz75bTHcEuIhGQUtAt78nNg
e+w0BnJ2AhnUkNaE2rlbyED4sn03EhMgHfA5jAaqn0It3uDc9JPodHwxQe/QTjLvsXgryAyx1jC1
U7PYYgEtZ6Zi1GnFrS/RCFRJszryb3uGSKY582UIz4Ep9YpQ2mNoHdxCgXtPddafp3gol/K1hntj
3DniWsMHIcZwGvgzyWv7UV3O3s4Tpze4Lameot6CBRcCilpkYt8VVIwVqqkjTNent2//3Lf1sMl4
eiyCPob8at17RYY3uempY+6+WkGmlTYoxmIobYdLszjVIU4xdfQ/dRPXMWxvZuI5ncdmzidD3vBM
LdtHlRTq3nMWTgYimLOOvTR509ZVWlKlSh/eEqxthOVrroX77mdZq7dX39WUkWcnEgyyA4eALc/0
fjt/nEaA+6tUCq+/w5TZbHZ1/78hAetmCLTO1MZAQqXDBA6ehfVGPRiun/MpBGWRrz6Ujw+mM9yO
xemW7vltoWsDHsNu8mZB5Vh4Nj3gHE/ono8MpjiSVxn/mUPbjQyy6YNma4KEQjtbF2YCfk5BLca+
MOmdTH3h6382zbUzr35rCL6xkLC9stqBxuEcuJa5p/bI+RBQo7kQZDqp5HBr/PryS4FSKr1uV8iT
t3L0ArIaollsath14YJl4pgxB6CSNt7eqhee/BOsfCb5AypkWY9Mr3b4YTQmjMehup2BCDgpU8Dv
RcBcjQ8poibT84ROPrUdE1596e+M2kUoF9AlXIAKeIVO/fJK+ozYt+tWUpX5MGl4DwAU0p9ejMj+
30FT/tp/Fq6zeuOxMPKA2MKlrH6jTxV4tJ4y46VDvAZcpPkM0AWgdysqs1uAU5eUfguRV28lKJ9/
2G5LblJzAQQ12F2/Dk9paNetfBe7Sjm2CA2ZcFb3bTYJqWirxg9R4zPYqwpmNJV2HdkK2v6o3MLi
F15q4m7Y81SRxO+imKn0FJXq9bl6yN33IfUNZkohBzcsqmsZALHZDFy9lNMbupn8fzwhSG+28gsr
LyFWf1xHOP5GqdUq+E/Lix4hemul1hot8v36mEn7xxrdzqcsAdOXXM3buMRo6KUpJRXv0/XlsAVy
8ZkTuHlQf2G/pJYy4I0TbdFQKfbgASa/JT0WM776lc4D59TDlQ4H6IQmTB6TvjuKWK/RjN7iEbKp
KPzb+Q+HeJcx1ZIEfZ3yk0K3fwLdJ/up9W4L7Y7gM7w9nipCDMXJnjgT+TfYfsIzcvexFT/vAsJw
F3YMin8jAGkcJnsGTb1sVTIFMKONVbrPbpS864HZUDXJnoED55G4gZsVYjHYPBf6W8m4WIKjdFiU
uD3T8Qh18+n8oK1Rw9SmIPsMAMGt6XwL7FK/fcbi9llnGG06dS/Ckqsee8Ry3DLF7fr47/K1QNke
Q4tWRTI9HyRbbQyt1uPRVg6E7kaTAtKLqmq1OpXIDcGxfLNHq8PYUVDPcC/uHxQFTfZGwnppmZ5P
nMmC1cfYd6T4COqfRz6HLNW2o1ddcIsPfJJT7khzWLZ3Cz/OHVUPE6Y2YYV9r8DJnf3E+QsUTP6K
oU5ojTfTVsRLO8xXUmIG4yPmj0425h2/2m1B/zBR+Icq5K+pJoQ65LILHv3nUfE81ql5dFPuQspY
TSFPE6aph9hwW0VYd7VSQHSGkNSS54FITg1Gq/HXe0MujDBLIOvFZ327SduOrL+zBJQ7zWG0Vcs1
3bfS5NUfyN/iYKwZFXmLIp1vursy/4md+7bRA12UaKFHdG4bKLxr+azxWR3nWeb6QK3R3Ap2XgWK
T8StTKWjs91TwrpdwAXqDiZ2tD1otQ9a26d9u1RgeBpn//yHAquiR1g3FJ3zPXlK7ZRhUkBD7P/i
rpQUOENbQrnAW9ACx10xo+sljsOCp5/nbGB5PLFR0oywcjDp/ub2DfXUOCwYnoENrlqfF1/epar2
aAaRJ6fyZu72vRttlK/F1/i86yfSti2vGMCxFKRxE/PyjkN81P70Yeiw56v5MS6x6ae0nYx8M/s4
gQkES9hfHEVBRiWSJXpsYQq0ubrcP/2FlUYTBeKaCmQiKfWwINAK+eFFf9T38j/9+AAxCmuOa+u9
eHfO7l9GtUpFkEnjJgSD4kF2KnlB9EjMFdg08yMPIo3/AMr+IhAtJBlRyL2Cvjc941+s9hBu1pT0
yr7V9bv4JH0LEL5gHe8+n4GHLkT+EE5wLkBCcIocsbhPP65TKTDF0TpNEHDOENMeY03vnqFy3+k4
ykYawURNcMP/EHNrpW1Ltv2kR9egolU8SbaLqcCOsR7YK1hBNYaIbgjv2n7hOse2BsXkLpLzOO6j
chnXh0pX3KC6tnTFUl7LUUzLLQvIBQ7C3zIJwCHpdLbtDK+4DiF8mhTO2Dn5FfPb14oODCMoaG96
N+ZugginGOLjFL88RPOW1x7XyFUYmTjSM9vkPn6qZbg1UvDMWtXzYqWhzmrISN8KRtQhczyo6Kxu
qVIYfrB9Xo4FRmq19ehpJ3rl3ByKWZyDVESkHktXpUrav4/ho8DlBIbye+qQTY7DYTorC9nDP8Cp
RwYseF2t9ZH0Vlokqr2uW1jFJ3ifaF/dq/3iV1fn1asQhCEWla6f85CBS5DAODb0zxTa14UFVwAB
d3m7fHgx+X4FeZDe3cCql4RNCkP/18luJsragCicz5E9LhDvD8/xEekVW/xN/fVLCt6BcSy6va4e
KZeJ4gB0HKZMN9C8YTXrPHe2CDlH3fHYnq8FSTauhCJOonMD3TjWzYJE1zwPQk/q2ClaygDUtpZl
qUmBNK+C2TiRxo+9LqutWmgHuGle0I1s1d9DqONEQ02SpgvEmFMnLWJw5QtK4t3YWXMMM/XfinnW
t2vBPh6KxEXXo4psBwmiNuUWG9amHx/Q9fX5+wA7hGuwKmn9usvzHCwRYABN4js55QJQhK/PDrZK
qtqzBDp7nq8gMZAKi3qixCQP9rtEehDNRgNlcU/mz/bU5GKxWlGwQlfwZ8nGdNac2ApK4WpMSrNa
kQDIbK82CiKkeG0lu8GtI6EXtus4n5JDMK3b0A1270rA02KvhVl5pOmZew5poUSmb7RAaIFMsnNO
dhOPMuZabEgtMEPfgHUYNOUOPUyEsMD1V5Ac8hY1sAXWNIe4ud1ejxMer890qPgx8P+cqDZ9LB6d
CDWWAyRfVuQ5sZtYHah6yGa+oE9CzOrHtZBPCZcPtR1SF6qIZxXhcasRXB74+FSHsHQKjENe+SFl
4jLf2KVC2HttPM8oove+2LMps+hEjjRXGDFxiX3/4CiAut/Rbw8FWgBeg3i7GcteNRXPmxxlJMUK
f7AJFiSpH5uoV2zV42vd0JKKpzldxqxJgnKSkTuIk30y6t1qZsVJVGh++gtb8G69G5bhc0zxjusN
8edkB1fdJVYufSCgNp9SCW3j5AmwCpPgpadTjhI0Fr1O03uD4ZhoTyJTNdIwduLYloJ46ch0+25b
F2dthDiKDX1nAySXAfNvWbzp6ejSEOfzJvjKrI/fzjtZvjVBAkDigq2HDGg1uscRJUJsiCpXymth
NJeOhgXwbjBN44RqwwKvcrJxzkv/dXbeyh4E6yqcsSRdVcWgFRZxdXzxQ94SKR/OgJPYs/v3NpQC
hRr+8dXuF/o5nBuq9l7rNqehmdyPUEAnhXqFk5t1P/VvwbxQnNN8LvCu/0z1qNsAre0FKQ/jGmDa
x7VzD02w/CBno/PLoL5Nai5GI/iV+0doGVodC7ZD0YdkFKFnzNJMKT6PMpu2n8i2ovi8669zhJCx
qGgJQVvhWiFFCdKrg87fsSM4wif7BnyewRiOr6YLHUOO0t1K2UFz1v082DUm9PRT/94D/uClJsdw
tZG4NN9DFS6Z/AmqLzp4xuQy/DAmkJEH3T6XoZAaROVbyTV3GcgT7TeXzmSMErsso1C0cpSTJHgN
IBMOAM5IVTsG0rX00BoMLf01L0pIZY73ABOFVARKOP/DT4lFYqcWS52er680D9sCirBbYmKW6aU2
FgNZ8fn75ezte6cIHAkRDitr26hE2IFwjffKdZ2/okJM3rtAxuAZaJgF7tjAm/GMn8uh3Xe1urVA
awLIc/t6GVi4+cuUFfTMNbBKRMwtYN3NV5LrngjzRp9+YN2JjMJwUj5aaq8dtDPn6WSR3LvlNw71
KTTe9VOamImbl2MKWDeAgNOT4USrGnHpgEYR/e+tysk+rlGNvAceRuOSGZv8FKOXqsiCSEQUjV9k
GnbF4nl7RVMC92fo6NkAhOBmgDQSySBjZD+vS3f3qu92wFCeudyELJw3EmM+cIkc8abO9KsUDUHf
xJMpQSw6TbCB7wu8eyI2vYPO1rE4XFN5cJMgGePhGQOU3ZrpeT9+Vihz1CpjCNXg429uXFGL/V7F
bVSU1OJGkEBPMyFsaj6n8t/jwkPZKgv97cbS5tikDVkTZGAYLQT8XXWy2GbMogfpB/ezeMXPcROY
whBsAtKrQeTIru1Qb4+2pzrUGCmfvSRcIuonh3Su4rdV3S0qEkbZvCoMDXmitNdw0elLTu6uAV1S
stDMtKHaC/Vl+ADCKvuonedl8FrBl98GNKVO8sUab/dfUusQhs561z8ClIwTGHaL5lYA0weus3KC
sMfm3avkf96tmtaUyTO7WTyms9qpHudPbdmvY4Dk9Xdt/Syp/diJYkVYvuhI27Jwu63m6qDAEB6n
SlKbRcP0DLtM325XdPzYg7hp7k57Jat07z5hb4K0rdsxONTNxfLOuYZ89sfPCnblPWA71D3veq6V
iYrkcnd8WaCqFHrz87gAW8lG/+RhBBJiyX4cYI4m/XpD3BW1Vn/F5o/M9l5+AoaKUIvFYf+7686D
ToBuBaivWcbc3nGll+KSjB3YuwA20SQ045zdypHrqdW2Bd67dEPylY6xCbOHG3Rj/KW6SjFzGqXc
0St5vMhV94dOKZHp53Nr+I7qqXlAJTJBG+yiXt2AFyDWqooZHJ+HS/sz3vMuE7NZuIs/m2MUewPe
+3z0Fu7jORy4Fg7nOJxHLMyIaG4K0V7zK2aoWKvJOTMfTH3oFyEyJsSehnKKrdupMSq5pa5Lu8Vm
sSKGKO2ZK+qXUz5ER5jXeSNakaCBzHsTPCHLH0TfTjohXM382gExiOmj6D36HHWXu2JADuPigFG5
OOE2WkRZSBw8slqzRkGbZSk/dw5JPPc/lH1aF64EYDuP3CMiAmbnPol7Rpl+l3JdVFNhxM7juw50
C4+voqnYc2k9FsiH6JK03uoobeQKSM7+ESxtBFCI8syvOW0cuoiL97omt+C8iVtFkr6Cj1ST8mey
caAxU6XR8WioVZBSwVXGNaV7Jc8P6A/obUcXVxjQnqXUkNKTujA0c6/cq7YV6Y9K0LwVOqkmu9n5
uRzNct+8tnyTab4+mGi+7X/Wabj6bnr/SsIIySQLzX51v5NaxHkSQiia4SV2Jxh4HhbpOg3/v2pA
FjoL+bT0UUoAWa3dszzczmKsRlnifHe+OZ/EFjQGDXtZN9ItbkyXqFY6eIAZnMK4hw+BcP0W+DL9
Et1vl4O0RX95ATb0JPUvi8z+cxP0iwy9OP3LlINidetmu4YjBnOjK32cXy+TNUX/HkozqT7yAj4R
unF3sX44+DmCLMBHjwbeQAhjMd/53dv8pgvgj58dcudJyzX+UokuReCIu4C/cKg06in2F7tdShSb
eAJdijnIXDLwY+yisKR2DDnOy6kxqqptgAJ0dN4L3m7Nh0icyXVrrCyo+Ilkz8E3NV2gdlQxKzEM
jGrkHSX2HSDwwIMKs07UV5hFxPzpeNlsBglEScTNZQV4Ug9nNja5LVRGtTajRKz2k/AWbaS5X2Oj
Ao1zG4RyZOttjCYOawuEdSgiJik4kKEtg3gIhw0oAfGGn35s14JbZx8W+htHE/uQRj4ihzc5Xos5
cqKW5ko1KjTAY42jAQ1Odrh7ZSqIwbm4lSPqdbkO+o+XzKsV9otL5BFUUIbeJFLSCQGF8vxE1IEL
o00bNAiP46IK9hajbm3GXi/dUlHuWrdTZ0PtRYWm+itMkcddpFOoIr9KRlFBKf6MbJugQDSCR3KE
PS597iLDOUMM4vmtKEsCegFN4FcZWQOU8WNB70wWZF/4pC4npRWROzAu+/mrNCK79YkZmwlNzhIJ
6L1jK5ARbDKP+I3AcfW3GxAtr8yrAglLnDwtqc9EYEtfnYmyr45aIcqhuh+3lrSx5WGbOXDkA3/R
xm4WxPPCRKQ07jgttQje4GSPQPSZyT4vFpqgCcwA3N6l8hwiVlFkOLcU+Xf7NTGBbrdP3dH/VsTs
ZtgJU8CRqwUNozmWrYy3RVqcTfUSCv623gDP4qRcWiBb85e4oB3mmzaxa+JeF0Roq5B8mmltJRUp
LuP/YkMVqPIN0JMWtK8QsDe4sEuTLsabuOwyjrcL47qy8Tf/2M3hPuM8zoSdz0HHIs5Hn5nnOCZ2
fmuKYV6ZMimVZaNY/OA0SN9f1t7tVXOEIIMQ0Zi/muPlE+65tp6D/tVw1Yrt+TN7H0mD1+OpBplW
m7sM5ZntqhmOFTVR3mvy4dUKzzbkbMHTeCJ7rrtfhHZ8oce5Hqu0sL0RiPJoPycVwMS2M36zsyAu
HyS0nI6F25aD0eJXsAGiqmRWCots7GTOljOmqzbvIe4oKdQgLcF0dVGiP8UoqKyCFGQ0qPfnW9vq
23Xkpm19+fxfYj1JaFSzOd+5L1ME/E2wgpg+AvmH5awrtlpAfAyp2Q7Wl38pA731LD9T4xqQARID
1Tl4IQ4nLlnn/cvBOd9rlrRytDehdGnKZS9IOt/ZQBIvpd8Xoi51yeH8RAEfaj5spePJylvXysR4
lXVCPf6SOoTFrj57MZHXWHAj7Qi/s5vtKtF7dbs2WcovzlmY+1WLyQIiVm/CZSX5RAF79yxoob30
wh4u8utDTx6842F4vFeYzjC11gub6AcB1B1Zb67/cwtb6GK0o9+ozdWaYDWBcE/53IAh6k/kw90q
VgeWWYeBu/EalubWL1KtpAaGZr8xslDHxzVQ0ra24F5s5Z/If7uhTWvfknpsK8t0UXuUnRxtFnD2
scq1ZyAtklXWoCNCcYgphh72NxGhriYXatjoTK5WvNejpMahJiYbWscO9VzkFZzs+nwohY934JlT
OI5H4z/HO63sBip6EuTs3UIMfcv5AcF0bOx3v7G3yQtKW/aMEbpbVW6fYaerc9fq7JNGkvUj5Fm1
h2i6DwvuvyzbQSMGT6aN3NmjHWbW6/fyqwGo7Y5YbudegBzOgTAcyEU2G76diZ0aIVknIRgskrlW
ZGwkTgMKeyXS98QRC5+IPj+yiGqr7WfcPFXZyxpOakMCHPSsXUMEvtPimgbwodQIhKzkhLeSRy5N
1VJPPs4nz6Li1CYBnLzh1XcDWBFEg0uTdTL4l5VqzFI/wNRTx3iTJsQ4Vx/umj7ck46q3NDnfLN/
nLHQqOGul2nVRvoCP8fz2cqyWHahBbR69klZnqNHUYfr64tdvbnANumviWzWDw4FVkdHCrF7Xah5
EshmkNSDoo4OTTUJImvAGK5pscYbfwEgf3/p2sKVnsxumarGxWGuFytGuP+ECkmRmKFYEHA7Qj9k
IqPm/KRa/DBWUWjOGKJjazurrgB0qFUg8v7MTEAj6fB7nMqapqf1sAaxPZfDd8N5CazpWb1rKG1n
Tj2t5jCNsLONiwGUFrO9uPMVkaVNLKRGBDUImAqMgc+TqIfHzQ8R45UPysFTpKGZJBQOlLamHGjT
aXx/WHKluM5TfI83ew31y2lI4kj/tQlSWO38GTabU9nzJNefbSv8WIxF83r6Mw2UqZlu8vRnkz7c
o37bB8daI7s3WT3OxH418JZJwWKV95hfbYO6aI1sGmIQVcU7ifFO1Trx0aqdfVTaFJmIuJ5LgbbL
gnViKo1ygociEZ+gJ+qp54yVk4XeQXHIBNbNF7/aEopm2755ogunoW1LBueB0K2Q0MLF3fg7wC2s
+Fx11Vuj6U+EI0pe1iPd5iexL60BWnpKku8bXKnjQxaZqKAwmHsHdyo4C7nCFjDptlHa+Uaf+3H/
QarYYC9h0wylYQlnLwfrxmsIQ2AkrB/bxIkAhNx15pJm5t1gViTMyrdl45c5nY+RbUixza/4mUFX
3/lTZE2Li67FL7KiI3MZ9iBqSYsxPR2LxhpmuIl1NvkEzh2SN6ut6TKAMk1rVWY0l1b9I0ZkPPqh
h9UpxpVSEe4Ro2zp48w+UAi1MgKSP1z3rNLY5I5cy89eEdl45adG7vrS8tjjqD1oHoDDccnFmLJm
ttLYaDmIUSvNIgY9VPvHAkxVRwiIUhFJURZR8vwd9IX9yIH9hS2g6cTfkUmdrOv747DLDknThI3a
m3dm3de5NcNmS8iZgqO0x7HJ+deKc/VIorUr3Wrwss4Z7K7E7uWuWY+YJDikO8olwUJaCFA+8Fsy
ExD+CZxX4BIGEF07pdBb7G8/n9FJvR6wTwsr9BADdOyIUAW2kd9hR+DfsdP3WQ2yEedC1cW01gsj
vY+K2liz+cdoeEIBLnqFS9wpByYzLRnhgGxHUMN926ylvRV5LKYJTdAcBQ2Mbs/ichlNdA0n/roh
TzY1A/ACVFNdKDqprEHcsRJVN1jA6icRF3ozW9188ETP0A2yHmHi/kk2xjQ+g3A9neuvTkQLIMLL
d9kRYhTGPjpFzDhDea0xT3/y/isRFq56vf4+GhV9f7490ll3WaHp4PGfUFk6Fid9xtO5ntphKOxM
kWzSSkhHcF3s37SvNawmyVqhMeFWHwS636W3j2vujryuxuD/5iwvaqRGETOXCru2204kxPFjPQPb
olOhu9piUDG/UELN9NfAwGfS0Q3zU5We3+PGplH11tDmB/9AffCTB+u9nWMHdnJMB8rV+vnga2hL
stRqdcrUAuvfeEyzQC14grjTaKl+aSIfzfHdxq1YM02AtTf2lFdjoY4KooOaO1NAgmLhO9yOOE0d
tOmIGt2V5f7wesfogGCqYekc1d0QBEhtuAH5geXuDe6jyyHrTtC/mG+Rc4Tq8uLS2crXH7sMaW1N
M5Gs5fbcf5df1gNpY3tQesHAOKAU5sObwSeHlPQrZ4R6IX5aHsjmIAhkSyP4Xco0kZRaKi3JyQyL
ZDYyteyFJg4N3Nqe2OvH+H9aHByjXwXskcDhrI273vSphP4bYWpOXSZEpXeO1gC05NQ6cKBzwSAS
Zpa8BUcg9umdrnmPy6dTtpdtdXsbFnMJabK4gmg+Ld9rmMJrn/FHJLRTZnaXGMTYyuImcRChGrQm
pHxRFSR7I36jeX4e2YxyyfO1uY9oedKhY5j7/E76OgLCpxPc7Mnbuf3sU1z8d6RJNObyV+hdPKf0
C2xs0QEi7X29IoWam4iV+c2WgcR6auxcwLpgrdyEuxVUSLtMJBUUFHOYlKY3V2OUgs3KHN0nv6PL
qbvtrSSBxDkqLtYCvv83RdaIShSvvccc2qn8rBwd7OuvogoYmxiNG1e1Vd/jC9Xpr1LnRKnb+yK4
xVv2mUbq1U0sZOTJRUVB44jkT/KMBcWLITTGPro81M52WgwiaZJp+aHJpC2OC1DjO2eVENLI5RJg
ZZT7sQTQh4KBTQKh/WvH0HemczFoWHN9ZYm4td9X/mizhD2Pl7z7Z3oPppvyacowd1sqETtcWJcg
qm9GHTSA3666fOtPGTOr11pZmi2RLPF020csK+C+CpKSbtAT6r/XqYMj4Xii8qAGYsaqClNKkzKh
dXEqzume+wD+3iRC9lKSqZe5biE3C4vIpUMwBpoZugC3qXuehVhk20VWdZf07XXRqiTFX41f6BYX
ZsW0iIohudHbrDuiuMR/B78WLLqxcRUF67yVBVcm2b48suC22kRQtPsF0wLT8nxKusfgyb4HPH7i
bPuSbar3sO1ObIO0nDupOR5OPsnNP03ciK4xfDsM41I3wdLQR/PGU8TEcZsqmWfFRuN5KjowJScW
ZyjOJ+T91u/cYV3abZF+qVtSuK3S0k3KcLbmR5aORyJTsKd9h+DRMBCN37ahew8HrCPCA2Y4qmpz
IPS77rbo65NJmSu/4EDpsg1ouds7W1xeFWc4hx9UI6YdRk9Go9wX5iOJX1TNG4cI2ld87MdCeqbF
TPlgAOABCozIQWTluwU+r7pjGl8yHfUxiE0AJMPXoAOtSa33Eec61lSVf1u+DM16A6O4gtjf3+7u
nbJEM6LTuSBYhPau4Koc+nu1k47+p8MIALLt71n615cU9tQRo9R+5RDQvljzEDuSsuYg9houLnr0
xxVJoZd7hP3zMnhlizObL40QRcNQQcURllyBC8bWSW8xGRmXAMW5Hdv7eY85UywH6vnVaJ2rGO4R
JYa5h+Q1ZkwRyGSuOfRBzLU2HbjUgklIu9E8NvAoe441tCaCSo6TGuI/MUauaqiXrFZBTo+xwO+i
fZou+mKQ37ocXTWKRZVDhOu4g9TfIJrxJBfXGl+uVXSZqRkNOzM3tIkiWdCyVh5RI3LgWe7p5CML
jfOE9FHJOoXzM6e9j5tDlILFd3k2bFz84Jq6zseTkacclt/HkkTCiKeAZt52WrjaOK7YC7TvS4mK
wO2DkOu6oGE4+SwQ+tpy9VHPEdKJ2uCg9NgZLSdXLxFvXmAcQ4gf1YOU0ZHw9ojfdyNAlNxDJgOI
vHQvZ5VFTky/4AptH7Yg+n16ArDZz9oJ07VrqEB116wLi5yQ0GQsfU/Q0oWxEWcRy60SJjB4jgeE
K1bBoYnFgpY5f9MfTbgqtkCp/Igukz0baeStGqpQdpRMAnLi6oKELf/VsPVLKf51OCyhVBX975C4
9z/CbN1Q1Z15lI+Lkr9ZtLiPKNxEvoPFb7bdWCoIjnITRMVKltR0yLOMr8Tu33D8Q1eeBRAyuFZr
Fw071fHhEV9lBJbkx4bYqUQJiAovA6ncYtRZZpxmaJhSXaLs8W69hUw1w4oTqUQsXFBdJnxq3+Rw
7soq7GxSABxyFxzIvUXwDB2+JKrAOuGZ0Cja1WwRTcD5vY74qilymvophrZgyBg6ZHBUAgm20vbG
ECuAmjQPg6+LjSro7f+5V+7DM0HBdrPQB6APogjXO8ZuGY/IZQTRE8fhkr8tL5ACA31HI0zEUSB+
JyZpZu3BSO2uCltpCTcmhXviebPnZJhTU+tbJZdM21q1ul5KkDStnY0r2Kl1speZKMh9gXs+eRrG
o/pMtXGb+uElP+meqLO7RxKn/fdZ/x//zXocfFqe7cfqzCnR7cd1IyBVUOk8fOpFooIa1TN6Y3vW
3AvBZr1v9RAOVxVrIWqV/EU4JpnuBvJR+zy//SA8lUcI0agrQ6R5JHbCbEYip1lFy94bRKdNwSiS
dCAe2pz6toaxhM2Xrg3FvQh2eeFpWrfZsXB8RxBKbmtcoEsUFtbsSReKcElMGqK50/ZQNp7NaSe5
CsfWpvyldOHwnSzAr530gv36sMBOfCeqV+qgh2C2LFSkDn3LTPjL53VFBJOlNqzLznThYFMGVhVz
1RUhEolKZkGe+ai5UAK0OBi0GcYJSZx1XkMJX0sYoJ4eQbe2HpfIokiF/5Br6yWgSVtF6hStk8GD
pzMFf4oPtP8xbXvDUHFx2mzH5pidtX+0C7MkWgmsaBLOz8ljUMM9A9gLVmF6jBCq8wnsUAu+8sV0
7TH3xBBaWCqpYCk0lsztdf3Xhr6a+vLEkaA+nsEHgAJwxqWD95mY+iGn+b8wyfiFHG4aQiUxqqVh
OXfCFE4RD5GnfC/cchwlnN+pbCJlYQyH/j9MlgR/rrbmNBiPVMhUID5kDGHKW6SRf/+D72BViFoA
pG2bi5lfvnXMC7xzuUyRhqdB8xidnjiW5itcZAsIMM4+s8MD8dhlNqMcGiKHBgtnZHn0sXV7RXes
2vC6weDbiHWP9X2suO2xhsRirq7Ln8gkEw31efpP9q+KkWOpmCjLc7u7TaXQVd0+H+THfepU6eKB
EhRE61UlAqq02PW4jm11JLSJ8k3ocFKykWVYzPZzANZIkx2U+eJtRgmFkfbh7TFwh5QaDRpfvG9V
chEiXIpUsQueNUP+OZWXbKO2U2S5yuKJ9EmsKQvPLScqbbah3QawWnLyaYXJQBYA0OO2pD2OUypA
Y5pF/WzswZp0x1hWalvnB5bqTmgAZtlwYHb6/rKpNmh66anXxEC6f0Lxlwe/k/USCIOTnTbuhWwy
UC5R0M4HUEA/OM4O3+hZesMuIRY5ry9nsDidCGRWMhGKJPL2qD9DWklF0mRYgSnEIuhbmqTPapjo
jQ4/D0pst2DvASO8GTETtrVTNa6Ma1sSWUkkM37c03r8xfF7H83w6BazMJobOdrylDUsy3+BvJvH
1D2PVC28gegtxtWbcwGUWY4C17z8xcr2+7YqArY7Y/p+XCJ75pmrLx8S5mcbrtOpFwypYW5xRMBm
FniX2Lj3X9hDhdrTtNbQY1jXvixhjrSTYZ4mRx1yin00eI9c8NMUbQjAzLUBPFQmPdaushFhF8LS
81ySrIdQ0Il1e/RBrzBkJPgp4iflFoYROt2aDbcWivlGgT1eyuRylgmdBa8BPARSTwN8cxyfw9ty
rEvt+nd3n4XA7/0obZWk7Jahv4JDxNT0G9M4pJUUHJtU9DFf9H6vB1aHeZFIHBbn4sR7r8RY4N3Q
ThHYXWRFB2UWIuADf+rH2ULdpBwXdMK/CDaYf3iKA17rKSyevTuJLMTa67Xgk2SpHPMPU2ZF5+Fr
1X7tESUYAZLGRS2yhQiLGY80lqmIBp3Rn4XB78m4oxW3bDjaNGSukKv94/kx3ykEl31Oca3iQ/m8
kmvnDGJJxX/+cPBiRo5eGPGBvagljqT4+lirAfb4HrIMWgnvY1/08m3vyju+5lBvBQFzeXbgbHKx
PmkAwRZK1zKtyIG5YbUAXczP8+ULTJjLChq6PhzeNjRWqBZk2nP18q01PEWlZ83TkrLOn/rc1OQX
0MIEykTMaRH5jAHjpwbuk+JrU/KZ8c32hHxv7RLxQMxchShGIDorwzwqMNflNs+djeVn5R4lEIjm
gIz9z/S/lCagkCIGNogmXG+vciKDNAXQZLBO/LlIo+z8/7/qZPNxrHIIGQ8cZg7MxR3xfbwF2YTW
CQE/OzQTthwzvQcILmfV2dZU9V4/p889jQ3cq8jq0yUXe1Erfa13Cx1QAamFRQOus75mRAAWq5OQ
5iI2MvLhIDet/YJUkanMVyC88/svvneeo5dj1i8wbNP3cGFed8MgdHyMF35BDkcORq5DyLoxhbns
0sgniT3bMacWqWVRCL5ZWUbSU01E0k6iUmiMCriFpO9w7hcROoR1hDyjIrQrqxBzfRwAUGBJ8V7r
uWamjiB3WzJxQc3iMqM/wxBZS+swggKVT2DrPYMjvZQuBj62FkTE7ejkdSwQm6msHvM9Bb+y/mD3
sro256S69SgL1gDrgzMlMyLI3clleVg37ExbOsoMFprinwW0prO8F/N2r0SYZ3Or/1WaDtfTAm+e
tavYl97HNcOeW9x3ZJAX0Y1uf8Ew3T9/AmDaOcMXHLYmXm1qE3i7V70DvNPUPDMA7ck4ax8Uq5jl
C7KBrgvfar9AVEr6F1GGS2BtNgvanTHHxUxNtDRA5AOWsKMXQQWV2zCLf/jzTA8WeaKrGWgA9Kkt
rT/zgdlg/45zlXQCKGikSGejbnJyZBP/F58hqUR4au4/5lXLV0gEVL7dREf51VAlRQWKCSY9xRPP
CY03FOOt7ePZfSpN3ZY9nvf6nO1akk9ekAzCDgp+nDBXurpV0vgq8xDsHA9mJ0yXTWMk3AIUD4UU
gImHpKHyc1PTPQPvdAJbMdHWrVW6Gca7x5vyEsH3p2aPCWCPOjK5HM06TwANENO/fPvD7ARQiIp6
wIwSjSeWDsaR171zAMswMHA4IXa8RwDztWp5j7T3YOacSBn4ARtLk55jPZcgGhhvLdSqdbQhUbc/
FbIoDxTvIbfOCCbLtzXCK8Y3q5XwK+W7dUXPQTCwm5LHnS9eIgjOhPhtBsQgkBiIm+ijW+mciJf9
SFvAg56LW0thX/D4rfUzG8N0IFYNYvfERf6JbqlzVniVQzRMFScOtQ3ChE70b8AACa6R25Z1/wBn
sgf7I2OmwEErWqlD5Tozxv67yli5gIuksIkLGuQLmOr/rTzJRF7yynvT+XNNmLLo42EVR8J2WkfC
b4yTX8WAdUJwl+iSmvepQcz8oiM3sJ/mAvUBvsfFoLe7N2m3xO/ypTe1zIhoO70pU5mDmXR/Qhhw
GBD3G2taeee46DlfVkqVf8Pk/0ZdjSdMsnkrpmZ7qBKfn5Qv+mlItr/XLxcI1TA6Ia4eqDClCfXk
mXTBwFcJVQYdcGhYeh6gKn3Zi9IN9JwQJokZiEodOGAkrLsihIdzCWRoKWr+qUKRrFfoq5pdXpfa
rAYUcuplyatU+SU8Rz1tfq477yy5IechpJxJywwgTX4Oq9olUJkqceIatnJR1gi8eZn6ZG8JODD/
2M22gXz9QCIqY1hHbavg1E9XM94zNjAszwqMJhNtt8T7Lyt4UgU9UxhrfLPB4YZdBSeiyghT3b3z
sBP+EFUp7faD14972/Gfh4iVcvggFs7Dc8zM+fyto1ilzVFmhqDH0d0+Fw5xE8ht8kWMXqZKJAEP
d+gCjKr0D4xcUx27K72Ga38qAbfpdDiTti+snY98tbY9ZXZaXbZ7yE4DIPxiCb37ldm+YTY5sqUL
15b6Iz3hJh4eIunw7bHqG3g08Vsljaeh+tsg40UGOBUHhxSC1DGTJEm8FFKfMmdI40+TddtzvWdh
NhC6B+vyXTq5L688YPijNeQ1bgQckc1XX1G15+zNswwR3np6Sa6RgGfH/kaj+zayWRMRAD2Z9gI/
oGKgfZj7pPkUUVU1xq89luIc4FwEkqBBnx1APjL4tPelEA40n6imkJJgmgUJ2FDDalmJDnjoHu3s
D3xHYOtTAowog7wYLXl5XQkxU/PipTc1dGBSx+J0o9VE1Sz2h+A8yYuTYV6g1OUjsMBAqwhzUjrY
uVWt+T+f1rf351ZpyH4SVaHh86jt6qfyI/cvxPxJhXYyL0sA1DV8UYO0Q44UDYbkFM2t7XumLHpS
t7QgGAdCmWmqIMFs+Ya7mqHzlT3kuENHYbrbRJQdUmSyJKLwOREr9T9bG2dpZKf6bIY3sseVn14X
TdwClHG8hFPoMtw8SbkqiNXiS8Mdebfl1pQ1GwuhkfmTpPfb7RFvUhTOvxbOMhPRVm322IbNnajx
rDbJPBXm5KT0nei8rVQhv1Os7OlcI2uJHV4Stb4eLhSEtoQPFVYdIQn1HAxT1WnQ6uj9/vRAMAkT
BdhU3mDYMDfRUAsgvuZKnP7JdPWpiv22XKtE4MWFbnza8pfnAKHffNOCRx0zQm3+tb2Q2tYwpJt9
ESmpHQZ2vLGOUpjZUtO4ncathYoiTD0I6Awp2iv7CIddZFIxd4+/7G05Vzpe2uioIOD4eTuhotHo
llpsEQCD893AuUv13A0GWAql4CCzoN5NysNF30aiakRw1S5XjOkE4iTeej4b46D+LSQA11PS+4cn
t1rDr2fb7DpTLFFuFxa0tHnIPhc5mYQCYrDAAI1DJQQCAa2gpIDpW5LP4cIJhmgrmRO93TffPgCp
6iW3RbZIZjEir2r5ST4y8u3WnzmpLLV/l6zWIK9Ly/hFHEfHIDHbJ1ooVQcejF3J5NccEPUa4iBx
tqBoq8nqqCCI1AC3ESz9oKdI4ToVTMYbZMEZJZUtL5WG4vlT80TcUJ2BOmY2AYhIULB+wubQTzYe
q3mAFBYgGPf6w5PkbTeMBmSvf9kG0BzXjsKWFTDN2PI3p1Ic8LfZjUTTqXVpVao5E7F5tfj1n1VF
sOFc2fRDPhnpCy/oNZFK3liilVaUu6JkW+MvipHrW29ntYnViUAVq8Sl2LU709cQx/YExcwRwHB/
JsvpgoOdRvqUUk2CNtZMdZTsm+iX7VCypVPwHSIMb8/4Gn9MlYJNwWXTwCDMjnDZJxCj7hBktgOA
l+DYZ8Civ2qaEcpprcwIExES5PIlbS0kBe9t4ov66cezgjWxJoKDAHYQovdjc18HCuCBX3aFenmw
+BMfwvM6828Ym5nYHxllQyIECsauixYi/Hk8/Illr+UZQjttQUmV+sAkw8liDhXdu+Mv05DcbpYT
LRtXG6aJf0Ze49/FIDs7GVDPV+Cw1yJBRhmbM8hWlf5CzcuCC9i69z0dFa5pwXpKBjMV4HC8mdvJ
DoIDcaqs8dAl5vIkurCvqGusJrlWsGwZ8hEThobFfwIHtLG4DULCjjOTkSE1KMW9RCGpMS9uY3AD
9/dmMpagroPCWYFnwN+vcmhd99ntBiozjaNSdcvwA0aAChkFMBTSm6shqLrqH/LKQVTMhB/Cz4MB
vDa+F4wD01TLwS/EQbquaLFtCEw+E4vNwr9998Bcj15xNwsZo06w2+jfRGE/SldVWS5ZNnbiKhyI
/RjYTRYHvZCjiyyMBZJRw4FMFd/qvIRpb6HjVvi26mRTBCuv48c4+6B0f/MHkYHYgvd60oQK+958
sh91qTtOAO1S2F26Xqt8AXcVzHsDfrT7kGvnPRKmgo1lK2JTZCFpoiw0eInPZd2cMn00JwTR9omW
RVYWpD5CvJM66IZBccoEIX2wlMgbjFn+WtBYtrhAVo+BTJj7VrNsx3UcYgMoPVHt0B6zDwLhMFL3
hz7hY+Ph5KgDZQX4WXMefu9YDJhE/t31RwX3ildHIeMQLlr4EwfN3NLeQTLjAGdn7VtsLUKUaDg7
uw+b3XwGol23QKtZmjz8p7ERBFFG22bZg0D55jSqc+hujkzh4yPiQgRkl5KWnMaiHGyQHMNVs0+F
0oTBigcMRcU6IqEaVCf/H0FmJ8rrYjcJ7UNOH6M6ZV34nUl+eIsYAlfNj/3M1/UiKKo/k5kkkm0F
EXREmwVrcXcx+LPd0oGwAmILUs8JCepT7DUX+xlXr2K+R/NowsrRsFQ3zv+tG60mJHHPVvXQym4O
yRyKVWdEFJVGWw1Dhwz/Hifr+X12nNMUt5LJ6w4UD/fg1FAqm1CQ7hiBi9SwRTumJ5q+4L26XI66
Ydt9B2RcvQOhtzFB8UHvfJszzuhHracKjfYS5CtaenSCjjtuQeaNgTzPlR/cAGF4GiBscNkEUSrT
jNkOtAC6Wn0gs7lhGZ2nw4EQxUNuhezEr+PFkdwPGJJCFmcy/EO6OeelLzrWPFOvv+BZ9UL8TOJy
8ND5LXm8bAF5w+WtI99qzg62gRsjkPlTs3b5JhnLyaJFum+HlQoVp/ydcDSsAxZTdGSTohKQUH/h
L8mnu+SC1ggVYZ7WvRQ+7q3M9m7OSihFcfBwF7lOntIwHpEPs7SjWVfT9pk4E3Lzh7GHs9uO9vyO
2NJBInPBhd63TtVE5VUHiRoA0GJw8A8KS5Bn0yVm8WSJvsAyQHFE/6BD6fqdfi00LzdKz/3igXwu
AjZCZr/wCs1ugoCXEhV+8+JDTyQZ/ZjcSchRb+xPOsmNHgLeGVa6P4eQJT96KXCnmR9oCAtAQR5s
UZlyq8wEBnpIbtzxNcK50CZ6f8kNuAkZodx1+6UkMOqCN7+sQC9D99diRwaWSG/J8dvdFvu7PzvB
fz5ECkObAGxzaL58eih3e9eQPgTTZeS1PP4FpsJyNp7+kc2ni9Q3a0niYDWGJJl2s/Yj9zWA6UYm
B1GaB9RGcOLdTVGzy89DqHXjpJH3Y4V7BgOaRzt01U+xEGRZjHasca0SgTUqHzwVSpoMhebnM0t9
z3+/8AEOMUY0zXLR8H+Br9U9DYnqpcK3kQKu17fwyhxnZpJ8mSE5BrhgNox2IxkZKV5iYCj5sBrh
/OM/E5ehiclTs8b2bZzzXR3OnbzK7WKmqILK9E6+dDzrrterv6yWp8U+UDRDskTv0UXwT2TOWEFT
8xaKA7q2SIsx6y3AvSgT0Vt/PonevAPbMRGJwtttPzsO2VUY41CRXlUHLRakie2Y6BguohIYSigM
yYxeJ+/1yzr25eRsE76pVE6tTJmf3nsH3omuPJ1y55k9cvX15QcEqXGQplqOMdYCAV98CMhy061C
38HjT9nq7iFewXOn5FiRaZV24hPXMviY0XITe3pXvvnOgPLzHgU7z4zpyWzjfF5KHZlE+eoMctog
AMkp61OaUN+W0AcShFbQHAKc4HLfWS5ALm35Vjdnw8Le1xXhKAuY3unZr3S3CRdj7kDrSwak3Aj3
kUGVol+qTWLPyaE5jR1Vi93I2x9vERTMmsHxIk06MrhP9SYb3bXUzC377Opv/DTlGS5nyU4Y3pTf
OWRhBucmSrFO9v0ELTbCFerbZhEDim/J0k9kItLpkNCi5tObSZU5+DdnQs9ZM3nYEOz1H9FeH0/M
NbyV7ouLRKZvDyLiIHTN45fOujK1bOdWD9ABWnkboirRa9MBb9z5PkESnlDOUfs4WvF2EDBCl/3o
Pr/c+OraFp6usy7WKUCuC4pBa/ti2LLwAf0WfeR7xK2VEKpDI6zqf+VIILuwY3xf8eLapIVHnaBF
msntKpSmVOq7ZzddClvCfOEAo1Ruk9HGNALVlhnPpXdaP4vcbfKZEPzxkBKkDBpR0hHPY/2hLN0+
EBvlcrPWcZg2OHMFYjJo4NJxWAR8E9e5HLERkXfhLQ6t0pEZk8lLVJkAMuhazlyphbC+pzclQAN9
5PfxvLwYHGDO4DeLBXQt74gp6j81+zD3HAslPcec0WhykF2LftcD708KnNmBW1gqCIe+et1InqFh
JJ0wRq8pUwpwdEPVanieByGkJIt/RVIC1AtIVgP2DtS7Im2dvpYr1mESv28Wv0N4qPmJyEQSqmfv
zFZvsTemHN60amSEvc4XGMKCmYlF6KVpQRnNv9hbHg8TTHSKNSMBQdsZ266PFlEWBvRdh8/hHGL4
XXhxta6XS8HWOp98OVr5AH1E1IUo/z7KNK1tTgVedT3ueKzB5hQg0Wj+ueFMX4Sh5sgSPd37Y5Ez
YoJV2bAvzZMM92MSH8r+IBiQhx2078RFMIo7M4y6CHkkJn0ucClyBudqraR6uuZU3VfmBmcEfS+f
aWcoQgcSfry1Z13dKmOCdrl/PJfUKl9YlZTxqQPO4kZ994P6nyMD+2O+qc1B3IR3eaf1UBGfXiEr
yVtYtFTcgBPqTuCesQpLoj77rJRBUJj9KfoRaBKoJjjGknpIPz2s5SiwXmN4w1XbdPANMdFst7nl
2V5ISNqdQP258a66xc/CLMpW5zH0dfbOqvGdKDV5r3fuPDPH0j/a9dLpriBaSxzB8VyeyrplYWpd
kMtmhkgK9MIAXxHAId7huUG/uHv9rG7Z3RcdlgSqpgCh799g99Yzb4iGmu5zcue+buK9Znw4s0RU
vybcMd94qrbV2hON1d7vVkUKrHNgeWl1o47qBF3J75mxljurEm62UODGJpcJaoZYWGmFHLdGSAUn
Yew9EmCA/oEfPkLNdcH7rspUrvqIqV4YKeJPFvC++ti9CvgroI7+So457TMmdrDGNp5AawAcW/bR
UZ7wu74rRaLyxVN7Otxe4av8c2qDZQAGRXFScMMMIADrcV5MPu1Qd6m+SbInSwGS5jrXtqd+HiRP
noqvINno7GhSHD0XRWjBdaELbpGE1dgMhpeI4vxQOgED6Plmvu28pKG87PCpb6OZIm75ESmcLL7y
7K0GJlr0D2WCD0xtiwZOe+QEjZVfR5wQTiaWeOhJ5jKRhFc6X0a6yMuTbpPgMQaOQ/kOYMMADuQ/
pSl58BEeRnwVDIm5QLKG09xlpV4m9F2iobGs9/bu42nCqlCmuVQSl0MLWSBK0AZ5CMGbhWtmiQC4
+d5Xbp8SNP7wG4GnkWWxwtOI2yKAKsnacxv1YltduIogkWrUWGoj/gxAQJkbD48nZiHSvUOJo464
2ozO2NqNrWvYvKwVJAOluhdKzooW/hfDXB1zJf7ueRLR+gkcBm439dYoV5fdOFoQXg8AtDiOENRn
4ebrdi2nfk2mJRocdidJtv4AHsY8NJGxheoaCfAwt8ajGQi8b0hhYns+vPrNq/XFU5otlqs68/Ay
tfLPHmW5e2sSdOSQOh+AnGMxtdUk/UUq6kOEBOVG3aPhMjBximbsV2xXbYSMKPx8S4L4KNadmSvz
DVGAO3vyudPj4N1YimwDKe45fphSAsd+Tp+Qo+kqobrk42zPVbhb9LOE+ZhF/mpWy/oChiLVL5b4
rHvkgsztsznMyXOx7Gx2vz+KTCo8BpODDcKRBWixNgSKY5smHgDJgj2Ia3RDu6N0wdqDQuSJmaQA
dfMh9LL53LT4qvH0mjNa9FU2A0SL71fyPDQhnIWPRq5E48p7bDB8D9gfdBIjJ9WO8GMMVUtFnZld
cS6ORhb1w33Z+cg/nr6ERGvRUvvF1se5Y44Ebk1O9dy1FrsCwB5SYeFkLhZcpQW7cO5ysPEvDDt1
Eyf6mlpi2yLd9lBNHDVs8csIig0lq5N13+p/OLh5b8Zabup3k+vuJ5JIK5snEjifpjPu7DdAI8yH
VxP6stXKu479pziGjE958L5rjuJVrh1IUxGkOOWUOZENjtBTP0T+V8MOOE7qWlCohM5KfZ4GhJC7
fgCG7WSxmM8x2ttHJRcY1DQBESWFo+n5Vs8uusGs+tuIU0KukqZsJ+gUQglT4idKUivJGHzXbhX+
MM2IaSSetpfSt7+/hh1j5olAW//1IJP1hAXDZQ80FiEdslFPUFyj6hb9t+CRNdvXjkEzM/2YgmHZ
Nnkwde703k9QcWMmwNO2GVlzvBxkzbWdKnbQxVngdw9tbGDgwIPZeHOpoJmtxf5uqxR/oYjaceig
zrA1xTZ7J7M0JBgJ0kQKYMiMGVcRxGR8a4a+OC2wcSi1EOm6r1dFvtmnPnruU2srhz4JQOt8rrHf
fhnoTSjlOlXD1OdEFVvLddr+LyqnY3Q2TH/Tp3V+Gve0c77ZCy24hZg673K4+uLEseIvjM+qHvlM
H2kZ+syMERgev01VT8eBeqtROIG7yv3pkLW/RuLbZ4hD9bX2AEvYq9Yi7aokI9sP86/FFtaUgreV
l/NGx1I2Z2qa+t3hfmYJBHhzeHKJwJTgfOrSK4lcthigRQSMFDuG7hARvkXrr6rk4u8bEY8/Xucv
28+7rGXo2jE2obrSREhAj1ZCUcX3Vp+eCeLsbmuUJN4awDHaFg8dYdAJMZh/atMcqC/b+fV/kuqk
h827/INpvQ2WsDQUY6bx4Z5g8AuawembVyMf25cX4I5m92BNYPrOZNwiGraOikTeC0VsJfHbagRB
bU3+ULoq5TidqOlipFIjIdDQBRwIddZAPAyrJ1lUZe5WaOSwrS/a5SYeaJXhi2U0b4rIYV3C9yRh
3s7B/grPSxqObKtifrSKW58HwCLVGJh08PToWn8PqaFbGW0ZT8SwQEJZzU6MkOVXZcnCZR1woss5
HBJX3nlyo0XFOCjcgXk25cHVt+E99VAlTsjP40nGtBAZPXNbBMTYF3rg6mtlyXEobfa/pV5cdgyj
LbxiOwnPn0CO/Za0k4gCfQ4i+vWHFDgKf9mh93mc11D5IV0RNJwyrQjEfctG1YVG+kcfiYoPQgHN
QXlUvB5hp2Dxz2EJU1w/NPGac38nyIEbMVbmLNJQp+mg1JzguJ036Abv5uDkWGm3lgFWmtUjeCwK
OylWhBlm77ddIjhW6SOzRpwIcwIwp1BKb70/gF+XEki5tk97kilC0NXAqInASAJNhRyZFOQGGmPm
VD8Se6XDQPi/3hAAO4MrHGzXqaYYcDVhwpj/aKUaL1smzq1B9Gy6A1bCSBgMpQOVuc04wcJsYOD/
cLHt328Ze8mVDzjCuNzIN/q72B8ki//ktVlVrls8mGfUCOTg7hfhLZUZMvnMEAbcTG3kFEP4id/p
JCQ+YsXPeVhuyUcmNgG6FFKECn+0c1pvjdfZ3mtkw2921MtygYgo/G7vtin8ToWh9ISUVpXR3E9v
ZGeW6NioPKlExsaNC418nfo8iSg+rU8WuwDLJjVpHVwhRQj94GqZ7eLd3L+c2cnpHF7t8bww1lDU
edrnrHykeMzmuz46u6sgkGt+R3avzRMapdFwMesQ6owH3v7/TrIDNBZteRHN+6qRqodA5Zlg5+s6
/rKpnhSUw9zcptpEjB9sUIyTZp+KRp/TjEIpaL2PGBz79tm0br+WobHu34u9feoGXaQRR2fHl58r
rngiOetIINPDkUz5KH4tTHmihjVvgKpj8GF9EF6Ukkr2KIO5Xe0H2eqnt50j6kdk2KLcEwrSN8V1
VXhLdwVXSypAB/DakIuYT1x021o5ybbqsLyBOJ5TP//aKIa2nIQmaBP8W+T2fx+HcoaUX7Unae9o
4fyO571ey8vICh981/RQmUnNXdOtXE4XtPmUIrIZK1mU8+gg4Dxy4C4VJeDO+fRm2M3Rm4glU7Ns
2t9Pxiyl+7mBnV3cohP2XTM1qz1N+Gw01CwufKvmoq+5wd7OsjRmy0ZWW068TMvq9b8ChhQD1i6w
7bFjMRXOH3xd0HAAeYIBwcutgcJNpkn08yjtgfWIYs2s7hUkpRVXf+yad967KZJSif6T3f8tO0Zc
KriFX7GJ22Rkv+lfiFSqnL/2BkQRCYX6q9mM8JQQi7dqw3XrQTIS+9ljq8DsUiSfNqVNLv4BCRNU
J3lUC6/eGy29ozBg82fNAuncU1E2g/c4CB6cih067iwwWm1ttTklMztqUAEKzSgeUbvhS/AV50s4
2Tzop9W7fqklrIAdp8M65nRQME0X1jvsjsjItPliy8HxsgFtxeyOBY4Af+JQ8LPkjJwi0DuvvJnM
CckiERE3mHnONJjolEOdj1gMd5TNxwEqgB4V2OvaYgxdlm10KM8t5KWfpkvqEO1AjFTeAsDq8QyR
SaZbKQP/8Z5BeKFpKUOrpxNlkBfJlPYpF0lZvqMrxnotafiEMq9o2vTt9PM9RAxhF+xgoioYyF5w
bi9j0FojXNqJALFUZrD2DigJFYdDaqxtE5t4Xi6TlO2AlWHoUv5YWe8P20+eFG9vYSZ6kG8yJHTS
p6VnFGERTjG5QD63dkQoZ5lQ7xfxb61nI7Z9pY7JA012adksoPZ6N36o6Hugu6Hx2ob0QjuKG+xG
WK88SeIwsqubh8Dl5twSB36cD/JxxeHbjfWSj/FhLDPngKt89abx1qU1FD+VaLTsFxSx0U9RQ4A/
QNP0pw/pD/uX/5jkbHoLq5YvqxVksqvH5E4IhR6ZRGoM9cwaR3tT3QIN2Io611PgVoRLxWM68sQ6
sZTWaZmiEpdAAmB7cCp93/38eNr6qY/JrDzLJnCV17mggtohIoIPkWyguMVV0XfN6UDw7sWN8k2M
knlel/zSQd0lR4UkNpedAa0GPvZXd+UuIqw86okNQO72HhaFC3bx1jnRVhJtFDzZ/ugblOLwE4Am
Wjqca6jP+hZNMncMNVB1vRawS/UurwUruoB/MVrloLh8rxl5w+xB1fz1vBm1nDy/PGTBnZvZu4ro
HBqoLuSSaV0IVSj+PQkH0y/w3QLAuV8oPpqhz8d6tAcHLxONJx1uYogcZP00EJ+fcP3zZs4I8FRW
rW3shqmLuIYWQFUOkCPffvzBgt66XT8Bj+SxMYrnoyAV+YJVkg3nYEnDvKmcudchgIPOJ0k3K9Dq
NsTL46Dw0RWaswy9LM1F/K9Tr45uK26mwDbR1wypHsYzkRtyUmZZr8jl1snlRnQfc/y8xRfv0ArA
0dp0cBOBb7oTW2Mwjfi5W0y8eZ3c+DIR2nrDJztm9SXdv6r2C/VqU91ZqtZki9u17vK+gSUo4S0T
ig+g2wG3sqMJfof1MPVQiDbNLJtYRJmZMzls3FsWcbdVe5+vzxAh79stJiwlNZrvKf3b6vGVQbTk
hA40R8dIumrH7ukdGg560R/vsABdaBOYsyhEi20aBYgNpk3nYSyvPwhCfq/n3GH8sSiwO3k6C6vP
OoJVQ1PxTl42bvuF/tOowzJicWeLX99ynuCgD2kS+4er2tMrNQsDpr2+GpdvvMVphiadaOOWmW1g
zhCeWHuxRAAXFsL7QWLEEBwwgY7NOL8v9PUcsa7v9sLIsm/xLSJPJkF4+H7wGZh0/0jXCZNNzWml
0hEjuL62KVcCHYQycARTQxHlcUAPTXmUXyz/9BupB1WRU0ppek1inM8wp6YIn9f8v8WzsY5bRAJl
fMoimWhdg0OvSsJW2RD95h7Z/+FhzeO6UkKnXF6OwL3t8xd+EyvX0vuK+nIx3Z57Yrf6QmocAxFU
TPrvvPRsrt4OlmihYtgSMX4Mw1mAfxfZpatz/xOost4vvvW/SRn73bHwH+9KZvgYFgf6Bsyg/AR5
rP8GfYLqLEGtduo7R4J2fJajU9TR81hV8JRseJgsbxpxO3K1VnsjDaHUKiLM7b7behjSUHI3pbMi
HGZ6mQOwv9cx0nKZ3UQAmaJ2Nqv6VFUVakVFgkMtzIBq2u7049fO0Ry8uzJ6FkuCedn5wzienXMV
ljyVTYD+tt1kBej14E5dkMI6FHCMKoSmbOkuECVXYyx5Bu/HToe/U/1YTtvyHThr8iYLNooDp7QA
gRJmlK5HSkIpzvJ8A9wIdE8TUEFPXR7BBT05MvuCGHdVxOjhS5a/1QuGx6CG37q6YFr9kZFuTfOw
lPn04mKDNWgOEL61flYvzCLtjNH4f0v3UVg+PHG7TdxniAg4TB2+FB0wrDR8OE5c8WaBXZL/b9KH
wvEaJ+9inJUErDoDO7c5jhjiuwB0oIlT1u1j7qDCai9kJEsSh+hNBADb0N1HSt0+xEY3K+E3kSBL
Hse2HJlR49j7a5blkX1CMEupyaOiQZUnFSJS4RPmqRTcgR9X1qeu/NqXh7tnUUlWZwT3y+rqKHXZ
1CT2JsWckI2r+vDPgiTIC3rjxW8dpcNqyCVJqPDjOLLWOqcJNy2hcjv2veDPuLJ8IDG/0vkIQ4Mt
UqpozwjAtW4aziCT8qqMniRl3Z6jld67G6Ek1kcn+vxpJ/aW8XDCLVAu01T1xanxjoBEXdZkcSgS
HyKco/85ybLSjjAzNU0AZ7x8chNcoGYDd2D1zfhK8ggZhtGqUrWbChYpuElZOmP10LYV93mA3EhD
IEjFGTXFS+WCPTeNcB/edjG8fjS48CwBSZxS4r92Cp4F98g58EKqtJN0T7rirDoKUQ4CzN7ojBJo
XKEykTg+qsjh3aPJPsC+SXeXH3G7iHStJRrUzhugdy4yrjD8Z1R9h8X5WkMCNqKDRc279Rz2BSLf
AyjJzwXpb0b4ITR7+OJb2J1tXn4ZUbhtuDu81jWs6xiCLwS3qs3yGCvfvKVgBn2C8bmxFTjcjkPW
D2oDQ/isTuz12lDe7Q0RdFcSTl0iYA4m1xZzUgkNtuSOyxxVRS17nenzdrqwRD5DT87dlLdlomEt
Bnpw6MTJcFFc1w00/ViUbGG3vRdt7ZbkB6ruXg9HOjQ6+uHAgpKa+Nrm1j4IWvO5lCc3uLv571dI
q/MzRSfaSfdAg4DKnEkF1Agt0K0EaTHrskWLTpLNL5ZRqnC9WvOUC5fW1UcQ6tli4aWYJrf6To/M
j0/AAw9Wf2JPrOeGiSvrOv3pONZvzF0HlEq6IvFh5dw5EsZJxCbiVmCJc7gm+3HBimUw1gitZStf
gJ+nT4wwK9YU861HHvBllczQPbsNhVTszK8FayjX0i6ZBb++VQh8zPETWQss+/mENlbZkiEyY7+r
XAIxJS8SCqVyKNNmgOkMVCydrRW2MfnMudPndxcEXmeY95gxNhMup/POfGYV7iZQ1gYCB8kMGYrY
rDsdRxEJwsclpAa3SL3H4IDB0oY5FF4D2NVWrbOT4i3jGLj4HN+DYrr0sZ9D9C5hUwhWc1Psi+4o
cJmXqwDFjrCiuzPuPxHGnE5A/44y5XGxVQ8nHx0icUHrJDjeld1y/1klG6V4G5zBnFxq+eKER9aw
Ev4ILca1nO+qfNRP+L9Lmp8G2pIjcFuV72h5W6O6jzonTJodCVBHRED2usL2lYCF/aWa1MoOsUI2
bkTYY04JaxkAovllsKMAi99txkkApUP5eXAOXC3tt/M5/GtVznH8ScIWkmYw6F0KIMkOqG3U/DFa
QHWZoZ7fDrVgQsZ0TNCcTab/Y9DP6p5TU+ba8HmgR5PamMdUe1jrNHQxwRz79xOtVhFnTeEdaMmF
6cl+FfH2Yhov1+2qaqELpNDPe6xB4G00ZNrrWyy7/91HGSxsJz9R9dqH29DZ1IAOsIsY2WUh+86R
CtDJRd0xYdnaZpHDvNiIxeX18As83kB1D9n71FO8qIGRc7eLJu9ciegybOi+sxGuH4Fvo+hX/PDd
OycWgt5BCYJ7SYUXxUxFx/9aRYF2R+TpHgqRZh0oulL4aTNFSGrN2SdcDkxUpVffpVsXte6sXXu8
LxYKReEY6MpFOneTbSRlyPmfxgtQGq2u7cjPhaAxg1m11dCYLhI7tCifCWpfSENSreN1r2JHIEUb
Hma+Jl/YR0+qSldYjQSfl9yo+DIvXuF6XXHsaolZJ0uRkBav228v1FK9wiZdgsO6LpTVcOPVJBqj
EcWlqZTxZJ/2Sy1yX6x+k5sOHimLIoVc1bR3IeeIjc32w1mSuK8VxKOiCNaCFXtjSU1Wj09rxlre
FlI4ru8XsYiwKTZClwj2zVYQI2AcLXWdSCq/iZNyD7vXp536tfOmyI804wy60kTM42YOOVaXWbHU
fn8qIUCV1wjJKQ08mK2jjORmLe7h7lqHPm5bsMIc2/lcrgrMmNwI62WFPqKnUSU00vjktAdspzIH
LFMQ/zUSCA6C7WJhE0zagcOg/pjqOHLoFQoV/ITXxI37thnojojefcWPBZqXgQHEqXwSL8h9Dg3f
hOkU6c6WbeY648jZD6CgIpiADJKNsCwk5F5+l2IfPGT1Z4POiA9PW7fCjkotS5qaDIGNeDuK2zu1
rKgPJ7vIDeirA4AbqaFetioGQRVEfgW10/DfeuA43my/D+XLZ4SCFbm/cvaBidhNT4a3ET+RJR6r
H3Np/2yI26SQfsD7v1AddOnG/xqzcybRsvID72Bk4gdk2gTqvWGNWPC9jvhdoY7ejt6ipogXGZlQ
vLVDqbixuVZYHCg8dy2zLJvw17qFJkn3UhRN2fUd6CQSxR+K1et0Y3Jn0em/2Sf1/cFLpro1ttjF
Ux7w9qRrmJlDSZP0POfspJqQxdE4y3FtRsMCf+bSbQGlpwQlSHK790GV2ux8GH7tLvlcCK3+9fhc
5zRIjYR/gFwPGHnqkvuS/Kde+dQz3/xQwNhm6WAzAnlFN/mQtvZSoO/qVdiGi1rszSGw0vwc3q7C
SUxl/RqESBnMPURUHyPVmaIIB33eu1sRt0wHvG3556KMBYWjYSAGU44r3bf12uFErqTqV/Q1vWvH
FYOPVuR9W5lSm6/ikXsbecMG7ln/DcfjbiVgYaFBXuxt52ao+FsB+T7Z3C6WoRhN3oWj7qgVpEr4
flMPP/EGumTfvPsddmBN2125+gBqRf2cm5lqpGVj+ZUa9bAXMiafhkV9Efof9LKJvAicpe2axaAP
N0unELTcT1tf0h6V/Mg2GmcQW0IT6ZV3xbDtWQPuXnGitP+lxqz3pOJnupcfiIcy+KmLiFHKz9Ly
EMAppLHq7r/vrgHrqMf6vTTlWsvdvP57/w871hIyarWIJrMIOHWEcj9oAf1ShgeXuDXmw14gIIPV
Phvn51BOivwpam9C5aj0Gu7hNVSZIqBmDIUeaQDSKD74gxnNP9dPpA2ZpMDKBLF7VIqTxMG1wjrA
uTa6rwcplxvrYC5ilfVo84R+9ZVbjheEPSjIHW6ecPKFN5YwpV4b/PUMxyYxfHqZ852ILuwIwMef
uwplIevDOlpwSMccU2bFD4fz6k87oBuS1omECd7V+5aKVhQyRkOUym3TTwD81zYRDKvwtJu2Q0Rj
upfWCdsFXwU1j0BB/PetQjdzIX8qAELcsbMpJqL6sB70WYXpj4BW4XDciWd0ANYG8MQZz+jI6P9Z
+SupPXwhiyGYJYyAr11+5/7XZnHSPL39yIhNjb+pxM2Svc++uAzQuz2gFT6pX8aQH2Kb5WyMf7RJ
ns8X5VyoQ1l19FqIPZuhn0f21+BJb2FIhBdjuY0e5/khE2mJhDlnBKEZK2b/zKrfXNH8qA/+ASEw
ysMz0oNhbK7lKUhhxAbbUABELN0RyAm589IudwzbtYFqu8xbWdEHTO7rWFgw+rRV1d+N4ud2ZfSq
tJAlcLYkQ7KuG7Js3Rav4gKLQSEGqh7Wfe3Yt6NoNd/tbqgQkV/I9wR52sGQNxqqt7k72Kfu4iXt
qW8YzBD4rFikKGouu0UwNz3nFRDKcMBX5jjlMjhG7iGdMMVeJBuaPIinMcZxoZa+dtxclcj4miyN
FHWgtsQZp5Uke6fjvniIEr7HgmAg/mflM7yfLBHm8jQ1bAkQwRY1+gjFUpOcV7+fGRLnNAD9+Za4
Gi3xpBBrn8nIPOoN05Mzl/oaezDEXCX7iLdRbNkOgK9GvJWgfC6Jgod7lGJg3CP61Bf9pQlpb9sh
ETp24CuEYMk4/uHpgM9tkJ6615w/T8gwEFyeCXx7IUv33mWPktn7MIIV6uegk9XmwoE0jQaokGyJ
7/tC3K9NXTOF5im7wFmshE7LsCytvQW3KMQjc2jLFalspVSgLb9iEC4jf4cJf3eTOrJhcDWB/xEV
b61azLSacZwFiEUNbLbu44FtA5FIV7N0dx9gfSV1yWb2wHNFag0B+tB7uoS7ioNXCnq4QaNh93xW
3hJXHCRCIaZUpc8v87RTX4XBm7zsguCIlto/GZVcqY90EBPm/IbFwyGacQDQAMqyx7ZaNQbqwVGY
eh4li+sjJBFcyaESY2P/XEIuxQa3ArJYrLjoLBLNPELtKap18yhPM0b7P8F9RelMDWdCljmT75vi
KCICzQGvBRjZpBFKDGEWAdSTzzu1mAFZkaGeDIFWCPHjSqS5mWe2Xtciun9VHXkrOqUsfihl4zeQ
d67MF0ezIV82jIQH+A039Uu6amG/ZRq2LNFl0l4bCMAGyph1gVXBF2Pw5Engn3CFK1xGaW6yXrcz
kKfi9iS4y5SjMPhUqGLThTUtXIg2CZwzUqWCRD/q7DNo39HOyj5XpPVlykWdx8wNHPRmz2qzckGp
0nvs1MibCFZYKyLAeDaDMD66fTjjMN9BOuc+w7BPWliZzI7XnYZcZROp6wwLy5dO+4NcnHkTBh7X
QXSmhVfTN46VJCGzE3IaSIfIk76FUPfC6jifTrOsJBlC01b9GOZ40hWaeULKGYgskJMLgxD/P/iR
3ro3ZXolxGMBV5dQ11lQINjZcZTd1HabnY+/0/dXNtYPXIp9OMVqnWxRw4W0zFd0JVlEeJSvsWOl
WE38/ki704dQVr/S2gVDNiNmc11a8fpH6b8AEZu/URw5e7RQab7cJCWzqAlUXW+on2vmv4a4eGnl
j9mMJCtlnwo8JwBs7lukBgo5BQ6+KZ2OE/TOSaD/CTiQHJ1eVSdaakn8kFnw7utntiG+h3KQ4AZl
IHxYT3wzZl86JoPLJdiqOoGwH9GU5SRwK94gmQIarevmHi5NwNgsme2RnBmPB5+3WKx1UZfuHA48
YFx7Wbbw0Qailyi9skMdSmicG+/XSDVG02UZ+pjqFboSrDVlEQ+Kq4wucg/mALpjWW9Pje3BXYho
sF9LsD6n/+RdksmKejYe5JX5FBY1QwVM757wQG6phSUQ7UnOKn3kqTGOUDRBLWHFP/bJ0wG01gXi
CQVbdYVclYKF8AtJKv4X6VUUshYhpUEo3ZDNVVREbBot7lnNAN7AsaSPdaajTpL2XMLul2mUbbMD
2IBMxyTofaLwfuaFz4kKw6HQG5crkukWdT2M3OGKHspwYEOC5iLZW6B1ksc1TDUGZMRDYiQTYTw6
VIhXIqt7NRd9unfqDyfyN2hYQImeaN9aXPdiyzVX9KFSlscuolruOyq6u5QOBCswG/K7KwHtq0Ko
cQ3RtFJ3tvzcOQQ/gxtBymcfH4DDJScb1TzPSMkFKAs16ZScsPIo4QaqNZjLVzp0EgBq3LZmUJfO
CmNNa1gKm3US0Txyw+/f6B6hSFss+B3rgGwc+iHQF3LRRPiA5up9v2d8kZAJm9bFOoLnQmqDto0h
qKX+k1rKTX5ebBWZk+NALnnEFGtVOBDSrvdo8fZAA4jK5tmBx6cC0e6pahJLG/091lwZU5CGGWIf
TLv5i9F6BXh1QMdmT5KT5Kr9ubzMFlZcDpCMp4ECUY89J6lGo4yEvLv+a4SFUKdJ8EM02aUSGZtg
CJCzekRQrt2beI59bI+mhIWmLc0JASymuNPY03f1VEdqCp9iqkxUMHZJpBletWzFPHDgLkj8OmhF
hETM6T3ePj59KCoIOdqrBWk9ziKaXSNN0EPAW3hRGUwQanWOGoBOVOwqoTRHTSlZk7mbLwlVGa/1
t9W2fa1J+FjTIfY5xEivlJAoEx82zK5ps48+5QuIt2y4VtPrDm+pwa7/Xt/521M2EWJm4R8V9ZDS
gyhBO0+FTysMNjqWIuc6hMeh6zP9MmlsVrWLLVTLW5PIbDRmHczyUIkV3Ag4t6SfHGOxxzrBrTjm
Iug9i0AYi8oCzLDYiN5HLWLxdG2XREUgbb5KAbR0NxgGJtQQjQ6/dXHqhFHfhZs1JgnjjjxCbk8X
/GopVTKzKaOsT6fy+QvXXdMWsd8EqlNVvgGzYMHWJBNmPmD1VYd8DlMG/2gcOtJsIwUvflRCC6m8
QfmqY6aTERKINFWKK8gKaA9zXRUcXwrCuhDQM9J13c4LvQV1+3jqh8FWUTrATNYXFFWUoJPl04pd
HR88gZSc+YiuXD3N57GNbApsjhQfxef+eZYAAZiu0Sow8cxmBeu7UbaG7/oyyewxUa2sAPHH1gtw
hAHh6Hcbznl/T4MVfjYgDtbULC6I8a8bCPlSRmFbpsuxe4ssDo1o/dVedxm3PM6yTCRx7NwxB91Y
SSuruRipBlmzleWYROXpLI8Y+zp1Q3MMxJ1ZJA3r8k6GnTvhZrW4DPm5FbE579w6w8/KHdZNS++d
dDToxI7hUU9ZmzwCT2pHHEvUh02vlTQQyTkGPmsqeNCSVSvM24ckyKwfXhTgNO2D32W1lN1fKtA7
13K8IDUPlFWZdZ46OL3Ae0TkwwxhFAKmQqvs/M9KOnwmZw14nN9hwHgrNzIfbQprbgimnn0HZd1Z
+iFk/Q9kXGZzrKeAQQNqaS1Uj+DVbZci1VFhGI/kP8iVf3Tu+op5tbLXO7y2FKbjL5gqMYlTV1UD
nLjMZToQA7J3r9H9BzBV5jEQLP7shQB42vjvmm2RVHW7m7NJtgyYZdIwsm7GvfAXin5eFx3J87NM
7lcvfYnT2IBm9aJgGKKrYkmLCWdakieREq4wd2Va+A/AO9VdfaI4DDeioLjhB9LuvJ6B+Mwrkd/K
uxOGrXQixfvp6oqD7mlGbGFNFyDQ2vjmEgyXu5PUQ8RlHicsxHbhsKWE9zxp3QPPu4P85afL4gfC
aXTVxtb4MnISmdG0irw/ng/0XOgaQ+oMCkHXqRTExG4iVMdEuUqMUimgM28eSl4cFceb4slW15iX
dozIDVq1NJndqT8d+2dB5ShVAXkwMD9HOcdMTIu4P4XpUxmXjalQ14R10fDZYa57xruzJVGd/ATe
Nbhi2PKgsguEXFdfJJ4qcl+Xsi5MwtEL5C9QZ5TVghPbHANxUKw5uQXyqkDxbmOlCjRU8kTiFYig
r+KeMUqbxtdh5KVd0rNBkEKj5IJLvZEQ95A9z9y+vG1aWUhd55GfnN5BFK7ai6FQy2COqYcMBjcd
iUI+G3ScRVitLtfjPTG7Q2RLq24+/HU5eUvYaHtEttj1ymVlbMAaGHOh5OElFmEDIm32VUVoR27+
8S+9uEgajT0KReHpXZbnHZMl1VZxRpZ1dEGCvdthqrz5OYtvKbT4N/RAGFnIZ5OunY2L7HPHT2g0
ozZY5zOp30zyOIxWZX//6JnTgmhWAhtrTtZXAUAuPjEtX1Cw9vpEKQv957WiTE0Y2mzhj3zzgi2o
vLUHvhl1T0atpxIJHZRB6RsNvCfk14LKkN8ttmWhMTwTHRFNPD69UvNz64TIofl2ZjOPkocoeGbP
F/xBD7cMe3j71imT+Wa1Rs/FZ0AxMhqze+s5SmF0waeKbnm9u86PzCM/tEsLfEH6eDVjOSpUii2v
n7KqMDbBX2cBm3o3bqBZVQ2rplQhhqP83cdfTh8ljVldxrafmC8HsShIJJVwqO966fgmFjPDKPtt
mxb+vNGfS6mFOrX+SqSK1a5DfjBFLojkUc1hlX8mlKbxHQh4eGi2Yfcf9j/WIK53yQRoutkhTM/u
b4WKl/PtBc3PXrkipradvwvK42qJv+fgwRAcdp4t+fAcy01QcQEwiF0lzcJHzQoh5WycMRiN69yN
9XhqA8V4oRUcbBTimOuIBzfoWdhb1Mr33rZJiyqtwlKo5tlZWZYyKGpLphXHjkx1uRlSCEKFgOxD
97WRP3p0MDYKhKdcmrL5VNQLYgIolzgrL2EJckEK5vEy+BI+eY/W3qpEgaXvND8Mu79Al3KKslYa
OjoNj8ejD2vBMA8k007kBoWbqQLFGwRx1R0XH13z1OJ/qzEAbKT1jPRUs59SovLFKdU1aX8I3mcA
oeQsUPcEqD8KOQ7R5Isv/5Q7U+fj+rXsACRFl4YSvjVmrrw7siMcdLhvAvQWZOc4mqzCuQkgnw+L
8WkGSJqbfP3/4Em4yQFgx13LYOHg3AHOmOwJEatPGJohCt77uPXNBYc6ouekcltss67wULrnpRqU
e+1pLwsJSIfRxDhb7BnmhyQveqQJaI2uCLRthc4x2XDGR+Cr1utlYH8wtJArK21zqTCUYW94+jgI
8dRxuCShCMrEzEyQmdEMl3G1hxqHbAazw4BrFiGtVGkiTOrXGpIeqSo5PkNjq5pWjRRrHZt6Y5bW
R9ENElO4PSm7rqqZppaq6Pg0M+agQNgko3YE/lBjj+2QC+yOs77uNxpmMlj7Il6FE4yYBEPW9USu
D/9YPRfPQvtVQUULFpxzMtu7i5Mz0h4KMlH2qW8LNuIji/CecjS7sjJA+jIW2rQT0NS83kOTgTUA
4gyVpKPSRvIfMusxGX4+BOB8GiGSt2sYwbb54rEP2riYDBejMWmxxB2vc3exvSxiaQ2/lUVE4L0h
9M8kvcd2bUFk3Rwbia8l/uKP6xVgBtX9Xqsi3wJwlv/WI/ONQ6xDX1smBjSyDAZ/bH5aNOlrTWmD
fG9XCwwyhZrolSiFLjZONHmPBNQEMn73bba1AJOasWfQbdLWymLyVBLktKpJqfseDkslr3sCh9Pz
8J0TJ4en8lagHEpcoY3DTdo50XLTmexS+b6mFj3t0LY1o52SdCtMcoriEg7CtrGH3wt1xpFdFml0
+ch3gO81Tzb14raG7ePi1N4/9jw3HcdfKdG/QfhmMe96dDXvRGTziTd0oMILFDbsivawZFYmSXW/
rfTnfwco3n5S7z++icripBFDpde7wc5jH2WLRoeXZTA1C2+YYTUYSjT1tmuKE3hv7RTXQlhBDkXn
/Sj20qvLHSkgKl56STQIeIJcvz4gwTeZgqYFSrbSNJUJ7HYPJAY+nSm8Bje836h2/VTLM4QqVxae
rDlLbY00uJSRxShRwWWjG4v9QtWTSsIlRAZnjVV3K0rIRFxkKyKkWGsgm1Prx31WWqotAJ/uJfdY
RlAgA6XEyUBDIoTfIuGv/N5Z2mwVnq/t/68piPofK3qGkSeXzYcch1UyKugX2LMVvssaZBVXg1e4
cveBhEr3taBCOxm6KQCZyaddjtm7oi3s4wMeQcyXF/90lh2eIu3JsnIfO581nTIVEhMml98e9LDW
2sO1Y6A8Lbwv8Lkg8fAnv3pATiSpOn6i3eDBJ/GzQjYZfvsRaJ5CSEn5bNf3OlDKWKzBa4U7mEuN
NxX8uGTPU674vXqJw88ZmCqwr2igkQKOKkJYUCuA3nC/9pIgxCgOh94ak66Lx30LZPb8PQTWoY6y
yid/p6FbjQxa+83oAvelRlCCJQ/wxcOShATDNXZdV6Ta9iBikJVZV/AFoeKFfu/rIcSDr6oNUE6/
qZlJAjrbWNRuh9Fo/OvHXtB1HX2UNK7F9qTgG6I1wZjrcATqzHvI+BZx3aT3skBqRGq7ddi0iQ92
O6+GYBYnVtpmxDg0MQYoCURcfOo51Szr3tJQsKLdNKn5d8vpobNxer6pLooXVrrQd4PRqUQC2upu
ytVA2eS94uyfkEqX9vHrbQHFvih9WqYVpMicvr8n+Tud4MWTHNHEo4YOgmb4iRj4r6n+Tz/+G7CF
70soU5eXQCNVQ4Dx9iY4yd+siULeF2dXPpszyEExm8W32CMG6+1l5i5IJJkkejAinWEOWs5Hbc/I
MNDVZCAprb86HnVQSC5/0krl2FzrBIy6UyBaRPTBaVSo45a4qZDg0Pg+R0fySUyQsvVZoV+BCUSw
4IFnBZWPh2w2Tm+Jsv2dYvEzRiuiGGMJ6lHsTO0A9VztaDHadnia45pcQfBEge58KwjaQPI2giJ/
vivEEw8ngHAI9oqPFqhfQCFRaMDXmaspmnQsxPRI7l3pDw+THwcRUB+Ixs7dUnx/FWGvBcxA93Jh
gSIr7sdUbBu5k44MSflJ3Kaeg1T5EYLEUXe0FQzM1YRI53MFCR6scC8ipd0JOXdayS4ZEtNSM8Zr
LO36fclQes0vOmyJbQ4xE9reScEZLWobvmq70vI0ZQVQJPGTdfRn/DkMs4y6WdNhrJG1wbQjx+v8
Qed0iJL1JXFwhppSmXZbUJ79YtwXLobPF7+0AO41R7v2A0NNLICCMtPjoIfh4OWj9ywTmt3xkXr7
DKErGjJppNJ6WkqgtkBrm6w7QNteS5FTF/Vpv8TuZ2pWfPzE6LueDYYFU2W8h2n1CNNjRXtfZR7g
D6V82RmDt0i1/fZf6c02NafKZb+QdD+XOE+3W3CAI9xIl3eFFSdOXeU+Em0i4lWn7e/BcWHcjLFR
Tdjzop3Yz85C3YWBqKDprZ5AqU8uBz3BWEzTTFuTmi937HDBrZAF04NFCW1OwIoubRwrhNmonbd/
C2SIJLc7cKJjsvnA+tWeKjwJuExllRDBYvQ3cxwrTBnxiWxslWMU8BM7Jk9rwgIDtQyeLdedtD8H
R0zw2A7Za+OTcnQThLdHj52sOam6H1XUg5finphFs4L5e1QDETZyC3BN2WfawVGYPosNtJPi3d+I
Q8XA+E/Mekssg0xj1atrNN+BAWIry0zLgTJTKFHgQZn+GYOLuBiN8AAplYgpK0oHgOVY88IwN6pw
gED+tAgyrPZd8dGDMUCrdLYe9XugPv0NzptLrjHNE4JeKHKsJTMrz1gSRdohj6kKtXuM2WhndApv
+MBCGlbgcwRv64l5FlKYcNtY4zdoqceXgtTqHth5/pv1j1EHwmcLGF3voKBrLPqbGIwPnXUxN/X/
DaXglWIuaa+JPy55BdXjwuTt7T8Tl8rh3nMfpwpOWwy3LzCK2XWVkeImy8CRfHyNTXzfV4wtiGKK
ooPY/iLpVy/z2hn8HgGNtDgAo1wR+iXv2Pw8R3qenIkMKhChiN75oBv+QrgU/lRyivgaJxLMTjDc
b3HpKwSnN8Vb2JVXQrndANPAxI6Hn44+xSKxvoyS6yzJgz8CrS00H+1MWD8HhWnWmpvIfVitA97g
Zlt4zhOscvvzgGVOcThBUxWhlkhN9QMeBNpdumo8x02LFqGgPDKxs0dZzosv9ur6BKAZpASNwsQH
/1I0mRutQsVaPIKk8T3gFecreR4hlDkXra4CtmRPIQZ+P7T/owjNzkYqrB/57L/0INBGy7lv/4AS
oizkECxZPLlfv1D1C4B/qQlhFqDzLKQ7vJazIdSq/HujZGKhcpuTBjxVczw7g+X9A4Tq9l1UMw/X
HiivNCaaQmF5U5JDBE9yKH+Gjru9O66TnVkjySnngtnJoycG6wwlJL/f7to+uCCk+WmnmFUN1ocC
71LyGrtAVgTdPassi4T49aB6nStsdHUzLM9mN6fVkKlBbL8yTH8M6PWdGW/w0+OZqXQGOgfjWYxe
Z3ebZdos0n2wJ517mKiawYb9MD/IeI1wIG447SHyXPkar14S2sEvOpxGI7h73uFTZW2OU4qAe+Gf
cUCzEIDC3qrsq5geL5j2AulAOmhjVmQuTw25qMdjH1O6Prau9uTF8zlla0kUr79O5ccx5kDLwEUM
+Y8+OWleD4QHK1s3iV7GTxwV/8QNpWb2Pj11+CLzMmaIuVdDFvq+88ufsM6IudNL4ySJieFMavTN
6VPwbJJDpmM1xI089nQ/bmabOo9RaI48VKy1u+mI2Q+iDpoWoZPKssU1EHM32BuTMaO+u4OTv0HL
cwUHTR/ycJYHTf4v84kf5rk9oJJaNra6dZMV5MAlmvC5N6ir1sLaWz8B7FTSMeip5+CgXjQvqIAO
Dl8KTbSgsswz4fCUEfeu6uf+f6g6gUwH7phBfoCd1nAth3XpKMah7sNCk50ppbkzxWYejsg9384+
UdTRHur/d63OB/qXjkoOEM4en1Og26FrNNmtIrQe7Qka9b5xxupmzp2C+hAqnH4Xe3GIrZRQ2Pcl
slnBYw5U0cQIVPX7veHazKXiTj6bTkfDVk98EGt8/A1Uel7pV4UI8bE8XmEOfTV98a7xY+lxSUzY
sRCbAM9ymZs6rx00JuO4lynglv9J3G6HCeL/pNqvV8GH6c/2dIH6To4qyW0r861AEeFdLOtH0deL
FDYWd0+RvQj+TMeTLnKtPA0VAR8NeIyI2F61P//5RXtWDO+Xn5kOCpcVIqGQhpepuGMK+J+zYhN4
+JWCXp3MbfQuDMkT8M5HZWN3VFUoPrp0mtzXBuzJkUW3SIR5l5np0QTVPFYl1fFdr2WYi56T2+Zi
70kag/1VESw4PREQHBY8cOi8AwlYVe+j1yIg3Uh3srI5QnQsIzs9EPyRhV/x50+ugSuQmdIuvIov
x0Dfu9UGxN+njFYVZtZbBNy/SYTJeH0ncKN0gQLnm17GAGwUiHVEdX0/NOAjdfVb/AQTvrXKV5tX
SXePDA0kiUamjpADfwZ0kI9SCYnG5k+MYC7ohOGilkDLZj/HFCCX0AQr+Y9SPUskmXpWwvgJKfU9
iXzDf2nOQvWsjKjRVlnadsbxfUTxbs0MHMq5iifRayLAXfQeH/KBDFGDPDexF/Jm7uHaSUY6waPB
EGJGPteqzG1z3r43iTs+2pryRu/pz7z1LM9c8cg0rnmkIFB6L7MiAeqKL/oiwZJnoztOvDLD1+3g
UBKPJcaMjXeftq73LHjoNV+ZWk84/qaXkpBtiVickr3/AfR/yHhzfZUGidqmQJ+Q+7Yua6wENFEH
n3STnctxI7nk0yJQWHeNz+tV/CfBbaFwD5JsfB4T48vlmVGtn/6EX47Pe+HyTAtY1f0Y4mO1df8b
d7OZH36ZeEpdhwv4KOGr9jR35UN6YYz519OUnSBdAu8EHbDtDnMJrqSBF7sUZGlhoZ+dMEi7pc7w
mPCs3uhSwI7bBMrr8njR45rmEH7NkOzjc2Hi/9mtkXZRtm9Yn4zueDvFFaaaEf3etoJkm6G4P1K1
UAfTSO/O3WEV3bRjBDbIXMIgabi9OpKYcxuG8h8havb7I7/Lc3C2jTso0A1NH05aVpOUSZjYjaxt
etih/ced3GMYPyq2x1xpKVnb61PfFQbdYv3v7DUlixNatmCR2AkGVDj5klwAtPTtaf4OWY3ei7Y3
bgfKK7aaWKbWMbv0kpezra+9k2VD1UQ6PPV9VTS3dKdZIVFPrUpxscdFuy3bJ1frYNLYrC1ovTHW
diOVo2ppw11nK/xYo8mCLIfTb6wjC3QNFuuqLQO9Me0QBK2sCCJoIDnBrYjPchizPzPO3Md+nIVU
J3z7BGoqREuGj6zlC0gQhPLG0VFfmj57CRSU2Lv13c8t9j7Z7PRq2nzx+smQjGo14ExYq6tIjNHt
ro3fHZGrXnqLKJNI7lq3yIYL7nBWbZ7LrMXTxfsrgxpdrCFG4VTuNSZYMZi3+BGdpZF46YagKiXc
JY959lvTmfn0hZ8oCpfdWYy1tFaKitznJ8CNv6OM4CkAHffgkuOJ/dn1suajx6SCfJPR/j90+Mkl
yD1OuWtz6Kxmokhi+IHFWWDUBai92KAyxC4nllLWFGOzlKk7o0060DEnnw787p9HzIto6wWZrcAs
nn8ajkPifpH/SnaAvLEC7BJXuJnoHOliIpBsP6Esk1pLebMnORoxSNRmS9Yluluo84xILgAFG1Pu
kzotRcGyN17SETPNCadPBxfclWd3T3nt8tQBWP6/bpuLs5IoBflH40ZzuJfUhbIciCgCkAwOhekL
P2OZIrbvdXPwfo8J0pOCuOv+fzDK6z2lQdi0DzsZ0SqqWLH9tEKXuAJuuGv2fcFKghDhNNAjbwy6
EJzyHxNs9Pe10KzBDIYYsWftDqHd1p6WqaDA20Qc/i59mPQp0r5VPOh+19fkRSe4p9T3VBODXSxy
9wvIwAlU4Gdt102T4QGaTqsQ5PyC3HDidEgU1JffMW7FB7qNc+m6Fu29JLJsIpRJ4d5eMcz8AvcN
btXMhlDpqF/mzcxNUxSxN/+Wb5x66WmhqhI2TXIEj6Zx3sg2A6xm9Qg7Y4S+CwAuGFGfk7DjuCcq
UpNB8dZJ2AmD+eU8Po0s4du0p00qyzhu1U5oCi9ZLR0Cm5q5GpX9+aUjT2mZJnK0sBzHV/dfWFN2
UNu8QCBIVqk5mW3sPiNjEfpbFzsNkw3Y31m7fnUZYvxKiv3SNXCKl73dOoL/5SdcmHUFkbPcmdDg
0MYjZl8r1mcyPdA9bnpv9mUGBlLyi13tTUP/os8qB9MSnV0FptHGNMMY44lnviy5/V/JEDky1VD3
ie52rzBuz7KTMTwZ0efhWXjT3KEckb+Uv72I87bdSbKON+2BTj8Bkh5Dh7lYfCw1pyMZsv2q/TEy
4bYTr6hB0AdpBFHyeKLAuFng8Dfjj02BF5PKH+KF4afSnCbBTAfKVSafcr+Pee5JcUo1BkK/TqbV
M89sjRdRoKeYpSzG0qHrpQ+yTX9uKG7BB9NgxUoM+6t4DemnxxQkwKtykugidmf3Q6QvvQQFGJS6
Kb5AzVI/O/4UxUZjRSMwWWQqF/++do47ZN5mjsur2KSZXfn6XhLhjqF4OZynauuxWZOqdVpDHwN/
MPLE/R/n90YZ5fPmHBRp1K+AA+ypf69h75V6y589kcti4/eyFlAzspmHZgz0I0y8NMwl8X8woRF+
0q+ZQ+dY/4CHOQnnjdKC4wABDdWA1ikn8t3AI7qj9Jrg3+fJj/qJnW1eh+jXNEjB/P52B8BaLxnZ
FXG5suqlxYFofc0KCQptqsoEPOa+hZJT65y/Dj+kjUTnyPGcG0ZPRAPfyV4rW6yFWXYXj45q9uLb
MIvF8ZL8ZXn8/YkCVoOy60g45x1rnkKO/QgscQvCIjebnpwudabp+SZBrmwnbatY+fxSrWh/0LvC
uMmqbuDZyDjM6ajhDhSNrghVSokZfU+7LpLylRLZoGg/rCatmvdKC3n63G/gQrmehxMfUhSV9XU1
KynVsOx7BTM6CKem6XzpCG1dLpQDTIBMNh7S95KaNgDmKKLXvTpI85tBgRB6MoDfFq1pt7lTxXbh
HxCNEV6J0PknB1LnXLng6Q69pa5FRADy5N8tNT7f103wsmdFdk31DzAA0rvKyfrLh2N+yIb1so7q
3L9IN52yZ7NUKwbpWISe0rpDjYDuko1wVfVYEVyXYzsmoq9rBWgjwZu5sL0OuoQb15NeY218uX0x
smDu8WFHNf0oKCY8KyUCoxdr3+sSRnG5ocJxRf5WCihm9PkXUAaBAXeh4O1cgznv+HnDNYdh4naL
Mu2LuECEHACUAT+eNGuXcnAvn1bELcJSS92qhWYDRtZKflpL7O779vF6+GvaXXwftbZfmYoqH/pM
eiwJhtp1mEyQPqgkz4M5KRsqNJLwR8DyLPM6MZBypa1ox9mMRCb16xsyXQxoSJAd1pPYSLtzG3S5
BFyleyRLhhHN3ZondvRbV5Oq70zafy5m7F/8ec4o5GM6Hgh5js8qBImOcsOE5BbE+RWDtTT3RnOY
pivNQiDSKn4PalOYOJ4tqqJLKCd2caYyGU1ry1GzdK0tpVdJ1PZUOHRUVQbXzD55mReHaie9jPR4
WGH8JdtOYx3A4h7E+XkuwLpGowQQpxSDXoTE+Tca6FfQGBCkM4qEHPFXxfbbUvDI0qgAtTN6qIm8
oyv+2cchsRYwEC9bcgdYF6dXKcssJHcdQj6ci/jZmCuhFSHGoJ/Sc9qJElTi0xskq1AJLJdi9Dqe
oHktndBXeq/wFj3m7GJBojNH4g1l+M3OVSjvSy/ECP4Qjo2JpcuON5C/RcBlN/Vb9bgPw09H6TtZ
pEyil/9C5mkPAYBuulU7jsnWIi/iDEo7OJuptfXNsxp32LlNV3JIIaYCfYNW8wZsL1ZfSO7jsa7e
ru3afltam9nt26oeoEW0eUT1fgfMAlgrOZi0OzDGgq+3m0eu5WPN8IEJyt6QcNdUIi9prdNvek28
g26O0Zq9iXmIhqRNLfdBrnMuTrAfMH+HS+WkfTvLg9tl+jsNZE6PVI8ztNAgKvbsQ0MG0ICUP4NJ
sGzLqoSzrOD3VFUoP9ldTQK5Tz2bDIOjI+BpQHuO4X029tJn//+Nw8BffPUJriga9yNgm/peDD3I
HtBW1U1nEueDuiHK8lUcVVHdiuFGiCJ5m0Y5bGNVPWtvxC+2GkGGSsaU3Shv5Ah+AclZOACsBLKZ
vm/DGHPABDzhXt5oJ/wh1eQWsd7h2OvFXFs4a2sI8+XbolNlUFUI2399u2AB101sYZos2iV0YYm4
6ti1T+i4dJ6LnH0JhTywmzvlii0MD/V+zcrfPI8TF6TXNpULQSIeOauUafHuAbAi/km7sMdC74BQ
1F+x0fAzOrMSTuneOsw8/hUAo5J3WyOAcqrIBsSBAqcOz2X75fnv8h2v59FANWUVzNS7ktdZ+hBn
Z95awqSV+XZC0p60FNsoUJktKwkgcMNgnrfzhKXA8GfHLzKzbNyZbeAnWeGbhmP8UDYnMpoNSgTw
D2tdxC4qocS8uKGxyVs0tsk/hqqdcbTsoTVSET+MP/VOsTCmGx2Ib34vUwr2WFUJ9KvO1cWjpKAs
cXeSxdphdqX9xUiWabM8aYX5SC3+ChunNg+xD0IwVdp8wtwLpK/GWYvO4/18X0LyxiNW/e9zMRIV
dU2VnVxSfMhaYlP/k7U5ZquE8Y2zSz+Lj6UzvZI7BSMs0xVXLJS94qwaGvRFVeo5onH/MEMbqkpq
OcuVos9dCiJgsCkERuTkwOESXHUX0QPtlL1r2K5e8f/Vz0UZWHZqHFt3BocmOaeRw2LQSQ9KLJlB
qA6R7gpypb4XBuS8kczhnPMuwrB4bHK4c6KJyhhI9mILymOm2qaJR+g8uP7NI/7rHlKIbhdrr6iw
f/MGG1rFYg1NfdkylyCfe0muJJ7lfP7Ssi/2Jytnh4QL3hm9aM6LEOZFUbXHFwpVdrN+EOBH5SDm
pNPj2m4DM76jkYwc8tRtZ+TiE9kNoWAqMdxNzBCqRf76zt5fIqy7/PmDQjWOZqC9z9SH7hyX4/9n
0t0kox6oj9zerZuBaMhaFRc2YlrkCbv5lONAwhN897Kk/z/E2uaH0hIoPwh7vW83M2EEDtUe6dKy
w+hYU8gN8pTvZFho9InM3nh7xFr5HbAKSDP39mnWbBq3oYRJRYXMkQ0LUmBYW9Tg8yu2z4oMiOsl
mhuVjeyTrJkmwYIzSslUGskHKyAWwVOhAE1G3CuxVCt66T4/QtFSKlJI24mgVxq5LG50bpF4rYKw
mFof1se7PqGtWIUCVHa1E0++qfpm0waqIFeH34Q+XqPx68H0xz/O2LHXrv/zXuTRLB0n3LRhxcex
ua5Wirq7AtQoYJG4TPtBJEa2WVC7cxaeIKXb+T3jhAVoi2c8KY7QfUmzmXAwfnEDVRgsZziI+/3T
K7Wo2i6t3VKc60MJMQFa7L2/jTMcIiX08kCVJVd6W1P+bwg/5bvM3brpLhulVj3DsPhhu+K/tikJ
M6BDPWLiq/2P3svv+0MiFONHsTIDcupN6IasnFd+4Vamr806YzCdIXjK2flo2mx8MgvF10q8bhA4
CuggInjHQWsQzNlu5iRvEp0mNdkyZlAKRBOhX3/JaPKsacs9RRDALiCk6+Okw7P3LR0rywmheMcJ
kxxDn3LidW5GdfFUuQ2Ov/7MdPl83ApUTrvNUVR80ajMKlvJ18C0WhxKnokBX2ngr+yty6hw4pFJ
i/qf6C1Z9/GNCEm3TA0NuY5eCkkt0oujNxkSfUqZ3eYbC7OhQag8doTUodo6TTw7LsMyncC3jykk
R91kuZoSKM5ee/Z9mVw1d2yaYomEoaLPOWYJYLePFdQoQ2qmZ9NBVnTTVuJIWqHtacaQIG86+p2X
vJSU99BaxBdDIZa0Db3i5n24DktRiNY6avETNAXPyiUjdT9XK1Eei63quNOHnRT7Sil8DGZYOXvJ
9zVsi6EOKjA8889EtByTsTYGVplTMFBIE6xVHSmXi+GGkseWB3O/5E8JotVachVkQu+oqUHsJU3v
vB+wzM3dwfjoO8IovVZrn/Gf2urgddEVNthVg7p/XfQGj3b1Iw0owXCRrBlC2H6vO+5RWsESSJOb
gI9HiRokA4gQ2uDjEDwG6U40TjFH+aJuHiSFB3IzNmznprCRTl+prEEZiMiZZGAoi4IXPn9p1Ydc
cJD1FUjyjFSGgsW19kjRc/fnvIkweV5EijmtVzbmWIlmV/WZzqCv2N4GX0kXRB8okjpe+gGdieOW
91GmvUqo0FFYh8ilUypuRQTdWxoaU+429knTZ0jN/nBk6QC/IKQRBECi5on0RTX4HCD0OHg4B8Bf
OxrYlx9uxB8ne706onh9nxOprWMQw4QTwYah3fxN2bqe6xkH8mKSD97EuFtaDpoeYP8yMWwn6oL8
H6Whndz9/WtDjLv6IA01MYsfKepR+Z9h+cB9vE10bp0aPYhAJqMLOnS6TNHn3zye8NtJM/SD5dKx
bXYDhxo5K0txBqg22cml0dZPmZKq9lwr2secAT4vIil0rfu6N4W8ej51RvDlzy+ERL0y6UOBqN7A
y45CWN1EsPWRZ4+gGfmTLdR98DubIGlxRA9eDny5bfC5Z3xk2yqt3VDfJ6+gTgppG81iUHPyB+0/
TYUb3jcgLSwecDDL7tioAQlHbc+3W/hneU8cfQ+WbZN8tcfcKvZB6DuATg6OVyaqDYOJCscFZZ5Y
93EBLjP2gm5Vlhv6l9GFWX/IMQchiKzG+T/BhvBuAAQlIhKCTEF7re7es0vTf1Z2nm/aHbxiNDon
GJz8yrMuYXx+AB/+ua/JZlp91PLayWwVXTOGYyZ5+XdeO+otylI/NMJ7iu6nADpR3A6y4SN+r4SM
568ZcFMFH2cPVM0L4mEuUQZzsTergywPJA2jqlLu+4FS6Dwn3YPWCBNS1RYP05ZZ0NNhL85kAJMr
twGunkIA59CrGHvaEVOfaPVDkskIcikWbspBeKqqRyh/VV5Qd3RCecBnQwYVv0wmA7ig7QBUvnY3
RMBTNTmSxszkU+MxhtmadjCZ9yoq+HKtm2FceZFgpnSWbqRv/nw1lWoKlnL0fg5yzgntxxpdC3+z
VmN1WX7X95P1QvtQn00Z/v/LAyFu+puG5SNDQfhZY4Ef3fb5Qab44pIeex+Sb4kJwGSnF8Iktqot
zakGsPq4xSqk8psLLwVteLkNOprkFCF91NTneDN8hIOKx5fIAi+pwRZErEplvvwYX/70T+7MI9V/
O+caMBmnU4hFEL00lOY0pRNnRqz9w2eqC55WZ+YuhQsHFdL3YevJZglRn0R87rpsay3Rjh5Vx77s
yqBA5GAPK3wW8dOxg6ieh51oJ69AZNZmg+jDiU538PJEVUhZscpCQhHEZL8JDEnGkVMJdR01hWTl
1AYRqHVQJeUJ6SWRyBhAZzy+azshBux5vJ9tF6QdwMuBBrZkQwNt7daLGW1hT88QZPKKIdEBbcmZ
fXhG3QDUFoJHPis6zfHNtFMSl3x+lIsb4t+9lbAhMgE9nfd05XBYYsRnKqqL1BjEUJfMyAsqs5gD
tuXyR4MfvwyZ5ug6RRk+6PwL1vXBxAHat+ofEpsZK4sLNbpr9uHQQlFgR4heiz6fYNBMOhbFKVqv
cW9Jjgj5xTGQesOFQEA8EFxGUip/0MyVKILMIi2AFSpbJUqup+u7RE0GHBrI+qTMwUpbG/1brZpa
E+wqJKUnjS0yWVVVwvYXzJqOXgUsqU2weezZNUdl0hPHQ5qr+pAuSxEjA/piXMK/MdjlAFIR13Y2
+2TngmOyYGHk5+MMMYpg1xx5bcwnH13T3EbPBCyIjPuTfbWbFW3cxLH4xUIYuYKoRxB2PBbAUGBf
ydlpB2ZrXwNYf4ouTS+poCvj9o9xZ6ayUCvtHOsAknLs6qBv040jVOc+rnePDdkvsmASBXi1Y7wz
CbVGOMNyc8FFeJn8Z+LpXyWczvZx0opin0BRfv9TMbD6cTban6xA0ceDr9Ln9qeMr9NBGY6D1Hr1
U51zVvtrvbmhsM4J6TrE++NnpgQLhgfrUcaN5Hxi8kF9nwTISm1qPnkLr3MF+MqHwWruuIjQCm7u
OHTiav8noKR1rD/3ngv0zxy9XZwCXsjdUfWn62vbSKiCkFHojCWxh1ev1LuWfp14WAIfeaf34EHp
wynp14Cw4rHvWEwy4ne4FgDeulq5/sN2Moq+jcbz3y2ZA4ChUQzrweG0/N/AKPU/elmZcWA+TTfy
IE9SBAZtUoDYgZQw0ST+yTmxwauJkCh+X7fOFXIvEunbWTuEwfUd0KsFDA2rTJ6RmHU+6ujre01t
9Ylq2SbnP5xBRetWWPDTDr3fdkVNLre/zxPfVlEv+x1IAeAOvahd74nUTjBK5Mk6b/M7Bsz1VnFA
gKzBk5LgeZf+kdyeU9M13iaBcMS1to725ENxWEgSB4dNohZYwFAoPXsNHvPkHFZU8dUonBmqJlg+
+n+42iO1x1o9otRp/ewEdweIkwwC40q6a+kfD9uRXLlkklaI7OT3eaoOmgzk6MXQYLz03LKZ94JL
BHnJYnodgc1/o78ZdFjXQRl6bDg5TnfRigPURe1DKlKG9SKiVdSDA/E60NRyx7ozuO8YwKOmoIWC
xaBGY5FMO1oQombR3rQHksnFTDF6Hdvsw/i1A6adaITRj2tlkVzww8KYpN0Y4jmVsben9OPV2RlS
k9xTfQyddeq9IUBREzJoVggZqiLJgK4JQVoAwjLzZ0gQvbBEdUwP/FDIczQzuuuUZptBGD1SdcZ5
2STNT6eHZ6VS8i70p6tH94FGduaDAmVCOfcKmH49MfTvUY3X/sQgdEklDubJrHHZx9R9pyT60O1z
2xosR78qRGBpwlm3Tfu42hDdmUIymWI7vPPD8rca/bX/1dmnzI5oiCqfSFOcr3zolL74Ax7R5QLB
hNZX7rGHJ/WE5rzX78qA4S+IH9H/zZ9FVzNa7/aix1Z5i77XP/zbaP2BcLyQrHoHbjmpd99fBNuP
f4/K9vXjVoNSIZKUzJmUKmnAomcOZ8vCktZtfJLqZ2Hrbph+7L82tK7FDRm/V+30+2q//tvz+9tD
oSn6ZTaN7h5NryKSZHUSOK8o39c5VLUuRhHJ4MI3cqC144qlerHZZ/s5g7lc5EyvVDaSqKLcSy96
hgQ4tytqnnBOS0XzsPuNoS3SOV5FnAvYo5GESTA/GY43a0rn6MQaWh6ZdIJR1M+2fvHIlhF2v/+w
Sw3FQnAW8irG9j+w2sUALwxfFJF5e6+9Ey6iPeei0bhGWTBVOUpUqAi5TBx/zbochmLvi6ROXqGC
/TRkiKJQM0jqcMkiyFrjKp89Ys39zPZqH/x1DVXz4lBF/q+oyNYGvu8LF6fYBk9a0yyQko0Tx4nu
3F/sQqOVOcmM8jmIW9KejyPPZl+5V+ZrAmCGS+Th2kGA8/QkygI5vEnMQ1VfodF2JJUV3PBtNMLi
x/ELNHPyRkwlJ235+mswLgFQpXSVKXuyjHgqWTsU37blmlgMQFr7fcDoSzQWP8dfPh4qE6Nb20hE
OX6MVDq0DrFIepVFlBZjl3Wh3L2Hoad8XcLxKcPlzSD0t0L49EENpQRyFpYHDiMDXfe525qXYmaD
V5kuG4M9r/GxPKSimahaFE5EMEgoGQJpONYivB5n6GJyJ7b8Zq4G6Ze+PQLrUwXh8WSChjMMgFrj
XWih03GqVhaqr28KiMsd92ENBRvZKXxX1vbRD/C8n7y/MlFQJQGvY1gyiB9TgmqGBMowCEb/DEr5
QgJZo8z1I0E9zvTLA2RfUgaKYU/xsVOre4svRjqmGhF/J28e8uOep6gMifH2Vg/n1ILWRZfoZL+g
D3idHwm+P9kO0fYvxRQxWGgnXFi1e2epcuoYDwjHcU0lJiIBmVE7RSudYmqjjAvKgYSGNFkOOiXA
lRx9E40StwB/I8RZGojIcyoHNyZ2sLKraA4ym1E1KUxPqUI79dISGNokwwbyQYZ2HnDE/ma6d/7A
Mrh9RFeEPUnxjHhU8CFE/cUSQrmixDj7pXSB6GXd8FmbZo7cCGggrrSHrgSwqlSXPRPXg+utK26v
Am2AllkTIiVvOT+UTCj0OTRnKu7+Xf6W+rpNoh/kt/lH59EuoXsNl03Q+vpFo1Vr7RBpVo2ll92U
zeeBqijfNmjgvNtIFb8qDmxTQ8xnNd0iGr6oYwUdxPe6AUAeYdRmVPg5M8c4sPPw0/EzwM9YCtrT
B4M4MiAbNHct1cOWny7kQQFcgqSlh4YuQhVTLSdjMz1LX4mK06nn64vzKu7hiIalFvLvQOyjQ9TB
h1SUhl7TXYdFyaoEjoR4LGIKuojEqrFizMu7FtQYpTH541bNRCcLCm6R6IrK3lMGygcSKtdvBgYC
m+lil3fTQgmxbPNh1EKWSs+xUss16yv2vLLoQPOEkY2s808wyjo6LefBuvt5tHMDxM/kgwU+yM3+
Ce9/XUY5BMn7nXoXr/kO3+q8MrKn+xoZ289on4utYbhElrVJlGGWo7GQAHVHh9CYF476V1EOV93z
Wvhj4QSeDbBZ9TF+XyqKeQ6E6Cj2ZG1zh4Oe3brFIWBNNU3v1ihUMCn0sh/eJgzK1hj9qwfTMLgv
aSOSB/AGatU5q1PlsXMMLgn9KizfUQ5/ycyN6OR4UZ8PpegUAj0jZJuc5ONZQwQgtON8KqWh4vGY
aop8J6FJAGPjymVajFN8h8XBFRe5rKulLBXgGQHlPABRkU2lxpCoLgi7UB+zFjaYtY2Xt8y3YIr3
AjqJoYjWdqulPBIL7lPbGyH571Z1WmpmYKy2ToB3Zlt4aigi+FEyVO5IiQJudj99Kgy612ly5bCM
spX3TL1SKx6woU61GAZZLI0hTj7t+LlvTWI3N+/V1BMgwQQmjxFOGVpp9oq76lItoY5ts4C8PhtT
q/svTYbHJh1nrn87qCZgpkXLy93twrFaLizjn0AMv8+6AA2z/ceB8aI9N0sjHqntp4G+EFvx0OGv
ac89SavWKpsMg88S11yZFIFOgutbKimunOm6t8CGdpb1vFsILYiTHZDZ496U6xKJaZa12/zl91fQ
mzQV2tGDCcIxK0LE1r9or8lre2VXRHI4rBy4yhYoPei+NAn3XJKDVygvfwS0gk7TfEIXOpCMsOok
tAy8J0I2w9gV4l5d01ztdrE2FrF5lGXJBd35Ogq3ABP7zgJheSgyjjxgDe5G97l5SPv3t8TkLmC8
FGYy4SCbutjfDDvZuqEt1gaOIE4W4gWjaQl5E8omkFXkVGh1OCcPj+sFyzbrpdXATxbzgP/ZUYo2
ox7jdEzUPYJTLz0D5HSs2nvQnaECi3PjQzpStsA4HBjv2wr2jRxvIon4uvREa9PEknsxx/cFhrbg
lxkbgy+ldWdKN0kI132orastpaHmPthOnRRJLE/Lgklg47cY0so+O6KHuQnJ4aEuAbtBFQ8EI/Yu
R4PShlPFOtQ8smLDCFl17yYqwIIbjp0CYk97Ft36vMmPCHqHcZUSI05qyJStIqEWqXgiZ2Z8vFNI
UHRgjB3Xcpn9aAr25szqwndiQ9H1px7SBriWgzv1Y+Y5Q67iz6OeNf9xjN+Kxk+KBG0zy8IXVxdS
pMls2mVO9bvKbcgwLUBxgg78zHcmX2rOj8jIwoOtJPqnvZjECKUFT67zhIdtlVGJy086B8uH5Lag
z2AtXoxaRKZA35K7saYpFMxkef3tqzbTLBHnJsoSOXSXnlqVnP/HSPEDpshZSTSwwZQIINMFvyeF
WlA8KO8tyHxfPggFTaqfZFhi1TDR4myMYtk73jX9ggGdmxo7COBLayDCJc03mOC7Pz9YjrNWy47Q
RLQwKYPBcFuT7PLqOXtFe1o7ZSNOfVMn6J3erodTq99T0srZHZqUa3VWAh9lU4hL5aJT5uThRsHS
2KcxbvuKujryZsr1gNK2M1sgViTnhWyLVdyIgbwtvUBIrVhBTa8WdQ2wF/o7xXU9U8rY3on29WQt
AtixyHck3wH9IGjcMKC9utcVy1+hF/dDv1CUD8NBy+6/Dh/ZVwi6QuUFpl9cxmB/l3me1OJaLjr9
q39U1e3eaVosRQB5N32u6J7tB0n59WYTCilWemPRnIc8LzT7Lj6QDlYUyaMocgmSTyk8RKiCMm0o
6PYZx7COcf2jhJ5UI8X168oeoA7rn6Vqf1YNQy4YZSw9bGBYC/IJAHXr8KtbibqRVNKVIce6AUXk
zRDyFfHIgU18WozkeKH9yWXMA0Dl2rUksg3+VeNCJcLfat6BIgwTwaT1uvBfuKdZeUy7oNfJZPnB
YhtMBHx7rr9R7NxxgTJHhUPFwFpZIHy7Um/JxoVsq+qT4kiI/vdkAqTsMaN3iFKozmrha1eGkFCv
FveivXl26iiRZLWqiP+rMKBsQNzAvwx53swZIdZHy4QpzvCCVti0XJhtlo+3uf5kA1Kg6vAYrCFf
oBczEYa4CflKyRl+5MSjugft6CsKEzYqLesmS3v+LUua627oJ4nrNrqJB41NCe8Mvlh7dECof70H
klWWUC7rZrbZW8Wbljh90pjdgQyIbXrxMJzcOj2fZSv8JpLEhuqyxNVhxKyvteDgdrv0mC4eBs0o
QmY6UlqM0zWoWXg5eDDbjCAKC33q2LkwHjA4vIW6Zc7cA++tGErpjzn/6/e/ygCjnvCQMSKGdCA7
Oq9uRT4o876LCAtWGM3ro2am/k+q25UkCzY2BdPVwdHimFRwoVDhmJjyKkRYvNVV6FjXs9yhCuUe
BRNfpRglTohwkYxR9Qk83OkuXSkmlnlESR8k0OSjWEqDwtAQUVxrUCCE3XIyGofuZ912h+9wjhWt
hddzHuN0fSJbvoovmcpRWTo7h09MPoMIuQDx44y3++2e86eBBNCR8qdy26USwF00tqBiXLbn0WXi
6qOoxMo7ihDe/C3/ncYyxwOaLCIiw+criAxeBFGmFXLa4TAQG/inWGFJ9DP3azs7aVPPSX/sS6EQ
3u9/lPr4jUqts8UnM/hqu8mR6XsMAiE4iKlGRZrLxV7MfEQm4AWIYXXtkswM4AImyaHESQYoji9e
Pzm9mYQhPpO0dqkxcsB+/RuZCLG4FF/8/aTS5fL0sVw4PiEf+3k09Gt3IVjgbE1r7yKqQBkyEgsa
sDhLHYQ6L3wtwptji/z4PmUmPQ/sHiJacWuuGJZsNDXgkP5iLEs3q9QMbNhIQJvcKEbeQrnCqh+C
noB8R/oIxZpym1ygYSurjZGLlRZ6/HgQLfWgh3Sm1Xl96ObGJ3idndQYB9oppCxMe3olva0ei9tN
RUjl4AXydjelEH4xP8KZEG3I37Osgs1PBZssuykSZtk8iDZIwjCGoYwY7nKYMVSO+tbUnrK1om5g
KUOaxQiorZiQQ7u9BPB4TE3T4HrzDjfC76uiKmW+aMXU5APhhB07+j8V7mO0fNES+An71/Qpp/81
nT55Oi2SkG5byTf0YmWy8TbkWuZ+xuDfOm8RIBR5RImhs6OljQEhNb5RuxofeUYldmy2i0yhdvbV
NLgRCVJfOBtranOXSfrVgTsRNoKmYiE5EQUx/+LhtzQL48too705lQFWb9MoPZ3e3CXvKywq9Sut
q2izpQwhT+P4WGVldwAmku4VAhHp1sZZq+nygR/5j+IUmuykJQfvjangKkztOo56xZs5t2Brxlfi
1W2Tz0bKznxZJQvxD/TA7NlQAn5naM31sKXD1nayV04etyDGpsrGGg+s+8XaRbghL8Id2QbyPxHU
0RTkJ3T6myk2H+O3wZI0y8pGld+qtpt0dnW+7dZjZj9W8kvfQRjLObG93aKMefhyoj9TL3BluP3n
bw2YwWM5IvEC8MBGGlU0oXmcnSigpMi07S8kQbEI84ccrsYoGQ4KKV5RUpL1NHLBivERuYM1T2O9
UJeLo7jOHnapCihbuSgBhgMsKVOP0qwdaUo2z5oJldNxWstMbOBUXUu/1Hiv8Er/BG/4G5nYdVgN
SG5kwCMuO0BLcMbOPW4wt1w/irlVCrgUIrtkcPWtIg9XeNa6eZSGaFikeBXX4gliEMIUC6cXg1jG
6iZmIjaTJKR2BUVZCXvt6BFiCDD3UegnMFJYrmOx5ZI6+52EfFE+tppCzcGhXY/wZDbZf7ygIWAp
k89HaLBmxEIhcGRh2ODsKJyGcfGutmwMe3jtUjtbdOm+m/FO5TULC4qmKwu969GNHwECdu2j8smf
mvocJATMPMUPfgysMMA2az9BUiaJdGZV6alpxzzIvOpAdS4c6UqHjaNCtfpoedkGFJTm5DqcRD86
IW+pQqxmpTn810dTSY25nnVar0NHijo0NiCIc3KnGGJWOaRNspmGqS0nybBP42wESH2UDbFvC3D8
I3P+ui8DgoICPeZSCNh/uPOCuGPg6L/mrovcN6ncgbSoCWWXGj5g6aPmaOnipQeCauuY81ajoe79
7NCzjS8eQpV66Gaqi/Ur8aMSg3Y+64HW+g0BxIMZM3b7u4NzO5cPI/NMaE6OlGkcIgF6JYUyaOUp
jpR0fphKaEDmAkptTbfCAiZZ9KIHaNSujFnE0fFrjSHUWnRvRUFuRLQ3bcmuMLPWL+MF7XxTD7LH
86PWDe/tDW3GNE8hkPMo9l1ODSFcJfuV4f8hawaWgYNp2c7rVZTe8d7te31v0xM715pE9ESXN8Qi
JFcwO7GnUBXgm+e2XXHUqQTkz1tK2vdsh9i7mKV3hdtCiOTnvvvuVLghaE7+tYldMHeuruGHB+hB
Z0r7PKD5OmyoDOwOMo0718+r94w+lzK8RBzYgzKfAjRkzIDBWl2JsBuug2FWRGsoZtW95NF/j18l
8yNoYelerecxjwMs3RmIxxW4n6GJ2DVUeDDtmy6cOFPc99qwx+mllLU+r4iJ5qdzTiki+ANdcLad
DtzMKhX8QRnQPYDYFJgrIu1bXUjFv/JSKtv3MgbNILb7ScGLkZ/zlqpiSymTgm83NZb4nTD/0D0D
o1xsyV+IebHKjlWx50nRrMBG5TKK3UUTZTP8PYOKnmwTJS+4mqKyNEPBFy04FtHGvTULkx5b8w83
/2lmIbS6ybS5GizlcXbS+dX19TgBbClvWT7MjFMVXOT8dXakPa6Vghef9Q1qackHbs4vKAZuUTTc
karZ4AhQUaOg61hNO7Pj7VQAex9OQimFJynr6RQcSbriR7waGyb8+yNwohi/36Ptpandhhn3SZkX
ALt/EOAf+VnzAaV6vaoSGWtBVJF5IzJ7WPEQanucLoFl5n4o4EiWFxyqhnTlAllCykDjUj2RQU+Q
Uo1jRiM3J7i8ER2DP9/0mrVjY3oNp6Bk/Z8elQcZydz+Mea6/Y9Mi2mZTFT6iqfW6ofGNdPCYPGG
xexPUXvLVnKzC1hZoMMEI5KhcJ27mPPfa0lwo74vlTSWh9z1HYeuIn/f2VBuwkIinrao/m97WCgD
VJJKmFFjQosdG9Gg+umCsLAS8lZy1w3x6aypiJV6TZBmNeVJzNNZR3m3JQdHELFAQdl+aitSs0BK
A6AuhP04CbZtgI/ZPwfVg0+F8zeQY/mZ5JwwFxH6Mht3a1x6nuJ9TfkhHhd4yr0/aP8B9NJtYJS2
aUCk9C++PVm7h4v4ajQ6EzAZvCTprhktaowrpczSWn8F2YC5oPZkQQQU27QZwibKo76OM+SmdSuc
5dklup2DuEYDbFy1bjrFwJnP+d8YT5FMxcR1VjdWBIUJjQHUvjwfBpGICZuPHmkysvsoMGY/cYLy
ZDX3RmCPG3bPFPJpTbFmC0Jkihn6vao4brnvANpbYFOmJN9+bgog8T9ZjaKDVEik91IjI3hgWQ93
aUNrn9n/XWBhtNbJ26OrrR0UAsXvDvfuDMNvkxZcLUqoOWO4WQ/npvyXAObG9zfQPq4jbLW11mTX
x+tMCzGo7YwP46ZL7hJclrwMFt2YLuNbnC5Xo3LdapxcPonbGQXsKpMZz/qdYAUGNqdqDJ04JqNv
oD+VxY1aZwfvT9jxE3o2HDUWJ2wJY3+tEW/Jhe9HAWegpS834z5NpOcU35SG7qdqu2m72JVOX6WT
y2wU4Rf9VV2qQsaiWt98Ex3lBgS1HUe9uRo9g7oT5qQqPjG7R1uOn4JIQ8D+ig1vd6AEPA5ilLKA
iUwkiPht2drJQ1bUcMH4XcMP4DE/dfHdl8Y0YTyeXA4ixhsxP7e+UBaBvtjGpFbE11K0DdZ7x4Lc
23msJQlQ7Zs1FnoQO3LThsI78Lsa7P+1R8qT5eWDyxcYo6nWpcZ1kvAmHTN0kYUgflfHEeGwsT6m
EY7IyYKJhtiJD5lJwjiQ8uOmp/E+mwAzd9Eyw1rh2ozU5zRxBe0GecVJjBI6hA/21q3HYEC9sIX7
7JgNFCxVEskIdvznC7bneOqUW+akYvbQVD0/cmC07QZ2n9G2MUX0eIuln7HV/AO8DiEQZjhhGs2H
ex4IxPiSW8bLird+wiHetOY/DTKINKylP6jxT6SzgJVFd1TXlu8GHPgMuuLaXoUFvYrCl+foBf/M
yg51A8mhG+fOyzK5SIwcH0fYytkklU8kdpugrLXLtk/QrJ9x+pen71LGb/WI91KlCxx1ZD6fnKsL
FyYdOnZPua1oeBdBr+dhnqftY52NcuzQOsBy+2WdsaMNOkjJey5OSqTeHDH5ipGCs/g7MVfOAazU
KFXGjOca8RTYUuvneMRoqIMGGCKstFVdXwTxTrTGRKtUi0jWG3z3B104C5BmDwDPHVCY2frTmosP
/vhocu1OAwLFHgqp6sULZhroUB/STGpVvbDUOw9Y993K6LfrM1YixjUuVI/omxsLr+nlIimPufHy
3dZuPENyqUH3rxgT/j4uKUYH5Ege8CbEPZHpbJcdD9QiXrcwMPvSqwrcgVeIIskUjMYDWb29SZRt
oyEO2gKFrTqwomE/WurPRw0zTfEbpJYd78lsybhGcd8HzFCn3LLiAWq9HzVKq9GmXikyqA/g5PJ5
F8fBO0WI2Q8+iGxGNSgCd5eMkx2cFyOGqk/55Lrrtd80rJUO2GsTihEsqWslLFy6GgeSAV+M7Wsu
qp0F/W7NmjK7qXT3H+5Cj2LCzH4oqxbQRwgilFqfr86ovlsQS9IaUFUxlquS13dJhVMudaC6H9DI
NbUs8hVcQeAjEfz9ZOmstaaEPvvKnF2BCm0eJBBwP081JnYBC9e8TmDoHAyTtGtGWIS2PiouCwSk
Co7KZFbgRwqxYGq5EXlOjqxxkTD6egTLYgMr4w3Akg7ZJTjP13y7Ad/SPcRiz7g7fvRcXakGWoST
yVIUZm0a8LUcOUBjp/HdHTjFuQWBvu3HuIVNTGVYks9tqT4u+W0QW5XyRyK/kBEBxrVvMqgB5q9s
ToL1Yeo1GFvBdyUFDeZn296YW4kmEAnW2OlUG101TvM7iH427hPylC+wrvIOozC8QKgIeypae3Gy
EeF55zuXLawTARSUrjpidhGr2pDUQ/68msRJbYdNGKvCNTQ0yMILwK/YV8/hdHwajXzXKAOzaCb1
C2K47JulO0xCVtJg4VPbhhGB3682k8471mWTP4ySTg9BbihFgN9Op/vVcDp9vRCV4ZWOxjN9ZuoB
LMEvXt0/Ci/OxE1TsQipQ1021Vonl3TfUdqLdV4fjLasvmrF4/biiEfTzOxBvR/jdQJelT73HRPe
7puLkznnfDYR4vOfAOJcFwZ84cvflKMM7sAt8DgEQyIymREb6shxJRWkF58ADBNwHLKViCneI9+Y
KicdIBi8brc8En4a7X7kaNi3uUW6BYiMULh/A6OC9mC352RsVBBp0TGjKwLEtd3n641BI39I88/W
TfvE5pNBlNCe0DtHPK1xF0B10lEGFv2uSjwHWHGxkoeEXF4bjfhOhz9YOkXmM/EzV3h7+8J4/ksn
c7oma8VUeo4zQvWxhU6ie8+/tDJHEJM8adGqUwFPAiD16y3HFTBEIc2ZAbC3YmhUupYNpkH6B4XW
xV0kYPU737nbcsDUjAVaWXUQ41eESRdKC+VyYHS/VBD27AlpAc969neOUTkbg/T9d7Qus64IHLpf
hvpebzrsyYoiVH5nySBQgG8xAOnVcT4pChZLKtneSbmstnAOGkZ8yq14mUNJ6dVaQbN/2SM6FDDJ
P+BSKBhmqWfeiV4xhjyb+bW6VQGCSNHCB+xUE83Krlrjh+93kaRTrKmlKliewThr4UYB9xAWXgjC
0BdXyh+CABV8gWOzrZGDBtukqyWjHT8dFW+rlyxEBrvGhO5vPi9gleIYuox6wXZRGnX5bjK71hP2
lAUG+m5J805VdnO5d6WOYpxNv78SKLRmcDbLiNLT7lbRbFejm/h4zo9f+eGgaFF8zXbUCf8v2J4d
mkW0+293usHxfSX024G2+SxzPXOhYKw7MzpL8ogFC0NL8u0BRoklzL2yjEhHc407wo8tNIEhw8HZ
ErRvqLHsdauIx/cdcoCJor3p3uQWPvsoYBahsOQpjn4rEgnITImMg/pgQibaZwqUCEtCirQKIprH
lmJKBdICtyb6qp9mkDR0cVnLWRQkox9TGqegfteRjH+DxXLwJln9sgydHPisQ+0nx4K40zdNTCOq
Qhf6f84eO23jEyj5XMVkSAAYQz+eq8aQ6Sav9jKU5Pm6v8hqpjOCcxAwx1iZh5YppBy35ddO1mt6
dGCF+lqeXeIYz5qgZi7VL+ESVTkMa1lplTwVjp1SCsaVdHOqz09cR+vhEnJP7adHNIGO8+xdyEMz
IctwMoDGGhsDy6bg1UEtnpRYfXVzuG/YtnVHcR9f5NZ16vAlFYOmNCH8063YjSdd7el0OoeJGvPs
xfh8z04podxJ16/NxpCtaUGVI60980iX6QwJ6DwNsyQ6B2rjs3aQI1BlgVMXe5N6UK4Rpfc+PFXJ
g14WPzHJdnLpGFzcUa7rm8VcJJ6mP0upqkzFd6cPsSaCTTq2cG1BeoJ10tcpKEGPLJxYENY/wMPn
cu0DzaTC8olYSNeIGyMxT1MKwoUAbq4r25tS+AAEkMJlhmL97dyByQXx5J1ElNrCUEiPurwfIP7E
zpJ223mscUz2Wua1seuzBKO9pPpXFkM+jfsnckBGU3MRGhlLVHGSnzz+93bsVbZlKd3SiD6gU45y
qw3+HZbEf2gX9GhmaIwuZ6TzPUa2hfAw9p/vXb1IOTv8DUy6r6h1e9hBAZVXwWbEcEGvs9ojdPxw
NXFckNHD19WzQnd9qqXOg4/RPRxrxYE2sU2ZAqolu0eMQ+IiBm9jQ+QIMfwFPZmzU2+qrYB2EcCX
ODxY8tv3cSI9me5yrohx886IYKOlfg/BNRHcvO2IzxIytZbhjTG/3LjOk0FpGq4xA6cxHOltWUPB
mXY/OYNxqA6d4ALcA9WAml4QvtjXjnjqLav/G7J0rS7NQmLWUmSOUvDYfJESA79OSzyhkoecvGkO
ChvIU40LbwuOXKLT1KFTFb/3qLooocjteC0knPG9akMqdJ2iMb02gAQ/eXEttSAcWPsBSqZyidR7
aG3mm/TY8G1Pr7spHooMkTXKLmwN/ZeIuNcszV6G3eyUgonKGU7RUZ/JcDXS9fwU8t4dgQYU5R4O
KqvxFNPCndrbIsz0q3AMLJlXRHhpS7WE5dBRE4yqWUe6AxxEQvs5lrSpuUhBbK09djlo+VlA+wpJ
Ho1P61ysXF95XwgLNHeoDA6zgOHqQYiavjexWqBaxfQ2xMaiK4o7Lfci0FurbuRDXBBFSV1PtOHo
zEv95z8JwHakE1XkFycI0Rlq7VY6BfK8l3F430e/Z1L/LZoL/b9hQwqpgDP/eDvvUs6/fE9ALjuF
1pytTvphHrH6tFLNyqsOx+j9k6rTPMGADdIzVQoz8megUSvrPRbq1ZXfTbHOUbr1eseP8/O4GOEj
24218O8nKLURbwjDCsFErvftBhGuShJrzAB4J/QFLuqxiQKOj60JtsEHvIPyxkaTwJfr8YxIchXH
mEOoJzPkyL2RLBOwEysexmneegTi71uevrhPkb/+9SoCU6XS9aNgnKQjtqPMaw7XlZyAp1dbaDfK
/LRcFzEK5yFEE/xOB+bwzLxBZ+fgGEcV4HbPGbz5v9eVf9VhpW/lfuIh8dHaBpIVcYeEStHau8mY
DRe5Gu3wsnsXyFCga5Szdtx+sk2srCsXyuRS8aCjarQ15BIOcIm2Vda55fnOivHMpwvBUuwMX5CM
ZqD4tujJKBeoZuwYkr728kkMbzXdvVhS2lRrvW8W6FocvtDc7TAJfxvVLLI/kF2M9NvWyKZpIqWf
RwBP4FYiCzizv9/o+3x8uG0ySEcVkSmAHX10a0P5JP0FpjTSs0bgJGG3CbUCNkyMQxAZzj29IQ2l
JPzctWGsCiaS9HUi3+pGoLELBjk7xI0i+nmfISRDhGKp4scDrK0xTKCAZLPvMxsh9WLb6tn1GLIS
wSmqn65dGcaWzk2ePFt7Aagl/qL2J1ZoTcDJeCS43WXxLIHX4AFZc83DtAOx3m03yD1jlQcZx5lR
Skwn/DZyoNCJPfUdPwVkK/mD+Jrqp9qN95AaqAnna94jcf1GryUbKVWXmStZcG4ZbMJBLWHuNF3d
NWqoG4DxNuPMeox9FYvaGFBbfyaDG4Xh2nklqDezgyIX88ZyskGztxho62ZN6G6vuP+IZjJxraGI
iWNxh5p7vMpkE6e2TpAtvnaTtwIdO1k0yPj6lk10lbQZLzzCX3bdLgixOfA4LbpZvATjmcD7Swid
LoS1ZQ1SxSYg6uJaCZK1Obtmno+qx43Y55QSKc9tXX9Z7/h6IsUIE+p9cvOYdr+4fuixS94SR4PB
BpSykP80f5YvvzjIJj2chqVvejOuxuHu93bs/H2M+WZPImSkBYh7nJ2pbxCCO4rT00YIDmOVsa/X
uMnu+T5YJ4dRFjHFJpfEDruFbDugpMyioB6n+cU/rpVyFQwTaYqOIbKherezplXL/muSg470F54X
fdsngx3RWvQug4zjUqs1jeC5tWljr1nLVYhx9SdQ0Go5jNEDDaWq4yaXFCn+oMYiXQ+na6I63s2R
WUJggBVrclbVdSndmYY2DhgrDe37cAgvSo2sh4fRZIlRwXoUcARVB3iiwl+9vDfXxL6LaHIq16MH
aECR2ny08B7CN2BuXxFPJG6epQpMvMktNiCk1pUK+z5hLL6NAJe8D/wnEd7pMuv3ZWhhA+U/BY7i
pztFpv63O2X+wI+k0daBdc0z5pTkfON4edFvZUCv52zzejU5s0Px8CWsvgjPafM1vqSiqjBN1MBq
VUFxV43ehdN4BiLzZQ505n8ZwqjEM3DKYPIvKktlBTrOUuEj8nN60pqs2MTvOsBBh6TOFB2FpiUJ
Ir1F7swzw2zXf3FqInn3qAtSaUbNaD3P/qj6KM7TdtF0a1qI1pxESAjk/x01UBrVJUp+VkLU345C
M0N4S008XWQSSofnG1jHISTAWJamnFtO/FI2F4ewk1KNZBfDdf7ePjBPV8ODkfRmwexI/3dMqrhE
iRPf2PunnwKQhkGaDf+l6dvvcDFMQuDX1HdVtzrHZD2Si27UFD7tIfwJ+ZYAetrcY5KeAS027iZN
mMd695PfvrfKyBF5CyyZIthcS7v9S/8ZsEXPmfixkc+WmkG8A3QhrbRtLvxN57puAz8svKgrUbEq
l/84MC5bP07roDwwQmP47nQrXM/GYT5nz5yLnS9L2F/j7wM2NDkFHUhC1vsj2dsrU34YcUGYY4zP
LuRtOgMNY5XoFA3tIgHWIAXWrCbyMeN1XahiVwbgnCkHusef79oiIKI2rx3qLmIcY6RxvGmDSxAM
j+KkIT94xW+/vPa52YpP43SZdyZn8QCvm+rGP50a/fjOPLYAZCMhyCEeBXkY/kbVg/FMoSfHsADf
lVSJ/9IIctj/dowEXZX2zP9y1A9DSLIGHmuK3hw2r6mXDEddNXMToYBD2LQ27TTwFDFVNQRD5zmU
2uJHs6eO40to/i2P9Y3D/CR1dZjLPGFQZ0R/q/XClZyQ9rrYLpueg6603dj0qNG5ThqHq7JyGYuL
6njueyCJHM8RwZszjWp19hzK0cymJCTCl6jFfd4a2RajRZN5URZdDfJXWIQ3DcsBs+Fren8u9mcl
nXmPGFTcQTJMhPsNs1BeJlMUridW1XDekCoolmykcjOGaTVEjSoYLuIBeS+kYBzxTOTkMg6c9hgn
QKxJ1q5wd1Hg3kdp00x8FD9FVRun7hTUIPu3fhnrf4iApk/IO49NaRkFcOXoaLAIXY5OOVsrduTV
RMsSZwfofhOuPugyNUPCLY1vlXK1sb5lOyIC8RvXSBxvGW/G8zztX6zIHJzKqb/bX31Vv/jN73Pl
lhFxtz6QZ4xSDUhRGdT8vGDVES3tcQUXsuhFA4M7ocgQrcVmUcrsOQd9AL/Wjb1s2v1Qx/ri5orM
PIZTWuyFvDM8nZeDGQnMKpKjtTY6jJ3Ra69ui62X1ug1f0c/eFCVwazJlk2Etm9YZMlYvgmIiZHq
z4KCO9EJzU2kRR3ntlQKdwxJhSEH+nzjijSW0sGLw7UDIAyjkNBt99l1R1tLjnmDZAWoNEN3mM3L
2vOccniCkwUriGrc1nyyslH/HS41FaLfFP7OJzYLLvaT61h6iVLd9kRgVHCau2iRor0jK23stgAQ
I4KIC3b4a0MAsLTYOBE6emHJuANxoiAcD1GvJkNfppUFKHzh486J6LHU4EhVrx5oMyeCfmjGcaTk
5Y4cfYMLJwpxHiouC9lq5iZJcJAnbUmMcl4ofpu9PfRIXqyLsZ0P/rY86cf7NcujQHafVmJZ6Gsv
C9uahptW+ZZuwFQLfWH6yryPPTU8lk3NSHmsLn6nFIs3qVoxwBtFF3+F0jemfHwS3yZj25TMA1Ir
3L1SM5a+FYulSh+RGMy5bsXQQbfmaJotyCAa/52qFBafZGz0qteNIKmvndhfq2v4ZvAH/b3fp6Gy
hFH4nHz/ydnJe2+890S8XLMHmBWyml49ZtRP4Jvma7tr2trxW968nG4eBJrAMUC7hTHjleRj79y8
gTvjwHA72Y4SzwSi/oImusBvs8HiDtDGnQXexMukUn7/UYUPvi1W9qWaA/pBwkOgJ+vYRoIKM+y7
z6DqfyCm8wVBL7OVmJ1avD9MOdQ8QlsIF17OpgYMXZUXi9M2qmjy1UM+1L5kfVg7adPw2onGBya+
XEX/wDq1LIAlDat6vQ7U6Zja+1fVCTQxvpnRFJEkGOMSzPKJySgBRfkBY/gICNlxp3CvTOl3M4vR
gJrEnMY073VBY0lZ6o7zl7EGKDaH1PEjhO3uwMlOq5b/sJ+i+RYsjeqK7wwR2lcwh7SUq3mYbrQW
9yagCSfT/rYPRBhK2CfrGbpfj82OAjGsvufrZPBvzlwo65hLacgqrQ9RxiFgWSo7maU3bxWS5ka+
usTfD7+LggZSmwqRovSz2/7kchWFgqY5sHnSZhGS6ACz6C9wLmcdagYXp9pIKMDXMQPB7oNmj+RR
Em91fyBzkQ5jGIOepGlPpXBrsm8HSKVjGzKrXA9jFf68H8Nku4lPLmWUycn2rB58CLN7cEFc7HYy
b12cHnYA07tYa4KFWKEvQ+rpxq1v8qnAznV0SoWUlk8cXuJQDCQ+TJeRroXPJAPRvfisZwobeGxy
Cfyuz54R+ho5w+Bu1dF2CDMdo/QZojwr/BdUf9IupeV2+DuFDC3QSQwttLFwpy1JTbWv50d+T0nl
YnduGJ+AJ3QqgyShq4h4urSrHwCITFIZaWVjBcWl0HnygyHZ+oodoB2oMrAGdwNLwZvHd3XsBpzC
MXRkjs/S61aBR1xgg2ynCSK8zgHd4UMACH9Ae9JAvzwl8BEfj6TPvIYfrox7G6UjYRmiu90BMNp5
IOMwjlnIYNWoy6+sxFt7BQ/HkgLcE8AIDUAskKFXjDCyxsnQu2vz2jOfODI1q8uRlCBpE1obr4nj
aUSZhnCAy2nwGBn5dVTPODZ1aOKU7DUDoxUMw0PBWpzd2sGPrsrZpbjmMDrY19Mji/JiGUmkPV3d
o5MndNjRFE1flFr1xNUe7kqFQz/Z7TLIX3pNfsQKZvXVYckVB17mPDsrME4b+r4PYNMOOPg/aqce
yceOTSxume6+rqjAxy/gcEZ+l4n3wttMNRqQTWyiYDN2wZY5TEUxLBCEqofwUxw5jFZjt1zX1mG8
Z+Z56QT5PLwbieKKeqhL/i8xJQY9pAHovbHUxPGV1mGGycze4moOT8w00+1IVWCx647BbxkSz0ok
F81C7umqaz6n4aoZAxy/28mcjTh12cU4Xxd83e4Y3EoNiTrt+EVy0FmtYdHpEoFskdHBWxsGRDeN
2+u5CxFQGCVBldCsxIkZ28eFHRpob5dwmP/qvJX7+xJOnObvXMw7c3AfBMOR0QqIzfnG1AMXOVU9
YXLh/dHAbTsNVJ6eIqzZtI6pnPtguqSzgQw34aeA/K7HajkmkYKjUy1wbA8h9WlMU+QwTJGahckF
X278TYtKh9kM1rJRWDy8yQFzk0+L3AmUo2OjJOsVcxTDD3wHpkV4p2NBe1hqfqaBmYVyYV2sXaRT
mbqgRfHu6yhMnHqm4Med1uRTMtRE6ZN5uyXWh3Q6cHAlIOV9JWuuobGVOjVAX2pqo79wjkZalbD4
6LfHgeQf3Krq9Q1cLfhot9Au1/VlvBwpozHh4ExV68pHeXiwkgmlbvoxqzCTLm2oxQDqa8t48p0j
Qu130WUvBQcysRpDlnyPhHukzGAWl3Qqqs28kfxHZyi5rXQi59SYUWOu6M52VB0L20JSqD06aP8m
dDFNqvH5mm7g2Iy9bzHPJAb5WhHTuL1BnU21bZE+P2ewK9sQn2k+KWC1+yHHS9umH4U3I27uyQD5
XG5CNjNfqtr6C3/kgSojpsctk8V8SBWIUrCwNFuMnClQWhEV+x9RAOQVNq+IODA4t7ppWa/VbBrj
7D1gOrORHUZrLWpQjAxFbRPsS/H0MFS8B9Aplw+zK3EVt/AzJonOJllwGS7O29Rd61+EQdsHQCyg
h/B8kKKdvfJkULZZ4eLB7w2R/6qV3LtoHatLrUytDtp2cersMTGEq/ME4LiFgecbB1S/KF59Zg1S
XhXEjIs1em7jikIZQSeqww50rHw0+vTIU8fOwwEc5dzlQ1jP7giZ4I18+pcFjxaXlQNRVjiGXmIQ
llvY4l9YbGPHhPDnZ+iTpoEoeBzX3VDYT2GpMfNtblL5w5S3P2CGZV7P03HYKhrzCFY/4dMSlItM
h550sEypFYdVMoLQeD61J87j/HzW+HzDufbQjfvzk42SAKMTLb+loLTniMsk2B75EgJwU2KrLCLl
c/zMJTIwzwBoG/BkUb3pUYEmylypUehbUCInGZ1AeTo653a+bfB/f4l++wIVmcLJAKR+gu8yH55l
hnFNfjcJ2WyWCyNlq/7tCRnvDGkgqz2+NzrsP5GdxhWGdO5b/jMRq17q/QnR1NgklfuFt4uhXVSJ
4ihYkTSoFHyG9PosFLgy7iVhaKxwkiedkXgFnn8SPz4SDj/KlLjNc2tFuWWGYEHhVFF01J8lTd7u
jWeeQqv/HolhPiOFb9wKDJpQoX8INa35Lczb4JQqgr6Yio8cplOYs+efSZ/TSZZF1NTtBuYeP5+W
evhg2y0NlL34gn4Fc1r7I5dWuWNJ+N0o3V+VZVRQAG0aWs95DoU3RdOA4OaYNBA2fpnyrEKZt7Px
baOlKkXWAZQMeYxIX5pqAeNzr5iT+7Z/yJdZgHe3apM/Ni6jBww4yqaXkK6aadTRwJ4z0Rx/6TTU
ByxlHq+xQhBxFguZJU43cAgYhFCdJHaPbYkpzc1jkgH5AVkBeqiLntmhokDMWPTVCWJ5oWvLJyIz
sS4k5Sj7G85aywyfAhgBZG68G/n+bp3pLaHHfVba1rBKMU7bC842GCH4ANLcDrWgXpqzOLYfcn09
W47rWteF8c7mTXuB7DvD0PBAB34aHMMWGByfeFnuRRsZmwZPLBaL+09u9inf/o5Jst+ZVOPkW7WL
qHZNmGZxZibvRCbowwiKkaGEe5JIxHpZ5aTe6sRRUzjlISaWyAUp68VfWCAiksjNYfbIu3QmdS8S
uyTYkam9VOGlSaWK95Yu3t+CZw2S3QtOyMMNRNSnaSrnQTgN4DsemfO7+CPKoF/zOY4Tgq4Xnos/
A2FSJKXY4+RKC5XdjxSVNh1Qeq84IpQPEPPcLeJRnS3nGNyKbw587ieYVtz+lA7G+3+/g/Q8DEWI
P81SVjyUABdV7lbc2nouQEFsCbfsV8ZPRkI/UIvJYdno+MctV/d4VlnmNJ3xJw9JqGygXqvAEpmh
q4IpFz8fZ72+HKw+QmDbu/yr6Ka2xeSeUSeZzRdfxoiC1qfEU+zCx03UXaM6iH84yGl7fYB0totb
xqtGb+fcdFSbDP+jjrj7+NUqosmoVSSri/Yk5VECQivM9MxdBN9OuPlcbqoFxhs+qcSaqXgWknMy
NqUdoP8Eoigckqrw5FyCBbu5zgP6pU0FmHq3U49LrpNnN+rfLCt1Glg0uaNbA6NWZIYfK2kiMTs8
MJ3UWJteYRRlLwXj2DMDULuBbPs9bLJzcSt7aIPaANQ6YxGql0xEFNpL3Z5Iob/D1muto401j+/t
cJuKT3c8XVEEu//DSn9S6shy7bUJ95iNnBPEiWFpyglu/2/voZFOloUHCYZYBMpYF8dy5lehRFzN
d8K7mC3cbOAZbPHEBwh0fdBCuEBDpQqcKUwqwugyoz1G+19Oeoj1Hgb9iwjo43LAzKfTjgF1y2Yc
iQwO7D///2JSbShvCmdBAwJ/Mo5nHJuxL7+nzsL2rldZK5Qljf+d5Atni58A4UyAgrg2ZgSHvYDc
HaDjvgilrgb/HpQc3PYvBRDMnf4DxwbwaMpBg+3PaO2jUekTPTcukcvhIBY6clum4io8iNrV1kI3
5osDjm8aI40o122NlmDEfyQ0VN25X95EIFOJRSE0T2BUl+vOhz4zl0zzcjfrwGBnfCj2j8H49mi5
VRILxBkNH6erDgjPafi7ib6PnwYp4hbiTkT2BODjji9JCVzhRA3+LgysDHp4SnBvxokxDCuQGAS+
XFxv3mRF92n/Zg3h9eeNzE0oJu9U5dgkLEjuW9VmJKvE8KvJlALN2bEf0bQkwfWr2EwMuPGdQs2k
T7nkxixCXAV3IKRxC+4MkH/KfreqYsooM/TfiCSOxr3KKLjm0K/06WGa7r6x+h8fZoWP3AmwG3oT
UJnjStfe6OWDUw+WYt1U5+3TBdjnrH0kWi+qORliRe37gtGeUrKU6DEK2XvlU1VCyiSm0DIyZLyY
axuK/q69jCXyHiLY7FBfxI7ZM7AahiubXebRENMvp47Kdx9brtkjyzfj5WXmSqCkEDoHlXMsYG6G
6iwZQOM4tjVoAwGUBnn/hdvWSfeMXW9KL84vNYLujbvr8N6tUVw+ja+WvTT2mBbNBVS53MZ8/7/F
qX3XLNF75Az0W4pqsjvQCLCOWnJALItg8THMO38QMdQMRqUeczJgLVts0SWwkg6HtfQnQ8lq6YJn
MiA8YvGzI8m3JZaMRi0bL4q04sDB2W2Y55/nXnJ9Twf7WJ/1gpdDMkhIBXJZaKWLLN8U7wZ/aY+q
7xIepJNIzKO1Zn+W2KM8qpDGiYrZFfqGB+hztvOqRjxOrSqcV54bbxnMgNKlKXK7Qel9ZN0x4BAE
DD/5seCJ0joAge6zZchLRPfM42yIdINwzpf3GNP1/V4RfiOBYQqdQX7Hlo0FRVcTaLCpYKt3xew6
wjr+xZFUbsAehyjqOOws4nF8zyRNIa8Li+NwXm2ykds46lpl6LdBKlxxlFz5uYLgdYnhJgobEui9
r9gRuv/XlzG8firuIZ4xuWRdgljdFVf3y3J/u1ytQyTaptoHPdaAeqob6wCzicGKHwIHUiGk8SdH
JRtFfCwQU/Bbzrj1CHVrQ3ajxm2Gr1jxwgRqyqxdfx3elQj8K9vFFDHfEDQT7R79noHKfwhkxw7Y
onlB335Dm+EQO6akxrdAwMehH5C/69fBahBuyrUiKUxWavTx1Hk94RYjqKjIe9ERBhkk8YLeJAsP
QabgRxszBGj3mTOajZUmNdaBPiAa4Wzs45lHX1SkXbkezP2IwtU24VRp03EaOWnVyw9dWAlCoKQd
yldS62lk+nWsqBzWLzUNGQZ2WmKJ77Cc7O07tvlY4Up644c8NYoFQ8+kqKjgAipSrGJzntrwQOvy
OQNoi7qRJfP8Mo4adXpQjHCTe6JDrC7UzGUdMwNzGBppJ5Kizy5/ODzTuvUaKjNCvuG8lzc5of75
jmKnL67EB/JZwN/JN+VZQ11FN4UylCLl3tjvD3O5Om7Myef7iwE9OmqLy3bALqLt6mzFUkd3ZLYb
e7FMzZfVLMJ5uenGOtHYo7BgoqQ9r3NtvlQaTBJY/WJ1QW9LrxOriD3kphY4KRL8V4Y97XOph6xo
3Z58PAd03PUMattbDjDDuYnfDyzzy8zqkYuFJUaI1yC620CqJquM/ghXpcnKuYkzyFWSn6P2J/xG
LaNAvRWk4Un8QPYw8ojGOWNgyBihH3H4jHECsLZ6+9GBpZg0Th3+j/WgAnGGLZXrW2YlWcAckw+n
Xx58U6skCpl8xqDJnde27EUu9z8ySu3ixsfMQw/Ftc96QqfqddrekWCslxkuTdb/Vdj2+1yT/HE2
0FWdVy3/8oMV4vPtKsH7+h9BMFupVZLvCUo+2oEguXNrPeEepM8kaxNoSPwEs7Bd/UTP+g79AO15
D7jUaMdzGcllzHVS530vxzvMQVTafz3G2W1SQRzhQB3S9ynVRD253cxLG/mDI719C4h+ov4EyabE
9CWhPw7Xn+TbG7YzVpFRmLKMTXUGmwl9nGvaIWovZi9n8yMLBrYxmnIRDSS6AYJJGxVis0fJmYMq
Gqu4Fl88073jAOzLXKI88bR2OKCSsi1rt21L+ZHIg87bKiIS1qnaTZQBYcfYB5CmdbkBBWY/k7Wk
G/v+PBENhhjSxbFzKXKEH7U5WRQRhbRLCQYgiPeHawswwRZzvvmZ92jvWcPJwCJHI+GOv2podcsu
Hh4e4FjbdtIDSBSbYNmqRpG3mFi7eB0rUll8oXbIZvFMZnXXdEskGVni/3pOW9ijGE1r8H7EpaxL
G8eG8YwmPwl3yqdCTrVrJ4Kxe+D7amWQliCRiquGqu4B3JCUD0+/TJHdvd5L5tK0OiN3HKAC8cTk
uQVPEBxqc7+IRmG6w7wjjXYTxUqtiB8lq8PoWMguA4BYlLgL2o6Kw10s5Sibsq78Za2hg0vS6t9C
YaN2BRB7jeXxfYwZJZFPvVpm9r52VgLh9VWv0jq9yoiOVBqnGgOSda8pyOL/xa8o6NWhN8SLkflH
NFLokUHnSGqlov2asOrrXt7v/AmWMU6cKfXoWgUYkk1zdgP2c3DB6CfcfwsbDPEwkSK7Xdx50Xjy
swl3XvVzosB/25SUo7ztMxSoTYek7EZDOFSC9HalFR+zsR+6Ym2Mh4JbUdE5ZSUjaKxOXthvIt/K
3eh7px3Icn867I3keYeadKGARP77NiA84skrRFzKRb00wTRoZEnx3JIhwIYH39sn/8f8Um5fPKFt
vUgvgcySgbIicE3mpikcBIDcZXFQwZ8r8qQ+ZcCRNWYk5RdSKSznglZSaVTfC1GjGz5VHFsjm5gj
U9bsnBCqgS6F6XJijyJMUPlzkMlTn2HvFcz0MJUZiYMoLiH6/IBQcAeXxFpt+3bKPjOJ5xl0MmTg
Ur895JQcs8OSnup5w5LigpG1kYogyVE7ClbNLmH8aO+GL5Kx2cOIdTY8r3P6z/32T2SwX0J0xtkb
bxu/b2hW85eXMciNMrpLlhjCYl8U2FEENnIfzGp6WJE0zegpWfLTIHN98YYwmhPFyJN9CK4CfeTA
yMh/dulixP8vKN/V4SONuxmoZKe1Fe5ryri5oke/U3/4pBHTM0DBfphLrEdGceze6kHy9Gnhf1lg
ZXusoIKEb39pLkO+3Zz7LQiIZgxJ6wB/U2B/tKPbOoo7se2KNFIGUQZWldX1TFeQOAlx4kh+8eh9
/LZjSuNyE4h38M8YgUYf2tk/HwYKl/FYxEA7aNZjGhzDFNv768aPUBuGlwgm3fhr16Vyw1Y/Tyq3
xzffbI00VvWBV4ystGavP4NXvfwhRS6I90eIjBu207tJY/MWhjMwUAfxOC7VHlI2cIjiNjVYufxM
ZaID9zBy0kFYHSDheq6mBO66TfxmTU+by2gUjMEbnSraPbEMEoO03Iy0A1xO+oyzs12kWyU3wPjK
EYeIRoYxbrVTsdaEJZHOAB/J7fo2JmM9Brr5Djn7njOZNKN+3kj8JJERhehq7p/Wk/PAetV+wlo/
TT4wSeDTFpSdx+l6rYFkwYqdHk2HimMpxjVO/BWvi5mJxtqXCNH2wQhfQ0Q1y50PA3KQbg2d3SYu
SxLSqx41A+C3XpXBGt24UL7ZMrzF/8wk6sYVt6xaJtRu/iDmWoMllj/b2SpVR3Etr6wfPiIT5/v/
HBl6kOInofGDIpK0xCcnMftHeL4EJTwZQm3Kn/b9nO6kY7TR08hF8+4ikC60yYM3vvczA5iJ8xKK
0LkGgmkCXvcfKUunPqeMQNglT12PmOcyHe49s1Mq9uMIa30QH6Fmd20LYaWf4nkytNxNJhbUO18Q
zXQc+gmdP2to95v0Gzd+hf+3mgd15KDtmHA3TwGaSynxbF4DKhEXVYg/qs+6xEoqQazo9rBwvt/F
TA4JnUFlbDtK3xIfd5RGWNeoONKTcAOHCovbcT/9RHiIpvYzSFKDEWeSQoVhWVr0D3iyAQ3hpg3O
CC2xUBFaNOeM+Pw7Xqze7MS8xQxKCVnjzQ7l9VubUGqdtn/YKJ0zvZ701ujuKOdYf4kFykWFiWWI
LpOgEhUe1y06668IxzGlxn5Sr+HpkR+FkIukkSvBD75n8RBVSleIJkmd1gepR9nknVDj0Rc4eHr6
EY3ZVXXNujsPCUhdiQQf4OtoTVKqtP1mixjTedpSyr1ldsf1YRs72xMgsoOOwKScMOmLUeyJtqJu
JxSOI//MO+BzJC5jsP4KLfaOBwcuDMs1x2tzifzRbYV9nahOTNCt/MhGTJUPLhWKh5mExJ9o3xzk
awLZmweU6BfkeFV9emhmCulznsvTdlsBh5svClcF2q5vZV1RMMmBNdH4V/3Aj4+8jmrBK8BF+zpM
G720M4fQHNv0IUPEa3AJdRvP+6NDsVP2mtbjB8MRj3sBmG5i7tCCTwcv3NRiapViQgu3pVxw4zhy
dAPHVQ/SMKO/kzquG7iNug8lUIcq4CBA+6KuUjXNFqx3dEFf0Bup+PE6fdSZHQHgTDKQQ2bbBHPr
VeqrqwleJD4V6g3ewCrvWtwaip2ERNpr/XLEHAVDpvEdXvP+6po6boGdkJkbC0gcwJhmBmX2UrUw
3pOLMW1Yt3wSdttmCWYaCXAA6yZ5g4+q/SE+cs1JaxfbbbPOc3XEXBNXbf3wxZqOpq1X0mQwFMbN
iu+77SrbgUWXUnb9NPScHxVv8zWVUi2wfoIUmY2desqrju1LpKJoL+BUc375xfuaScH7Wic0IYhY
Zic1UXJofSJ7nLhE5B2MrWRPIXd3kOJaj6i+dr01SQzOo61/bzn9xjFy4YMMP/O9EfHcyBZRYX45
O6eFTZHo+CLruE2ciRqvatRNb1rV1e4L6OOt88mlxlJrJNxLTlNqKabfnorSSdeSvvhvT8UWHEnf
4CSJVChW1zYt6zbkzaz2kanCUAVymwJKbZF8XkffGLxHc1+VOKVceodjCCqpfjVBOYkxTLGEfDDo
8HoKHTeNfSKdUJbGAaA0rdkWTuPzOAiwXff/FM1vH723fyKIuMX/602iKDmD87VUlt6t6nJo5fWm
dz6W9BhqgbemKxkf0/msYFx5PHzBvorTmyxNoel802fPNdXaz7Pd6KtJhfIDAes+EpweEdXmYOBc
0YYU3KBn8VC2wli3yzzpic9t+9YlCOx/i1uA7rWyFwNY+GqaJTFeF53yng2nY88hGkDxXJvxJJoq
zCq0jDzpLmkngSMVpE1kk04NMCc3+I97P40s3qJg6J6CSu6PKW4Wqknn1ftIXXNTNV6rzWl/pZns
NkS3DNWY7urqp0WT3+02JN/FiSJYr9Wf4ULtxaPgf2W7NXoSIYYvXOy8w2dzo4VcWmNJPPdqA5dy
mxGVYgwjj5hhETRi4v3t2JCXbDLB0+Qk0rlHcQDFF3eYo8JC2ylvNAJcwQ8JLNWrvfFUkaZbxHTE
SCyytQoz8/kuL23uy+7x0uU4Vi9Y/Wns+54PDpxIVeZTN/t0cvOMxozho5p/MRsUWMC+kbSo+hcV
xUD2YcpWA/+ah6Wcyy4Kbr+ySrPgGK2ZVs30EXMvWTMo5o9d9VhSsQIaY9SqtgkxBl3PCrR71K+I
HjCfHzB2Awh3oi2CDbfdsivThaI8WucYBUdMMwUB8BfiSrg5fAGgNxJyG7h7VEh77JSyGb/qr9+J
lsmpJuxlBb3QVb1F5pYULbXSkIp1YUrcdw5e2Pru5n98LDVoy6z7vrShn/ih3mvixLwDuxMVQRH6
Gl1SoKJg2qVXZ6F+Bc/cFfqVvql1WVk57bckta2w9vAqZvFvnVfYzxwwoT9R3MlYXKJMFyRj7cWQ
Qd0jNczEWNK1tsiaF7XKJWRARcjYVJKRIUeCopJzWw6ofAHde+n/2q6/UHT9NlmAqE/+gPgupAKP
bZr/88+ULvSYGeDRVTmoiatXSxHB2+XRyyuokddewgU8fQ8e9gTt3aYVpA+UShDiSNbSm2IdfC4C
/rByiVJHi0bBV5mifeSba2jK3twl+3RDt/SKjK2jn2qKREuG8lpL4bp/2rbrcgGAfYuiGimOq34N
cAl9P2sNYYwH97luRzO9NX+9SkVBHKJmkx/0c7jfEdRrIslAD8XUy97jauK3KAlsXnlToZFAYqUM
wOSp+v4ZzXsBMipePYHMRS01Wng8oI2hLjl1nbNot1fkxrh7DMp9fraAeHKC1vOIvjuttmtiRHkd
qWxLXY51PR78Hp70O9gNJrzPAt465/M45crp7WeEtyS7VobTnRQKOfiZH30zDJ8sCG/jX6aYyspf
ltAODv/7IrNHzIOueEjpx97RrhH43lZe2jpGXWF1jRhrRgRnT1on4jhyOd4Z/wWtf7y5u5y4RWTa
RIToQ+UJ5afz22zID1jlbMQ7BXHZqj26j5nTYYsNgW3GDictS6JRh3TYVlZZ1siAkspMGeISn/Eh
BleuvD9f20nJTguAuhjw7rzEOrzQZhfzSsSpnqq8IfiaAlM9a855Yc7MgR6SzQyV/TnZtHcQJiP8
CGL2YQAzKOYOo80LYfSXH1ApTHwk6mRejnOJKCOwlYBVdh971OxYOMyFdCasYh9spF5EDWDSe2HN
NjLc9lYpuMPdMeLsh3J8wEKifsk7sDBjmOXQxIM85IWAEfEUBI2j5tQW3exPnAS6YCrf8n9ELKfY
i3ZYbjjyOuFREtr2z3UrHPaOIAI33AHy7ZFL0vM/4DDZmaMRqLKfaQP4I6Ol+qGo1qAfTVrwhw2w
1u/FzhtZgazEgbapszWt1E/U1HPR/LTHQiB8666jqYPc8r3i8Z8PqQ5xB07qLY3PD/b6UD1porup
IJhXAIJG5PL59jAyzb2v5Ikiwxdj0JsMqvx3GR6mxy7iKslUpyKXav08/Myi5AhAvMh0RvnVTMOV
uRkYX6PD2PMjpIqDbouTJm43OgSbxt0CsAPwy89wchUap65axBSlyzRKEe3wf4v+Q7utiAb/WTLB
wQ6ndc9M3AI68ElZawGuxxjnbAb/hNZWcEjqwB/aYAFWZKJ2Sex+GVI0iqzSGmM8qXJFpl3lz4ue
07WsueZXVTokM3uq3px92HFeIvvAZddxlAuyt0xpvn0z7xkHkuIWK/VwZBH9LNjzvj7xQQjXm3HL
/QQc6s4c5jxmD78dxN5II1Zl0yB05Wn1RuuVV7P8oGmyrSuOTBBAtjlS9qUtx78EdUNz+tjYXDNj
e+KqcVSQaGB8qzyVR7vxDW/QMc4g/lQ/4V8jglAGWW4WCN9PRvW4Kkqk4swFPRvVH83uoMGbLdk6
jUP07iAb+d8JyQ7mxWNECc0ZLTKKsoTp9cZ37eriZ6HbIGTOpQh3nS2y+uM4cHisClNzXP2D0BLz
KNNzqBBNKahRPVejccGAOlpq+pqq5pbUytby5U9OLYVhJy0nGEv+KYleR+PMOpofcVHu7zUYA8jv
9JtGJTA3/gMyUYbiNLTExRndziz6Sy4BnO+cSxbRJMhP/4MHDSKw+skFsaRuIIBlEyDHXGnA66X1
7uYFIJ1w7hkjfUN0j7fgZ7KUD3MIFPUO0lO8yJVQxk506ANy2elMEvMC7jPUH9FoO4shvTpoKLfH
j29unqvhf1rFOsJSutmeLjJv1eYvPIHzs7MB6d4thT3yoGrc2aYrvTe6RIIEHlmlKCr2rWiGt30+
UBbl67AqfK9ZFDVr+mvmjuxEw1gYo6jEe+GSkpefYUhPdvQHOzZmzdFXcwoZ4NRLyKEMA/E5M75n
88m530lMgEJO7c8XiS5yKDcU4bUzRqaZG3WVlaGAwg6hw31mHdltfDKQ26u+rfLZ71YlI7gAItqc
10pqFPapxV4kHqGjIBSD/i+4YUUha2hCu1MjvgCWJ8+Q7M9KpdENd9t1SjgE9ooh/xs6IkW7bl5l
1Zeb+NeN87YNXQ0CuBItVETDRf3FqvrZ1d+F3SyHTZxN9iDJIw3AEZehbACdbkc+sHD8JkRbvzgB
O6Cjofqpk1mHac1pAjRw5ClVlkwkdBAKubUIDO9b+Ic+GvBhjMYkDuGFsympptyA7hzY0IFcoh4t
1J99WWuNK5lev0OBuVaZEQKzQc3udePHYl8uaLPRplecF+QYy4y1UrR7vf3sCEivpvBxSXF97qxQ
9VT4kSLhMws86uwjjT0LM0RU2m6nK6Sm4zJi4EMVClSXGwqOREnFbi5fkeaJEY42cTP0E5kInTZ4
sjVpu6Tbzbr1wu8UNun3+PDFDr6XfkJ15BrU5P3qLYDnKftJ03XjHcm9gHN5oZ0Y29eTyHpCJSGe
lbd7edfkjUUWZxMcJpb8ooeF5PwUqQF62Br7IzW1Sy509BHqAnCBbBoH8DphzjZGkamy3EWv/L0n
t02jEDQb+RXx7qjTVEvnGIjmzAGa+ei9D0oR6WvvIlXa6B//M+ItDNkE95Fpr9LjPvB0sYEcudGW
C1CCyGr90Ln+4kxTqwBZoR/OrSZI0HpxAMZ2UUCd+WugbHugS4WKKexS+msXVavav5aNiyYRtIa5
1qo7o0XfI+GrX6UAD0crqAFuw1QDylEThmG6qhb9Oru8umTdEUstUt22sKM1zc8ecZvL6o0Z8h3o
ySgBkcvMDC21d8BZJvO23CFQm9QQR73kHfUkK9dKnTuGw7haT/JHGDoK9a9cqYkYcJd/y0vQTZ5e
4xQLWCcTgIWtPoTqSo7jgaDM/E8MxIL1nA046ElSBIxj0cQ0nkpJwJQDRhgVhhttBYG6ZRwb1D7/
+8bP89QtCtsjSbH94Ofz8B5hoqeDPdQggK3N7OqSzVG7Lu/YVhmWhn/0g9QUC5pg1vPBLcgD9jCd
GXLuKyjOwkKX6Bi2NNnKYtg09WBUckIgTMz2CAEdTqJ8gjNmZFs2Lq9P39EU0umXP2lWdPz4M9Tq
A/04Rg1RqpwscR9EUOUfUcolUnOfPeTdF8X8VUNprk/0O+jRJ9Ks9K1Agxtsffa5ZVsHvq2XSbKq
1SNYLgk9CFYBuu+or7e+83sHDAdwhu0gZpWRFTTnZqgHdrGV/36KKnyTaCmSimTKIDslK/yUt+40
T1rYcDM5GQq5t1hfuPZvVSz2yiMeLnQEyY/Nc5lU36hyH1obohvUcE4COagllu7OAU8e/iVOfXpG
HzezGBzPzQy3oQN6+8N4EyITt5skPMTeaHdoMkIW9T1hKFYZ0PIbFDHi64RNnclceS68pROzX4mq
QTfnU12eznuWjSZWtcCGsU1LNAVcwuapyOfdPtjLmhrsv1IfkHdJPFIedkjYQJQr055ndQ878aXe
1RNpKv46HmWCo2XkCp18n8FIU+hdNoSQ/I7i+Ro8aBRk8fI3J8++sv+JiIc+Q0Vn0KUYTr6GjS3r
HfnHUTfPDY+dkqjtT3a+IbXZSvOqBbnwBjlscCc14JAHWG/bFtg5pEOl09pasOMWGPoTNTscSJpU
P3ePjSZrL5Js4k0pEQwqT6uI/o4CypeXdJld3vjFA3QgoDdvHFx92LQZ5DaA1aEZvJvpwloo9vdo
6EJ32tYDE2Vbpj/TnFzNgDg9vU1/hnkB7jQOcBnWkVbgfyxoFdgOfwyE3ynJWuHRSwOhrWdu79jB
GUMPk25VGJvkKH+49ylyvLaegKU/829sPVqKA6R+uuLkEOMo2Dor6gEjtTTFSDCFhvFJK9lT/keP
Z8Cc+q4w8wcosNVHU2DpnENYaHaoNsMo4MLnzQ4824gSIWH4lI0Dk/GWoXKvPqv9jb+1ynMIFj/n
q2MGOTq/ORkX0zerFEhhqi9pOB26l6hEEpDWPJlMzIwOGId0wYMPaPOZ9mfPUGeuiltY3Fe95OKX
D5PrU5qLdu+84zNJiPrwQy/Ys4QSfJATZ+QDPwS8SX4dOJjJnWpOvpT88awlhuVNZp7SHjEO5siR
11BBV9xOAWIu8lF7185ofWjyQaErBQV+ls7qrXJNpewfMfgn7c/bXvMGmTfeH6EBea64ph9UAH+V
TZPqLf3GOFkfdLWgxSVLlvAvYjlSYvbBF8842qeVSMBhuR09OIiZsHGyp0e5SHTe8e0t2aCX2/Ct
xBGjw9u47MegYjBY5Uw87L00G7Gq3sHQTcXfwEDaNOBZ32AziIAkNgclYzXyUHXZCmLLQVbxmNd0
MyOUI4lvDW2e4tOOWebf00jUzzO0l3mR1wiCc/vjae1umUb1NJmifaoctNsIMdaLPT3WYMSABQZE
uOWmlpY7pts0ZrdV+EsfMf88CnwVvbzLwXK8Njj4Dzf2AsZF1sPyQHuzFUxheIfUqEvmwsz3WbaG
ZQMTxM9c0LhGwxt0noL1lmNjWZFS6hFQWk7KKVvJnIAW4AioZE5tcrXLU/q1wWgS2xZ/9fXsiniU
DY3jslaNL9nKzopM7mikUlyVS0FOqkV9IRVIOpe9+X3lhcB6kN4p9Xq9Fojth6OATfxx6rsFAONK
mcqvEKIocty9AZT44T3amiOAKjxp+3RRPSgfkGAD0vDWoKdfyQHMXslePCAAKAYSGYfem4JiRatG
zh5bivzsZFquMjeRM6RX8NGovarJWhehj+pwXfXLXbjEVBUPIIzjDXYKhWm/Q7ocgWXlxfqimvl5
Dp5im6Tux14+2HVTbJKOqFaL48ZVPdSFglhqotWvBadWzSK0cK89IsK7HF89tExB75daOiWR9uF/
KY0FyA6VfI7vhkrRy0zhhRDd/RZs0td1vk+3QYawmqEbibFqJ1mUwcboBAb6RNXKzYEZPTNUQoyU
VvxyyEUSj8QOktluESOibmu3uVxuqZpBKsj3vSkhEHUDchyKoQ7VZum36whK0OSxEMTUrFT/KZ9C
QNUC/gx5byvwA+l1mBibXKT2eTx5NPohn3+xkNVGszX4pgyGrw77JtG1HgM1RkY1LCS3oOWlIlMp
u/fGiF+BuHJYXqUf9SAlnIP6cTM/KKM8otzomdc0FnEmXKu+W/PO2rDt/7RsVfibqORN6T85lcDm
XAhDKKJgXeRSpUf8XluX0H0kOWQnTglP/2b7A0TfRug+7DwDI0ke821ZbZhADPreWy+T8unuZ8Le
Bv3oznx8ZMbNeaRGF6mShCLkNzbWlTt3p6CPW4O45eBUctGX9FheAeC5l81vcAVHcSaRie3tHi04
ljNFgv919aO16alhvRfJeDBe0PSyGYZw8Q5u5gfIPIUt/ahrTmckvWKHOC4aW2AeX+Zkz3VBriv4
8FO20SQFphY+TPQv9jdnr9xmwGbVRm1jFVkNKwd/tHO9n1IP1kcE60exsnuaAZBB2cUE4JNFdUhV
iWG8gLfRa/uATSrUI6/eXsw7/wfjEoGXUykMi5wK+Xy+x6VOPM/mHHE8fepCK4UuOilkkCqST3W1
PJUTl0+Z+mMOuV7d5lIqSgzdNMr/akwK3ZX9VrruNpRgZ+LtOSb9/47ZxQWMuWHGeYI+gRDfK/uB
/lI0FCPGDqAadKJ98jFqJ1mlaGCKG3P0eNJg16BCKsnJyo3ovT/f7lOZgL22goJncCtd7u9gOXvt
HlTtL/NUd9vS1jK5xXFMr/9hDrn/iv5Iph7Ru/yxnVGUoyAJ1rtfG2gm98emo0HnswZdfaMhIgl1
cwNdTgrQsTshJr6w0bA4SjhXN+usavlDKa+BNJVlll2QcHT71xR5PYHm2z7UDv3jE/3Bkfy6domN
15MY+LhhnzlcR+iolas7Y0nHEIjBW/GtzMOYGLRU19QowkDnbHED4TTtB0uhKm0qRhyPFtvBiBjX
dDJ/EoPd8LMiQpLSr3bx+wSQ7Ium8BH0HOBmh2SqD+U8ZLA2NyUa7BPqof8n7ozxXP01qYlhKQyk
6jQHJLO67reaRt33YbyyUE8OdmSwOHNWSxuEUnsGPFUfDt0QDlJvTQFQO0M4bvDyOw33XtbFs/ZS
YAqY3R7yRNp5/+Z5RDO4a3Xr5o90+lUO2l9oZCiA6lquRReozRCLwpb1YxRFPEGXiHNVv9nP0p2O
NEkul1UwDVotarq0+BCMxolabOAxY6NjcWgHQz8jkjkkyz1+S5XyOB+TuNUIlEAS/rX7UBBHlJre
ekvjW75eCIMUP5K4xJcETHtzMRqiykEeloEUplzjJuRfVLjVpciYNdRfskFW2+7DKjX6ANNAVzTz
XMhGDbSAxG8WgaG1A2xhbjro+utQzhe47G1EWA83PguWyZwOJmsV6yIXMOP6m1Q1O7wfgtgwofGF
EVSBhHgjjsj2lzyLPmmWLs1NbImn5yST7Kmq59FIxmBszqJpRjBKmEIBdnjk00IXnX7bUbtv90lM
zOVj13N97/QFMS09o/aYjRAetc119HGcL84UVwNMLCY+m2S33y5F2LdMVdn6OQke3mLPnA6apaoZ
neV//rzUxKDrGwV4uqJiuvSQmzTeyzTve4dKvWEILDyzDAK2BRI1uapKE6Dwij91LqYgv43Nh69h
z5uZb3ZzBasIbtRONxtNPkqcGWCidGlMK+YumTq1Nvpd53y8onyltPGsq6ch0ueHOWAWOpw0mSCA
dDjqoa74c4HaLJlHoibTWsdrNI9XAf61AWYT+kaCavPIA07YxOs1qETsrzeQxXubr8wvGV+E9BrK
QUyK+/iyFHkY/HMtPYk+87giLaMNyiOY+8TbNL8AJ0n76lL4nuz7AuOAG33iA+NxWeU5xfuunoIg
WKUDLd1GMxWVBOJCy39OpHY5TGVggxF1vqFnxCfSKRHTjIRBNxAh0NdwvbmTrt6I49Sh3Iismno8
QhgLCEW/INwFRo/HoieHqimTKeU1K72j0fTMFGo9qKol/5zWD5Jl2y3+EizsLvXxQX6oeo59PhRU
o+eIL0HPUNQ5Kqc5NJVXA45ShjBLaxB0KE92qbE1rqHVYi7ASN3bBc8lKcA9RC5znYh2VpUuasXL
WlKgMESVmZnt1cWe717nDC9QH7g71lI3ziKOLyuwG/Se0wm/lDpQwWxNEv0VGr1xgEOhMYiiu9K0
vPtn2Zamkbybjetp0TfS9h0FOavKwXjXkrQVM98E3ZVfxHfLhmxf1RMBfuObWTlEYIcZoTTH+s2K
rIVYxwxhA7nRdPQH3K7AqLV0r6ngV8iZhtdMZ5BsqRRq+27LGryZvx1pHvtQoMA6j+dEONTPXlyN
kacYQ7wSNBycyPsWFfPqsoUyfNePhUyDeNDC8fsmGT72zl1p/+rnnzMnNqcOMiXq1kqGscnoDxJ6
pj9XwPBi4liUT7lUc7qY2fM5A3Mq+88i8lAfenJFNmOFJ6VmM37TG4yZ2GryU5a36ykP1AgZ+Nnw
noJ6F6BugwbEscjri7FKEfkWfTmgkyiX6DtA9hhAk5PxkUaeBucfm9j1ff5SGWBP+5lEFjvxyI2I
vnWKOxSeyuplVYQ6pkCZlQK4MVqMOHoZCLTQM9XqcC3owg4uNE1TEFmKGyPD+QJXmEJTV/hU3BST
RPbWWJrYPNuI+HQs9/U/ks5seBDeVEJnzcpn1uaRPdLmGgWTIT6zZ4RVlCR4Rkr1q5LAa0zQX0SU
1jjaIcBVTWpitdIjK45odVrVA+9bLejOHbUsUIVLN0Mt1oILYQHjb3WAg47miFFLj4+d2f9sp4Vh
TdcvCuUg7AmF109rFDso9wrNpHl0xdWC7gtPwAslZLJqItQoGZHyYSAAVNk2g0C8THUqhlDSTYOm
5vHVm5tZBwdcSCLRIQsuy3riSXihwrESpMItpuqsxLm33yv/ro021DXUbr/phyrpQxmCfbg9TFws
tWiu33KnRTXvQBcq2safaUNKf41Qwka5Nj8MeISzu6N2Y21sdnfMPbPLy+t7H+TGZznTjrIxvWyl
gN/uGng/Xno0AcaN6Sgl1EToSJpyVZX7R2Yo8TdC48UD8SserekBV6HTCA9af4RyWjlHdgL5Bvds
oudDNivLhKrbmnhR9AKfN2P+qo8OCKUI9BLTJvEJ9I/xKnjbl0L3YQ3u/uz7SUMo/Q/IWSCQG8MC
Q8Rot3bO/KDSalNrg5Pgkah9ewNs0eIhuAyrayLSOQYnUS7RX4uYQY25KlcBTIRQ/m8YLZTM3L5m
t+1Zs+XbLrmPMsYHbhzkH1y80GWYAlVnnn+0RXtAbJmQPwk7wGAQkh61suXDkHnxdclm0fYpw0yk
h1lj8PbTLaQsTICnwzb4lhbLUjWpcLhKKeh3Kd+z7RyoQHeuwOlzRab9AgNq4GH6FMgAhfyb11Ft
6N8VYpWEXwXIr//L8XqR6PAhkISFGWw9ap1erxT72fMsK7y9/9Vdov8Vi49W4IdpCueMH0K5fdSA
xuQSjBGXQm/MSneWo1E0tNW2BP9y6wl1Y3XuNdT4PSx+/nCQfZX/MkB8Ygf5in/8sLbHrDi2zRMe
4MXlP2rS6f7r08RjBs8yD6yx1EZSu1j5h08mPNOWf6RI0Cvdx6Co8tlEhmNVW4cE06wG6sIArDZ+
+7YhWfIFfjQaH9oZqxqTpqPsbMbB6UFQqkGcu38p7HoPvvulq3+1ARLpUCWe8OZMq1S1ggCXt4qG
8IvvjsGakLvOzTuysHlL4r4NbEV+fvgF/vkw3Hvb3kj/CHxjsH/oHWhKUa+IZ9WYBgQQaOGU9Cbj
tuG8RYEppm4G2ykPZdCmhhRJRMtMggNSyyDXB2SXQjCXzPR9K41F8Gp+NxQpkN4nBrNM2+LYlANj
obuAt9jeTznYa4cUp8o0QT+tOIfPbEiMGwuJzbZxqhecnKPFF8qYujDlgjTncx2COltgePoPoOao
8nkowtFv8LljYXke1x8FBd+b5G7t3oHk6FjBA3Ql0BbZNVMEe6U75XLAW5LswsXik75lL5EOPjX6
w6MrnCC0nGUpGKzHqEUNztQzbTP/UwcHLCVgRykefHKO5D7OMHiJNB+c2V8A9gQcriqnuuzJJtrG
FrGAtE0RpBsMPz2vy8EyqPru1P5GQ99cLX25rY/Xiq7ijxzVxirMntujVGV+BT6hvZ4sJDn6wqkz
Ty4ZpCj27XPNif3BROZiGkmF60onNVVG/EXzrBuXH7JgMBSAWD39qBJJmPbtZeV4hbUySTgmkjNk
AQWENtQo8N5COuKWxI/Ks7tulAv6ZC4h2Um/fhLyXbqJkaKR+p/tafvvP/T+AFM5YoLeBAEDAZ6j
mHwzEjLJ/dYce7fIvezBf0u1ko/DDDzE+we149yUvO7fDXfyNOBoiLCdXPmj07gQViqFUnZ16+tJ
YZRfMWshVC5490cMAxfn17Xlsz4EhWKQZQ8dpjZjwH8xd9+qemkcshnlsfmsz3MiSFvLno5VtLP+
SQsS1O7kii/WJdeSrYkHxSl2yI5aiu5KNZwXpBfOgR/waoqekQ8qzARFN1nm9Q5TwRB3O77hVECO
7/DD2VzIX2bYwSoBIBV8mX4cHI5k4jwrE/UzbNPHeIIupp4iPuJDlkowjc5CU1vTK25i59LnNJ3n
GER1hLJf3klW7sBNZIhr9TiWznE78OwcmRvdBrsXpNTsMMrkz5HqbaW8oZNGVjVeITpVtLSc5K5k
lZSumhVy1fZdLQvNHsAxZGQPz3rk1bz0wZbyyK2KzZeb9zh67w8Hs+BrbTUy6yBDL34sPuUsfaIV
3fqdEscPWoFG14r/6STQNcTGPPOHnLup+AH6bhhsJ02lZ/D9uBSE3WkSvn3vHsaQzQ85Yh6SmvTf
wo1ZeIUUjH+4s4ZG3FZaIOS/tTrIPwe1NmM3+SgKl4c5xGKqUpXfvXRuXd7xr3LINV/d8lW607/h
V+Txub7veqfCApSMv4ZpH5olPJACHwRgWYW77wugcpVcB3dl4c6ldK9/k8xcet01G1mkv5opg3s5
VYYEYGrMfBMGD6hh3LprmJFfpSlBhd7QYBQiN6Yg0nrPdZWTzqkq6gBWb376koVCSJ0IunKcXCg8
Lv+6p8Yd+MIv0zXktMqarvt+vb0lpZ7hWDaPgTfIOc5v5eR2Ulz2sGIrRI0Fmes9ygvzITz4/4vy
NLpuoPOJdb9FKvZRfE/dnZCodkTOBSCQGGncxEoCJOsUu22pRq87t3bpLOZhBdZA50uK3u/F4ym1
wTbz2AqvzTf5VM8OUr80R81ydUX3f0DS2A8Yf1cQ7kjrKxB3W8OF3PONx2Vt32awAICRG8ZCZj0q
Bk5EqC4kCKkpPQTXjYhBsoZfDBgbuh+ytK2BFE4oWprF9qgKJxovH3RRkyPNALaFes+QodsTf85M
Kp+Pb/wR7jkSux5tQ0BTIWRuPI7kVJfM0iTer5QGuXgsBg6jTHtpAV3loAehyL3b+dx6uB9Bnu69
7ovgP3YhudsM51GVS6gOdWLyCZ/tlUi+fN0k8DIhZc2pC+zriiGTU+UcxF36cJT6cO3u7vF/3H4E
hydNwZ54fl3rBPwdpPfY/m0VvJzhRrpoLMmwyXvgyUE65UXF032dYy3FwT76anf5sh6WMP+wI5gf
2oUeDaNQIX8UHToKeo40gG+PwkthIomnODC/gxjpeAJfJGXdjyy6zcQX3OU5usHWFNOTpExXPtvK
Rsww24eDlXn5Bp7Jgs/hSf6ZliOoKxVMODLkG9GJc0MhfUu0bBx5mHqjpYL+XBSMUXYsZhHGgYGv
MD14ZpltkuYY+rvaIsqjexE5l1pXFGRm2kIXc81+Y2gm+6jJew2LHLXqgTkpe2zWAaI0s+WozPiC
8l53k2KDCweE4kEjRRq4bW7LF3hbuoA3JtcyGu1jv5awy0TYjst0DAasg5HvbLj0YtN32+et3VKj
B6PFwy3b9tNyoP0me0S3ICVCl99ZMq+UXyGcgPGVMxIEWalQVXR3coWWI/HVqTYthQvhX7FtdtBP
XayXYr+pHs0zvS4KrUcfwQeuJddCYfWMjI/a+IZfcpjsUvplxlsE7ousWQ3FrR7rm/PMBcL5EFsZ
5x7uO8psO6GZCBMBEtUMvfB7j4JchUCb9auTg0nn8p4atg61n4gXHpaYewmqf0SthG0jj1j2zJrj
ivk+ZOpq/PtavIO5P6tqYffHFJnuUblSkrHEj89hTrRncFnyFbS8FaELVnIsue6nx+eNWQRwmzB2
081VM8xJZCmpvVfyMO8TTKesdMRH2zG2ZqKnT3ucTognIe1wTNkfhSPMYUXNx2n0sNw26c43daIQ
Nzp6z5LkSMbQhYJnKAb6Icq63f22MvHaMgonVlHoXdKB/oi3awV+oH+UGtrp0Fx7lV6C352sAFxp
iN5XIsEyL8X9wSqr4bmCUQaRHNDUFZh1AfspUqKNtrpr8UbwTY3Qc9/R7fBdk7dOihgmSN5jG7qG
JdnKqrr0Amh4zClQuHJ3oItWnXqulrZcJJlTt3pxFugwdwPuiQMD5Dg6V00lM0fBanvNtD2IGuzv
T/S7kgXGGmyME4TIg0stqYalSi6nbX8hdCJdJBABJARnBIn9TWIcZlBRl3yKbbY6So//IusYvR8N
cFzXKuEai1aAvOxVVTple3mG+tDUzYTIhfQi1vm8mEucuwhJsRheFHkCHOlL7I3U8zqcg1E7mq3m
VnLUdvBPrAR41grbcVy8GmXnpItYZyg4ol+mKSZg4tOTX61Otqnq/Y8feayw4FitIc+Hx+/VMyaY
1kCJVITENgj+mt96DliQsLNlxVRDq6yapkVC07bcOCozuLwCI0CoWYOMvZKwBiXl2hpDzzrKV7mo
fcdn+lZG5HXAjm9/lCXFWhcJKoxW60Z+GTgR4r5vfrdn3cUYh87nduJGLbzMEv0OFJy2EVCU25Fc
MvVyPld8vZ/yt25PPyjKfj444IGEdNwYJ7cc/wxYN+cySoTwJZhoWdvtg5HDoOM6yvvvIBuR67w6
k+5HX076j9bWYO7Nssd4TJkEaw9+LdRnMoLMLyvAqZPg1MY1qMzdF+iMXJuHDwMGHHu+BwUBZxMG
bZ7AHp85rqVBJkQ21mgrlgJlbk8Z/mV70OBYLJg8xTL69/pLExYZNuPpKYDVge38RJP13XOXVWa9
dfIJrWUf+9CvbkjyXHsHsDvGiIZHbb6b73IvdVD6wn3EE5F0kRfmZye0KE4yx1DG45XqiRzFOZge
urO4sdQljgjyYhTePIdP1YlocMghta1EeAjq1Hsvmnp+RA8akgBshOWRoxK9URURs2dafSdY7A8k
bwK/WKOaU4JjGu7gZ12JtItsXafmsY2uJncQB6LqWRtLPLt511H3sBsqWz8PJtxKMCAwxx2HCK4b
t351jkmfPDGciG7D7IIKPYcR7g4yGFKpknRLElj8QqPnYksoK6fxrXHUgg822TJoKhmaibrUhX8f
dVLYkCC50n36oOEAqgY7Cw1/mubUyvhHPr2w0akRAiwspDM3TBqU5N4iJB3cIjbWuIV8J3CUTFg/
m0CbVr6yqNfcq3WlUdw2Y2rmE3S/wvMhW09S15OzC81+Yu++euYMqhZmp8GMyylWZ0TuVfI34AQJ
5MiLJXKhJbUb0ffX2LFgX+4kaPMcmszcAieKsB/s9vV/NKZni/ycwb7zaHvzFlwK7lLI8I39nEeS
KwrxlGU7SRsbtXohLWV/F6vx7K16/MlnRJ4yoUtuQHhCR0MVFibsyKiMnVf/PqVMTo3xxvE/kYFk
7Ke6gE5NPXBW6K4vFa/SQXwTugxqu4Tmp7MlGZLzw2zP6iOVNrWIJF8RM11JiTWEksn9Towh7uMJ
4cKmc4aoPQLt/KRT/PAeH8OW4G0Ee+2AKY6mw97HCDd7e0lGfz+NzVLUZuUcXg3XU6YtFlUARs8N
fOe2Fsy6vE7HWFXntdpVW4TAdvZM7Ocyx/PC4sV6YCzeJLPvdtl9fKM4AlggOhZEbaxzKUiiu7nt
dPp92aPPX8jk9gYKtFf6N4IFUDJNnp1uJUk7wXXsgt5IBnBbMeMUhLY34G2HqxqN9MgKsZSC1hRC
Dilz3JIY/hxld9ijVBuad84UN3UV40S0TyNqdm0R6l4PYvCRdG1uHBz2E+F+Z9xomKisDQDSg5Yc
MOvb0pIZwVUHUnjfv1khB9sQ6ZZxWXsHhFeI9KPZPP86bRis65NE0CLBGlw3Og53/8C1hhAWHtII
mAMcRmM9+164uwuXxb7sRiajZ1VLEMCqq8uNp8LE3v8Z7Po3ToRk5oP9jj5V/Nl1dSzdJGElJxGN
UBFI8sf+GFf0+SHYRisstRRe7p8FYQ75kxXSgvkYlHzaiJngr/D/nJfH0KV76cUEFCylHXLRegKJ
hn7Qt5NL5sWF+p35Rk7h/8wHMcu2OXV57h4tFffbTqZEIxlvVVny1UNrJRTUmyKST9WTZV4v0ECd
7uwzzRXxxB9y2JbnZf/KQOGMR0bD7CSxuIkCPJm8lIGircHfkyunDXqg9G9x7Etcevo4MmDXFyLg
403zlsaOqEzdKafF/WhIEUGOS5SubL61rgsTx13h3tApZX9XBkdfFCNwcuUtRq5z0u8Mv2MfGRS1
c9f/nrFAZDEBw0FivOjMJB30RAzKUyeEiVYet3v3FQYxuA9jMljMjo+U8FTD6H6DRjKLOHS40l6x
4rdqbaqzwyYg+nbjNP7Kt5VexpDrY5YA2L/rrIU3zu5xD2opBRgk3Cqf0F1SWJZ+JlCtHYNFu52S
1HoVmNVyR0qprlSNetbSlD+jIgFYQinBqGbM9aPTTz1ZPvodAl6KWtwnC0bGcYpHcR3qDLIrCAAM
GofuQpUWFGFqNbBybhNn6TeaAJmTNQqbxAJT97mkgP0ZxR3m2CcD7qRQnIpo2Bmx7bqKGh/IRnHm
tjsTN51PdLuoNxQ3T/7KRHw75B44ar7f8cVtP2tZsPJ+nXE+PwwAjYNN+GgwDYcuDsn+L7l5eHXk
GHSnvP3wheQDyQL8Srf8jNnAGqgRGB3BvSiovg+yO1Eq/MH6BORm+RS1Gx87i6PpskeDCEr+Ms+2
ah+gIWaEQzORvcy6Efag8/Jt5SniQu+uxJZw5PX6FmDrlQHsxYE96UkTfuyOmA38IXdyxx1crH0V
T152tf3gC+tAlvWOzOUpl3M/Nch9PAdGYaD7YvpsKPacC+SjndO65Q+TnOcZ2riIuf07JI2p7CH/
NnyvTR+AF6XK0SQTqK25P3RxOwjZFCqSXJuvcro6P00ktoNqy9T4rtuU1Zaa3XHwXmK2YGbLWlMb
xCN7XpguwzTNMgIHuN01D1iajJI2edjQRnBadLjY4W1V1SqKHsEgs6Jizy+h+GZYOUSBUPam0mxl
xZOngeHNEmb+ElHjrucZTTHsQqUut0XrgUVYUgjqTXs+GeIpSwh8C4G8RTgtEy6Kxk2UXV5/pcs1
bc/d3yi6DPQTdPiBFN8NZoO5SXqCJx0R7KMNpvPuVHL7tKzcblQfFKKonz7K7dIxOe45mXt0Xtrs
LAMI2Sg9Ig0oiOIc8iifMJRRn+ZhQqove5RKfCS7WdyQfM5mMripnOZy+GB0GeJRH7EzPmf9IUtC
a13J5hWDVuqOXu4rmqBp/fABxtb+dCEcQ+NAHwseidQamQ2uygSaV4f1mnYEu8g+FRZqN6QUP/r+
6Y4EbP3Bd3Hi2lbdek/Vhn0Dv07XE79mHjOE5r5m80pMEuS739aje9emCPwJuisliUkf/QEJDAcB
tPk4E6pHnebzbmUv/j369otnYp7bJqXDZkeCv+A4ch2S9jYrh/JCDmfb+eQ3hC0fWbQM84snB0IO
93jtf6eaaPgUd4Fo2sXUIZLTi8dVmITeHPUik0zheTqFIO9ka6AD0AKn2ojEiAIpXjvwYMOfpsCm
TO4o4KHxik1xece3xXAxEF3OhU+2rEvKaO0+S12nt05qg/KGYbeKhv9cDWGNMYkZUJzU0vxuXouM
IjVFhpgFA9teyyBl9Q3sVvfdhGmyqkxpKLuzLHMLGtZXomgeAOH0916PIK3sThEdydkanUkptQie
WNTERuNC4XM2ANgAfdlF7jWcnBMcpaavBhqWszzzPbX/Wp3rkxLRQkJWr7++TfBh0Na4tpQKV871
iIYsrQ9m6Bt7sI6QBGwySFa9f/e0UpriS3n9rcx5sx5gnDo+3cs40hi3ffQ5eFoTt2KRRDKyShqT
J/9krI5WC2Qs+1VhKoQhDqsuybXFsasgLq+sL891thmaR7DB6VxMxXPBP2/+mB5VyjJw2kKSM3Cl
fRuCx+UMugHu88fVz/cMux4IHCI4nPS9W9FjMQKPyUBjD7uxirNFiyGTWtxqL/EWbhs8rQpLZKqn
/+1q4cns4/w/qNJb0prPgMXPNmAu0oqDXQJw6A+XkBB3Q6U0+Rk+fFviynTeLE5igVuqrBFDTCZX
SJF1yFgnVBLZ1NK+yYA6TN4n6dWXjUoWsOL+h72KW7W3hvu6a6yxNNw8ldRRIFPEBXmfs4kVBiKO
VFIRobuVsw7lpxdF2E3npgvFCsgPIFcqowblJR6h/C9Omg9hCizcrQlxQsY+ze05ZqO+RgACF8yn
PGS78HTAbnIzljVY97uZsyMatI4j2u+wf4iMWJ8m8snYkY3VHNUttizn8F0e5PwW8bmcgd4uNoGA
1LM7Cca2sqDusxsp9YTjiSwvSH3ngcfUT+LZQ5pS+QYyTtn0XDh2iRv15YrLMVmVMfnJHo9vrtjf
695zqYgQEemjv7zt82H9mbq8QXXgKP5J1IDxTPc4P/ExZHMiA8DnF04vSa83k0oFXLR8Pz+RxZMS
l5TFU/mYItePsOKoITJlaXzXIOHVD+SWko5aQsTUR0YcQizCePBiylTb4ePH+PqtUHvpE9DvzKHB
C7LBG/4idyI5yUZbOUsDkB/E52kj085OBcte8tYnSaC7HVdmmcBqCLeeX6YeCIIMV9k1+2lTCzsT
JBch291h6823Ncr3XDtu4twr/zvjl1K6yZ4rSpAq+JY4tgFb1E7KoPtIr17RlTmRGqxEV6qjwFbR
KZiV5Gfj+StlYJOuYuky7o4qE1fzZf6wnY5i32gF16yNRsHpiHZrf6AbUrYFx+XjDCUA8RJqLTBG
37gXcXE8K24h5uQLnUEhfxKBMIiygqVz75TaKdfGjCT9z212BnNc5CTE7Y+conOC9SHs3V10wIDq
ljZm1P+wYtNI/EIQg+9YKvOsAhXyfAmTlFol0NydcNIfPu0HXbVY7kQ3DukpTjV/DCaMRC+8v5JR
jU44h7BiU2q0OuiIMsuABa2UiNeAe2eInRgY7t0Dxf9DM6JOTi5xiEc27rl6nkL9NKmP+usq69LQ
/ka5l72wuim2bOqZ8KtP93YIr+b0B3xW3kTfAgVpVb+e+ab8Vv+0idPcRx8VDJhxfN/uGS+HIwkI
7oqkf3osHG91WvpohNVe0OqQ2Xv2ASKGy/UeA6tT8vWjtl7rSJXaZPPy96FERvpJOclyrclQZeya
cM9qPd0/+Kj44nwamUXXq5nidXmFN19yW3yqmgUv2j3owtHw2bqigHRb87TL4ZunY98BRzLX8ti8
kfvTGTn8zUWnYwYikxa7C9DfccODWdrQBR2qGG7rCY5acAddfrgHlFI/VL7Sy63NFiFzUJ5ba3b1
61Xc6lbaXf9yH4tJkRmj89tKtDwzBTY+dKsz0BE4qPZ3gWTlIbXwGO7k/x8zXknprA1uhHiIFelA
mRwtL70UJ9KQrT43rlCfBIR278tdZqT6Rn1c8TWPZHKN/2CEMKiq8j6owxq6tXG1sNL2OJAH6d6B
Luu2S5eGzzr5mrE1iWk7RixzLMzxm2E4IDizrhNWVcWQwoZcvE4ChGXFxFj0q+vECPDBtaFMSZGr
L5DNDB8jyiKm7QSFh24cBUvI3ceYJCP0QnVOPfRAm3h/1KFhnVOuTYIGYU44X60xm4tCPaR3lOhW
I4uw2kANo/3VyFXU4Wt+Dzsbd+/ogQ3WMIviBKiWv6mJTUhuIrrhW5/nDr28UdRh+Vnd46bWSBiR
PEScEH1vlnCjGMPLtIavjkX/HJGtjYfJOPI2wqC8B9plQN6jUK8u0AAhaopFQO1qzUNSf5wwpOvT
GoHwCi5sSVjnAf7NUCV6YBh2B2/s7C0XyfU+Ww9nKR6uvBHpCETe8lVu9s8OpjS5mHS/kJdMJUFF
gp9+OfCGP8AVMWWhaOB6etQbfMgypaUr+vku/JtT8D9Uf+ddp6YVlqzA8qU1DeZ4CXkHXBE8bgrV
5XEPoQClhIUe7f+dtW6FWOrkSNR/n79VTUA77MPcKWO2TLSaD50Du7EPJR8vPaL/7aoLpah/H7RA
Ah9XTdXW4eS6/pmXWJZQp5m2Lwdkn74+04J+KEzTr04mDgkev4/dFt+SwdKMAMYZ+QiU21Y6jMCN
Mwc0EFpvvNGqnwRrTzda8l9oRXueRK5I4XYoUdxLwlQQw2xb2CVZQUalKL9ZDBvep+Yt3itdvjYw
fmXpyEmXuVJzUxGF0+KoIFJTW3pVALSQWYXHx3zSLcxe9WJL/mCrwM5+1ffTyhShHbvukXniTDGc
kziFnMXbleEs2lA/J/o6yIeHbNracOFikWY6wIWedtVwl4TgOq+61rmGm3jEhp1c/t/5O5wGsJtZ
ucyIpuK5B6hEgg3TwKRj6q2I/HPxODGah4220/la8j2C2PlZK2K0Fm2R62FaRHFgagv7we4KSTis
lpRepYmVttgJAvicmfTFyCTT1oF2w9gwXdAidbkVvB5t34b1cIPQZ8LFMYtdp3dqyppAZk1iNvdQ
a0kSYpiJFwq2WRuXoeV9rS8gIhqprBVIrhxJ61mot+12/QDJfw1WKFnIcTGhc8AuS1YdFz3iCTn0
JokX3FBTEIFoQDkOMYrFsg/Mh1w6kB/g5r377MzL608jH/OPF32M6L3zzSkCWzfmfy9vOJML7Hnn
PSKs84Y7HRmPAqzH8kmbnGHaDwFgCjWueGwAv30yTjVO7l2ay6VERZlpVt2YPXF4xFlOE4piAXj/
Noyjqjwf1lJRVgQ2M9/65RQ9572pgbXZs0Q0OITduq6JlB8ZGbT67fRmW+xifR7OHmrFV+W7tRoW
KcbdLerF2Ae0AsWolxC6rElMf5eYXm2CWJqeF9XVLJKP+4xJTD0pjfK9I12ekKCuZfFX+fkGy+wV
X9DV8rgxq4Ax1jYfwztR1xFS6YKIqvjEvOri3HdRgHv/UEZ5EhnMzLQnnvt3nUxwcRZdhlu9UpZg
sFUsk3kETkqouOSF3FCU7+5QzWNRweHXd722jqVR7svJWze2Cser7RYlmObNkkMhwMTB8V4pYYE5
u17xB+rCeXI8zm+uRQAffPgRL65mrkz03FjdokAXSczGEjwP79Xma7RLKhOKKZoX9p1sgbEkbdeg
hp0D/QyNYIL2XrgmTK4A4e13Cf2/pQ8tkIooeU4zatMs7JQxsRFqWuNuj2BOtOoHvAdF+ZU54vOE
8pmQ2xaCqBO/ASJUqf3qJPaW26ZA5+jWRRlN8b9Q55qnRGsKZg9uZN6vR/zELvaaVj/pTQZ1EuEP
nP1DZt009/cehQlfx9Aav3XAh1Oi9JQMcqwQv4Zzrlq0ntYKEjZx/Ga8OSCCeH+Mcf0FgaasfFd+
so+fgQr2JjD3LE5Ud8/gkTXFvUK2pPLKXQLxPfH4uH1eBXrsu7U4rjIAh+zGrJyPQljuf+3MlqMa
2Bb3GKSEgfi5fJa1Fnf4oCE2nMMhnOKFFlxFJtZdRUubUOBglH/fRauPeoW6Mn95K+GXgHuzJj90
ZnJpYMA8AYM6vnoTVd3WpY03kGN3IN82gXvRVjTRM4UH21Hz+jn5MLHzWuH9TKdVAj0f11OV62Oy
8TQAf7PiXoTCjIgtLQf8UiHZNo1tLosFQzRT7LJls4eyrHgrkQ4XEYOSAZEaS8iXuE1eVrblskdZ
fB806AEOtfwMu3GzujlraY4vfX5iuOXob6eAgdIZlt2bGaWiwb0mCclot1jh2t/dO+0MY6/+wPEY
6ppkjcuS8O92f1VDIINW+9jojOxmvlH8rQF2IEbOeuGRoD5pk1YHOc7uGCbZP6ZAhGBTTNKVelFR
Lxv+hdkFfgbqpL+r1RkZ07Jbn5D4avDDuO1LTvPO0I0k2Q3AEzr4sdmVzWTx6FBtDNYzuuPbzBzO
D0YcAWdtt1GcUCYV+bqIDm6RG/DzlIjX0bGAMcp3SvHV/g8k8XQZUj65Ip231S9MaXOz7Vx6d5ul
2NVgScSGdNBRB7RoyDzGG/KVTnvqR0Wnj803BGwNX3LYJrsl3tl/Vxh2v5WR9Y+J3SRgUkgjqbyf
qPYt9WIPg8IQQVJ+IvDqd0VqLSjiQTTXy7VtYuHLwSa0pNV7xCTfyDSujATRdIo3aeZFMVhYRtoV
/k8y1HpsMNtBBTGUkDiHHNUWvOG8CkkwJk3zKviDG090QW/zLk+nh3aOMDcoVv2nfM1PfE3TWaO/
O2v+Rbo/WvFLeN0u8e3JgX56JSYJlyv4UWLmTWgpz3OHkgcEYlHA4CrpxjsGt+PdBEW88YDlgWpd
1OkIJxwX2psamhMKx6GcyxCzL90KxegxiKKL4vbwulal0oXJKReMTeYLFb3eG37nXg+qU2WUFpzJ
c4wr1Z5r2CJs6423TBI1DKU1zxfPloVXIYUsoX1UlcLFixNyODrSFvrXpAfgATMzf10ZfXNRN21k
9JGuQVuZVprNoidbsx+6C6A/3UFgKCID7gtkA39L8f4U4paELPMiThO3dfDb52y8ks0uCUNo5PG2
otMQW1Fz0vOCNSIvFSBDpkgy5JDW+VQeZamzbBYpPj4phakvq00WTJnWns2rqIqJTXeydkbUOY+2
2kgaFv8Xe5+wihq8Pv8WQEUxgNs1ZgsfwZxTdkhAtKg03p+P6WqZ+yhj8vWphVcyZYKwWldS1/2g
mulFKtnhxS6RSSASiM1WbtCzhOfZ3+Y2H8IrMcnuECu1TaU8qlfmPec+TD5x3EgfZiIBTaKcyuhl
rv2a8YWtFuyrs3+ysPVetf1jOHIE02zzm2iC2brnjTPg8HIE379khtpjt4Iv0kaL6+ZV6jn0R1DS
DnAYNmTKqkgPLyYLF7Dy04kRwlKZCfZlVtEFXGlqdQLQG9S5zhPKoOsERUap4J2X9516JYi5oCeq
aL4EOy0m4BDIoE27ilWI6RN7bt8fSYyWa1EWksIjqpfxOxZQFaxnRlpzhOxB3hn99sXI6J5fZqpX
rYxyXtMmNLm0P9Ap1TXb7FRUufmh6kTGdM6hlEzlrkUBczi3uHwatp1ZIl6uC7/wTabTXdM+Maf8
wGy5gSsmnF3+cGKBEHZZIHQVcAMWecd48WOtPBp9UxjbZ/YgAQkfyVw5MXaVJD8I6TTlJeQgIX8n
/v5QcmcgqOckAR0KS8WR4GqxGmwX9c0HFKb8jNQQyo4RNgo0uV1DXoeDyITisvYz93tCw7B8Khre
k30eLPHFFHUkPz2Um5M36RDP6VHHhpnbc7s+5qz5WFby6ywvB0xbXKLURtPpam7PWP2tH8dRw4kt
VZrI1sS3QtPIclxP9DSnSufNWnou5gKQTprlw/hW6HF3fps/PK92vD2dbx76szDHQX0qH6RlZoZz
D3Kawq9yqzIBwhnaPX4Gwt6VFtbexy5UJgdxJTIy+OiSLdazPuc6LPswdmflQLdjchf9vOzr1lU8
vjvIUUvWMaiKywIld3JeD9PDl+NCpPG1Ac7No0yJs+48sn+1SBt5eGp43JBgmRCE2Akq7H03A9Uy
qvvv4JgPd9/kM6V1ljfnEZ6auF4hZLgc8qC4GnvVhYuEM1AlFgGvK3eiD+iZkY5nzL832ajOrChK
dMXg02/3zKvJXxnsUcSPp2L3Lxj4zTGrkSiavbyj9gWnIv7cT0mcBa/b/8nm2f57uZHh3gZU/zv1
/fD091gVGFuGN9QB+eDZTp6XFLqZ1Tn1m/KBBZ6VM6QtuKAlHwb/18JavkcsrDmDWhUg5nzP5t/e
pwt0FBfkF5LfyUwXfi9b3Ebqsfoeov8Yjkxq2zsInbtujiEjc61ukrFJr2auoY39emwKMXbPlCss
kVu9xuq+h05Eg45tO2wJWQ9/TBbGuRy2Xgk5x+oPFlF9mlC9JKBliao0mmNATEDMSLH9VXjNNJr0
jMJUjAI3sAsO5/AbidjiEeKLakaNPxjf82dVNtjD02CrXPRqenhJIPCAZlJYxtjIhojCxmheI+hb
wQeKHYOes/hTERf6eFQe2sT+UfTPYZiTmOWpu++DXmlxQ7S5e4cXFPRuXCW8nBFVeMtHP0EMbHga
2RQwpTXM2Fc+d6z2AkRHysIASWnZQsU3xOX7qF7DAgQfQHGX6htudGxT8Ocx9y+tluxdQKE6VqsA
uqTX+H/mMVXgNM9yVqyEEmUvBdztJfqWB+4uIcKzjSJ4vc0XfnrUxgaS8YBRlkucBUO6TB3pLAv4
OhKcr5p0lM/jUMEbeqojy171K1hBamED8c7ZCe366Qm1MZpR2Qk8Pl6vpLxwyARxOKH3+kRIaw2i
XZF3Uxs40QlFlz0BPYtPkqAvJS6DEvls5micjl4nSJ+btYpl7v3wlnhjjH6zFlJQ4kvPQAsuesmh
WUB0Jrd0MDBd3mzm4bmF7PqP+LR38M4eVjryjE/rG84pmq7QX5/5rk6258FYIqS08vqM4f9U/2s/
O4K+eklDKq9WyWmuseHdtNwkgCnXLvSsawLeorp0QuIsRrl8IMsTRZVxnmhyWo11Ubjpc0TDLtwE
9KS5HhC+BNZ/gPnyXhgHrXDpxYKsygRXi2ya7OrzMUfdPgcu7ntdOwXDAOIHn0mvDCxpAAnonJiR
LknIXmwzwkSEkLR1BdvSvXOz2nHQnQKHLKZLg97CMihbbn4du6RhjgaKoVrYixL0K3bBcpQz4veG
zDcdWUj2S8P65ds0G7HcCS5ewEVZOxVMsaM3t8hS2oRHe6d6BbxVhxA5YivIVv/YKHyEKpVFIiQv
ejhN56vHa3Aux3Zzi8yFm9EH5hyb5WYmMXQhQlrE0c7dJuSL6HCrl7aYMrWQ90dGuVTZ882CejiH
MSrSS2prx8+Deg67kFlvgp61Yrp2JVaYZtXSUj6Uj5cuyiouv1NWUhECo9AOMTU35MqnhG6z99vL
gG8Uh2g7mAyFeLUJdH1vk4k7W+a3t6SuTNSbl+02Cx1h/mSZGwSp5vOGzx+cJ+yCbWwRm8L66qSy
aJ//E5KK/8UypIUFw+qMoiI9QMMGtndsSj4KnpZT7rpGDEwzI54sAYwYKLGgEfil/g3Zoi/xXOBB
lpwYVzblNTnwn4msQvunU8ZPsA9ft8Ttp/c3DXSUevxuNhi15VmvnL1gJcakAtDRoceFcso1ldd0
1QDSN85RV4W4Ghe/StsWwah5wWfdIDa1+IOWK98oRX+dtan6cpkBNdcclfraH8/0yO+rxsq3Nvh2
7ti5VbM9ExIJUZeCgyL5mYy+KwEea7pQ8O14l+sAoi+njQsMJYm2E+1svlElldlsm4kbydz+5UY3
QjoHD9Z3wdYAVC+4uqP8hUUAj19bV0g8tAjkvdlvQVbVKD0WU1AWnBff9ZZKBnGLEZUcWG4Uc++s
8ogbmOHh06Q7dZaFdJN+gS1wGKHL01RzalhLfn5kr3Cky/Vbv8JtdmdtiiXys61oNzYv2uQyDElh
hWnpWPmmQiTUxL79ZfVXB2QiquQZEMvpXNDDQ+F82x36CLvumn+auV9xn8ZaRZJnDoWB80I5zq+L
hfSpMHsxVTcPTBbvIOFNKuwN5++8nWb1IISXyHNPTFZxTdEoMUXXv4jR0UuWj8bULI291dWVZ7tf
SlUclMxpcw1Lf/7wE+QAUKNSVuzMZ90cwnUi6WaUrSTFPf3LK05sIJflrQhV6rVB50OJcBhQdpxf
tZUgNaGow0aLsqf3NF1o/h6o+CCbuWbMIS/Rm1ACPcgfEfke8ZLK8wPnf/47718hEpOCj6VZfQBj
PMEecCVBWyRkWnvDmAHPK6unuQ72dzV6/k3rK+2QglbiL4d1jCbvYWheuOzfDwZMNA2TuEwI3DB8
FAzIIce/ctZDc1kHZ0HeXhAumqVRV59K47p1IOT71SVWFLEB4aLWMnW0uTr+pbC5qXQ6SIn/091U
GbRpo+Bjoo2PrQKwVcspKBAMpn479bXR+mWGEG/wmJELiIZ5CwNHL93zEe/cadHHjTx2VYTCUV1k
vKKRSXyO5YOvKUiBwhFw99A0SWtl0ndnE33YtSkkXfeM+cIU66b8fNB59DJ9q0ZzpY/8Xfr8wBbg
z92AFfdsLNZSHMu8PtAamyWaU+bzP26sxlugaQxNgIkz2JY0NqGHdcqjOQivZ0jULUo9ibLev4rD
E+EPTRVDovgqCSACXZCWsVy6WPXXAsexo5rJkCK/MDIRtfG1rO5G0P6CfeortNtYjuNOzC0v3UFz
KtxfwMgEn11qBb72UHVaJ0mGSbIG4B1wDBkjCECa0f3+GirJV3q5diT41Z9r5Wxw02MbglDKo4Rf
Gn85ZgPOT/gKHZcEHIpCUrJeGD7DTFNM/OMqBkLJGzlp5c4CkD09/A9D0JNU5orrH5NIJBup20WH
UQk/IgAwmV95ye8Qmpa8m4Pj8ZXp0yMMH6jC/foJaBA1zr0/SLbSsnLdPO4RNccpmDAg7uLde/9r
onbBAmGOSuU8ThzkQURoJWPPzhK24DolGUB7de45KD/7iMJF3xDA+dU4zN/sz7ssULqWHrgdSf09
5Odkjrjaz5loTZ+4h1yEPKaXmUA9dXW3LYAGkBceCE/wQwSZZfKbA6DS9Sp6uHAgd5xfCg4catOq
jf+tLYWo1WdRPRMtshiVPoir4z+/nHQy6oPbYgXct5cxw2tCU5SvQRFJL4b1NA3sV4Bj31cHdwO9
L/9W1wTOE6oUDvbLR4pmFzNiTTcBFso4njMh3B6qXdg3zk9DiBTOBnn7sNnsqMLmvEW4y7vaV8ZZ
ASlkuFfRlwgioY/lbgy49Tc2VF3OJz7bBVFHGdgnf0qy80Fx1Caid3froREraEZj45OgeEEU6XET
i1Xv0yHk6mK1NLd1Xa68MNwnrdrZ3O9MVElfblb92TLY1X/8t2w5sxpjytI2BhBbvqu+sftokz2r
/HDw2Pxx0yw48QOzk6ZjNrUUa0vCFdfdE4hc7d75CD7hTQtN3YR/PUaRfGuXfp7ZtkGXzxBwgN8r
SSVPQLIk7vaahnBWbpAHMgfBVPjZAzvqswFdLbNcVwgqFkUAGORq+nIIq7HlHrgK9VEJjok7+vCT
7dBeywJhPAPeYZI4+Ct1I6+IPE2YnbcfsJZ7Qr7/w2ZTrCHmpLjC10NDqNiOSU+RXR/h46fL8W83
E9s9NYrtgDkBxYM1cHYwhZifLAa1/+r0Os//Matw4qsEnhRh74CuBJQgx+tY9brKpFKi8nkSttJ9
w/3ldKKf3meeipKe9qUFBmcjpXsjWEu64pRvs/lsBCNNrucJjIv9pbXIBHzjnubibYGFhnL4dZ+w
MmT/lEZc9IJUZ+oKn1SAEb22otKVS2jupprLNt8Hac7eB+SaBl8Sz6OfT8ht3+wKLAYw3ux7ajhU
+Ls1K+Ly5D+3y4uhoftSMFBuncjzU5s0/Gs5o1BD7sMhP4gMKGJie4+SXuve71YChFoi7l4xmzBx
T0sIO/4MHB+8crTVD3JjLsZksYsf4jOZDxLUpAUC/iasEUzb6ktp5HgDeVx4JckVlRAoGMu+UvGq
7rTvp2cxLNnrJWl7jbZ1EwqIxpAtUJAGqWNzIo08cvtaL6Qv4Qoe5ejEU/xBK6NLEjw3L0fFwRMz
AWXh5M95oGse8/GN0vBw2NV9E+QhLnyyTDGwU53s3NKwPOTTJXToFOcTpYfGgF2YL0vW19ZKKMnE
YlZRI2qcxX5a6kEP/wKbPmwaTyQd7Cjw5pHnahEVBSndHlvfyAVl8Bga7KvM0xwKTawa/fMa5DfH
oVXGGB8kxI84AdF4zyDaHYBnUGmTiGkvMpmkoLwbugpHoNJ4ddYZrG5syqoH5LX2jN1IekLuZeQw
jxxG8k7y/5tV495OS++ejb8cg3UD8X1O3BKVqrTZqBP9qo/70Uy2jWC8yOx4Pb9NblKl+eg+isko
XVvYjW8QpctcwfEWaQAxG0XnYllf7Jqa468/0tmr8dNIJ/aSmVCWqIdsccraAfnR+ol2ywYfal3v
PGVt1bZm2sn6Vq6VPapm8RnkWOY2rkOX02Wg8TIacnKJ8n+TCUxuKU9HP/h5VBabjUBSRZpBI4iI
oaLgwXPcF7/qvVlOX0EU6/JcNtL6erpaOiV4xUTF/bxU9ebbMw12wz8jCscRAAa7a9ndL06I033o
sUA5bb3i0Fih1nOc7ZgZyFDmD/7qYacgvOSWP/u4+JBxUE4vlow2mv+hQ/sGotZRBICvsjJnx8h7
T2ecfdlTyn16VYhHFGa/NyEYcEJfYwJQfp8fS9JIhPy19rvR9/h1PgmM1/jwlfxoaXlI9DsxylsC
4MFfVkLOuh3J1fMdADCqnBNbmAWwO7v9r5IsPoxsovZx3bLK9PmOgvmWf1e4lEjGNnD5eJ+DKMQC
QriaQC+Rp06Jegdx750W3xlpXKldSi3PZWn635xVhMDOK3Mvk5/DOMjpTy9ipBaAFKhGMUmOEoxM
SGi2MCZEhxPwEvVDKccw+2BMhG9MHUMT1sXQcns3N5XLcvV9yCM+hoyEqgGZaIX7D76MBKIeR4Ks
pkve5fL635OYIh2Myc5mqxfTL9EnBmvv1hfYRSM8CFU49O5Vp//p3l8sAn86yfVDqMJh1G5amtuW
sFGI6l75JYKi2Tbd2973U2inI8oAebtqSJKozOd9FWQDksP4KPJRx78eG1Svr2h/9zRxcUhAUBCs
lhT9MlgRG4dZ/kW//TmYwbcIKevHnBaUGVluX/f6S/CoDcm9zTh6P3M8XsSbAIwk6qVTk/FYJWem
rz87xo+0Pkq1cUNaZuUEJ807jlgqX5pdGN7apC8J9DV8JEDU3sqj0XCKpidaKa/OPPUDk88KRwWe
X3RIaM7cLVhfC2h3bbYv5x0RxxeFjnbJaWeFx90yDytbLqW/VCXJNxMxmNQMllHQrgFVjnVouEtk
ldNp+/iE0MCdxO66N63maA0X8HTGU6Soo04ehnOQ6wunsKIVgoyA+bVBCC9HKpCHwlg8UMvzsIBw
jUpGtCIY7MyyDTtT/oRljgj+VGDM4OsOb1enB6v6JhHULfdfq4I+H5NCiUEdqxN7BvE+NMpemHV6
OP3XpSqtaEvABiyUiXwHkN3KQzjRl9qy7rj56yVtFhYIfeg1FP38XS7q1URHWP/gCfkbtyddW+cv
VhAdPWIM2pPRL3pFxCKzYM39G6bMLhTjiizKi24VCBVqZs+e638hBi86K5liqAPNRydJSMXttbpM
32KzxbT3YXPyWopDFvnTQQF9f7K18RfERMuasHRSDlblLb548KnNzlDLOjtc52FqmtFVhOhwJvN0
Jd2WC+0dlJZV0N2PcDDkWHitGcH++0gw9cd7Ff9M7P//suU7XjaG8xrr9m9uUxwlPovODbB7lL5i
LfMR84YN7NLizNFMl2C2nvtFc6asTkVI0QeGgZwPbNATFwCKUZ105Lpf4d3CzRKabx5vrIQ3YpPa
e/S7baOhiEB1yx2MCGYiORWLRNstwZq3W1YKcoy+nZHSzW7hsjuuW+95xuS1H6/Ryru6fzbWRB0O
ok6phEQI2HQTPqfByKTI2rW5eDbkOh4YeUXahV4US9VGFEtlOfAC0Pwtk+nK43Q3OZma0itvOrQx
0di4cBn7FW+b+0qwGcokR+05MojGQYKZt18ItME026P/RpsFyrrmecHseClau7OwkBo4sy80S4Nq
UIbZ0lvx+VCx7584jXQ1J7ubc4/JWj6rlUoDd+gfXiGMgx/Q+av9tWY40NleWrCGApAtZ2j/IslT
Q2KuBA3cKvcICTDUw7BUEsCLxA7/cV5edKZl18X48WDcifzyXEaIxPoJf2afIGAZ66qryGE5KeAA
MG1poQeEKephLZhBQgU2ntXVd3gGaa1QeL159aWjyVLPSwx43uw/KQ9bdX39ZdcExUNDLan1hcTO
N8h1mHvniWfnRPrzjkRAhGwm1JjjuwgHH7OX0jd6j58oB0cykM3cMNsEiNEFMbT3GHmDYCkENcUN
psnU1wzfclB07BK/vl3zK7A5oA9tBGgjUaLV/kHUXNkekioADodrMIPD68j4MFcpVB8NqH2/RQRZ
9ptrXOsyzm8TmCnH0yGmPYXppERPMZFU8gW4CPkmm4p9sdX3g4vzNaOYWxWM5wMreTPb6i1g7wBV
fu7/csML+Ci4CRNcA818vAauUUN27kCNQRRZuoil97h3aT58f8n0nIewe1gwsXJ6vvPBSzRvc7l+
9en/7ZFwT89aa+xaMZbeCxWV4b7DEOXdaTgs33VObtTpCOyajNy0O2JMJS39MtO6NiMk1v+2rpB1
io1+bqJtY1a9SaRFt0W83NEMPnmLHvFXqce0LPKGKdDGfYMzMN2yXZ9f+17eM72YqeIhUJOggmnx
bJZiKOv4m079rCfsRnNwkH7QFCsAO+Msi3nzcUaps7Otlc2f1SGwc11drnHeQe8cpBQcJF/8SHC6
mClnjkldlLd7QPWS2HvTvbMhvHzJT/zuueWBQbonCRmnl3Ce3iz0Ly7mJSFGClO/ukFjiNUT4a6N
Y73eCXmwxr77WLj8jif8TGFd9zrjuVLFAug+nIxEswnGLA3+OAoUi5H/+lChhylcqhtKXDkm3CT5
2BsIJQgTpW5reo89vnbApJJAfHZhObEnOZhxWsiUa9jfeFPSJZJsxRA4LYMGaJM9ZgtkG/UrqmyR
1bcw0V3Zv7OMrcskzl+AEyyKjQ+CPMSxyXqDhvCJj+Ym/N/YDaNFmyYMr+mh6ASPpS+tD/gHVHaZ
fe9gPKb4/kfhtLy4gi5xY9T7mu7Yo0VgqCnU3mGhE6HtrCZxOrgtV9AYgMy5SLb91wd8xCq3gm/B
Y4Tn55IxYjUtKKZlpS4xtyPENaXBqEKxRyUNjILNDgBjynSslKSnOHmihCMoO6AHr4qOGo/ahXwL
Vooci4O2ysAz1OGDx5pVJEZBWb2k4jbHToew5mMCUrQpGTgEXGJR9Y8Cn4LYRokUv/Taf+ZjnOc4
zJGbibJDoMbQ2JIWoQYjisjpXtLJhkHBMKr+mfU1iTVzs1Io8dORQ6Hu93tX5w2rhd+8F8nkkZrm
qJZJPCWjJGXHJBWUGfZ1iXsoWeiNEJMaGavcuXfRV1xMSjbBs1qMB/Iznfc3lmMatwoU0p044Xvd
/E09nSMiRnqzf3nc+eK4xHAJOmxjqK4gy1dm6FZrYkuTuu22umNqZJ0NoUuJ7uBppT06yDBeRBB3
BfeSZ68V5ppr2RedyNyizUiTuJP/G3iBUAsrdHgQUIPx3ExVb/SJOV5hpZHiKOyS06gXweIH0dQk
k0NjIrbXcL/XMR1zyrPdsQvbIoK/qQED9DgLMaCZGw21bNdYuKALS59O65X9MMfYYIf2VTKb1kIW
psdAXjj64w5hvTJ/6ZF/9KV8alwMw6uzYx4DEtxWhzjNwFPwNf1+otSO0Y+qZ0xzb+Z0xPDVqKRy
GweNgVjNX+0ZxJ0bhff76eV9mTpLPERGlfUAMEDzsYOFFYdRoaNPJpXeZMiSgq2mlv6xt6+V/93f
kyYLFMrgdWXPDkSNnPYxJpyIzrd3Z96jVJN3zbFNMGwr0isD0mnThnN0L3qvdVV3tgWJIE8L/LNa
og0LwyhFqXLUHEeApMjXcZy0uvZHb4ejr3pz//4V9deW/PtVBVqWzJHTC72ulK0StGaqv8mxdZvm
Tl+rJt1Z+kSIlgKUXdPVe5WkfA9YpQw1XsZ39b4j67NjQoJGP5J75u/JqCVT2KxH51IGxm/6+0Yy
WGNtPG0f8cDEJdUepEOYRzp6+odH/0cl6vyBQgcXl0sYScHYo4hLhwdrshzxfZIR4lfpHmIzuwW+
npSfyJzSk8wH8Li2bqmnGgTeNw304ij/oN/xVYbEbaET7U6yh5oP/5lEwQx5GON+FWQ9ZKg3lAv/
s9n3ATB7jUtrDPqciMmp+sYRE+IAKex7B9jvvB7kdWs5xPgRLLbq4TVbKVpDO1D7FgPov4g6wNhr
VIN6I1994/o9WlIvvgNL3DnjTxlRMRZpIe+Stkr9HxRAIGFDknhyhyle2GNHR+Ezzk5Jn0d/js1b
kVQON7kpQfk1C30BTtEn7v4RbBAW97FVp7umzhCnea4n5ScrW3XRgUKeORXgXDVPFLqJm9kAO0Y2
LonjfN+WQkSWYxyiw4S0wOWdkTmy7eatA8rhW1Bjb7/Ag+c0ACddDFdYfru1U5WbfnQ71WudAOub
MqRzp7r33pB96RGIDwIQHSTEwPlTTMIT10QeLHM1rzmBqO8Bo1hleox4CADnAr33Rf24C1/Lr8mC
FGH8njjFFwugNpt1pEZm0K7u498TIzVFFgkOMIzl6Z44/eTr0E412B7NYMfYPfiu/NiQUNd0FsoB
ttYTyLyhA/StWOh400Yvo2BSfmB9RXu54l+0MUMeCUb6vaHAk1zpSCVwCpAKPh5J+ZymOIDCB49l
CSBv4ydrRzQn5BYWZlttzU0Lz3fCZsnGmxevlytxss7WYv4acU0BxCd2m+3zUXOED4MS57H36QDL
vDmsRsucwLrd4D/UzhfxfwaPm71JcO4ClwZnHDneNIEDK/okZgNRxv3bU2oA0+Mvaa76RTXqwUKi
hy/f5tWuUFilSaAXlkaFcmlXJaxgtSDYEqpRk1AxUNGyqGT7tYFiy26Sji54PNlb0kWQl8S+OGhr
89Z3494oOh7em69m5fohFiEr5wA7fiR8y3OgL0eLLF0h4KQ2BhB4hGXUMCLZ/8YZR434DbtvHy96
Le+EyKJKQJIPKMQPGnQ+7BLwZmJSlmg1QRxlnBg0b0uH4/X19UCcOmOudglaumANaCrcld3Caqh3
oQTwG5do6+KtzbVm8jAzorqqJJFvbbOaWcmay2bT1pupF6QV8dKNPV1eaXkz9f9G/rMBDVL9PURY
tVNFgbuQFmVI91NsKlzVAzJxDtB2IJJgVnH0AJRU+Hg/C8o+TKIKqZaZ6RNVhjD1YnFdKwozh+2a
MSBK4IBjsIWJe8zb/jVOOrqdrS+LYDNbdxS5DJIM6Qm3j/AtpG0ur9zZwHywH9/jsyiUEz0TsDv5
dTweXprdtmWmJ5whRihXyR/NaD9KDb/BvFPLpmhnSOwXmQz0OKFiywz80vL7Xal+za13NCOAjH7N
iMQWZO1/0sA+Ju7mqLmF3AJfjoXQOvOTh633FjbK9+Shn4IXSh599dfsKT2xgdJ6IMY2DMxlbsjH
B2u39liHay+zUlvo+NBNRJStcsis8vjYG7Xw1zn6388A4/faN7ktXWBlKjrd6Q8iN4/eBUb12LEf
0iIXp9H8QtV5ah/9TXImGT0C1MMk+aaNr/io4ogLa20OX6BftHidoicjuojP/sNUW+5Wou38uez7
exqYNCOK/3LTwkDl3naHpl/hO7uLN04DsItzLQahi0parVeOlhlYAewpQjLIucEdOnURh1XtBq/V
LTRhZ6WrR6jG5SM3B2zNzF7KsjYXDFwR0QBrrGceVcBPJQC8h5lt4vjhgs6O7UW9Oa9VloDS7doA
S1WI/pdrRRBENTDm7m4SAU3H9opBHP0a4Jiq1UIKPlovV2dd0x3yP9+gz2FaGmo0aj5URsMjrcH0
vKKy+kPYnZIbuvPJIjjx4R76o7eXvrLK2rc5T3nTh27aVMXbM2cAK2FayZf4NBy74sLAahkKGkha
6DvaFOer+C5p84BtGDBoAGz54Rc5FG4Uz8KomB6P7hszmkPFziq/mp7HFdwyioTXnL5x84fdHFI3
u5GPht1VhhE0PyNkvqodu2nF5q5Qqzp94WKeSaGJTn0ZLfsQyfSNegMvBXS5jjs/iw1YU3Jf/Gaa
tHI6eabblE7/SwQO+gxd0PofzJwofkslz2lDD2oI5Jzy6rb7FkCZ6PRwpNHIIMtnab4L7xoPf3Lp
2EDCSjFnP8WlxwALKFxrFZ8NCt5JRgmKrvmhUSBW3GHCVmmxxS8xnaQeoxPpPQQlKhBk1uvXuG3A
7Pe4ppYrxpPLb0K/H0FW0/eQcuFHX8h+kCngiUwYoYxaEjW+WsmBb/USTs09muqjx2HMY4vkz81W
orrW44toJJroo2+gyvtBkyhz6AiaERjE5Kp1MHyQJvXJYQHmvA+pqE9gVuATB1S0mPVYGRvRNv90
dDPLgqwyWd3sXDF4yZ7rDTQYjGgoJ+r+FMnttN6bmEujW858FRH2iwyS8iURWs78tOurIYy4YF+U
GstMMRE6zJVJDRxhsUqTOdQIXfMnv6TqOADk+nLxLg6ckzvb3qXYe+BEmYiotRM94rNWYzBCnmZT
L9GfT+yUh3Wwt40la+pPps2dn05Zbon3NBabOk9ZL6dBgM1lnTSldpme0JhWlEnyZohr1/wp5qus
j6QkYch4SfMAiehbbTZay4mxBAIaa+B61YzwV+7kdJX1/Tw84+Ew3GoEId8ZOaN8DzrSDdeVHsZs
/Q+422GLrSYsKFhkMIzzBbWeaPLIYWaBKkB9hX5o/6DKooSPY3UG5j4rQVlWlL4vp8OM9aDkycR5
Qs7GW1tUH3a0fWCQwb41OMB1c97z/DoTDrzKKdH1JBPia+Zkw778kMHKXFxmsCyP4usx9DMKF+A5
ezFFdYd88m5FEaQSGjMZMf0GcqTsZx0u8dMxBg8ZzUZHNQzhPB2iv5ZoxhufpXR4A3pQzpGsOTkl
yb6PRiQqGWGX+3LZzzV1Xh5s8USFlBv8iIDLTx8YzO0dlGPXdzbMBzdsE2nQZyIVAd7Yu/hN29kH
PKVGv1mMbmAuaDMksGwTPG/i19DBkZ19BKpMVRSAPeDmIDZI+4IV++dbXIRqAOtjaJXf9QZiW+4U
rn+bM8aUKUqshGHlE9yJ5Lr+rzgQfhcpAUiiwxyD3WMMW/7NC6TEcYxW4roTtQOjUu7CzEZA60DZ
K+vczyWdbjK55dlJIRsDAvc02lfsOt8VFB8inCnUbomGXkNw/RZ8Aw02ocqQLG6a30UD5wt/uei+
czI0gezoC7KI3RHHdFmYRonTIsDY/uN08zi7Blzs9Tfj2cfNPJokckXNkeIa7/GnFiZDY8Ht7a3F
i3K9x+/WECWZiUT4yePLISVNc8yapX9J+bZee9afHqje2thY8JngSLHOXfI8ntBfsxWJLph7NgTd
TIVOFbK/P1msSIFZ2h6jqjq2S8tDoWklcxS/9INIsC/KFmL3iZq2SZy8dWY8eaIbeLrFedy2gzaS
BvGATXqdCN56Zx9SyPhX4w1FnzuyWIQkGvyoreaAahehCGTevXx+OOoDdae2qM870b76/jYTSuTj
0AouC3AlmJhTHCFAplC6xzDmeDes+X7dFpMT8/iodb8ZqIBzI9rEhA3F0KWrNgBATvGLrXDoS3HJ
UPWiGdtRflXwZFquBoqsw3ag1vGZSQ5UvZ9rezq1I4VohZ4Uhq+PQ5hFzqmzTCHcrYKtTEtyQsWg
91kzN+EgZub8MFxGT8sMkisYQJoAYjMGTyx5a9FWflyTv6oIjqPDE6NAnAg/HQWz+FMboen/KVYr
P4/aM0luzNEl/gTqTuueBqs7XHxpHhz4t57BuQ0hYfrep5KKrMmwDBqnSyCbk2p3D2Irb+By0tXp
4CtFc3SM1lZ0gRutkki1Xic76/4ugd9//+XyE9a+/Vs3yvMmUBdiOCZkyEu8+ji99Tzd4QrOjVNa
MKNC71pSw1j45xgxz4GBJRK+Js3TLlUBAxsoeAHbyjAmwzGBxG089nKroaw6fVJ1TivEzaq8NSqh
z8pmDFHEUS5mqJ8X5o+FflZXZ0CWlbF+qymsFP6QLKsLKzZLUKmMRTOKWOjKS3M428HLYcy0LJDB
x7/pChKDgZ0U7TlEZi0wISCayuLsZQVQz4vbe0kkDgMZpNuGk04Y2gX7i908rJZ7ilIpHYmjGyzJ
n92dI+TD7dYsvYQhOmTIOSZ3n/8FrsuficFBM9exa2uZIXmdM0fsjwNVjhix4XcuMfICw3xmaMo3
S4ghCXvYg53baHfYv2Nho+YK1xVME4v16E/4dixM/Ez1joOOifBCJ8hUPaYYkseQoT2j8SEGF/vf
GuS+6LyopZh2Di7SOxTYXce/oTIfe3v5Q30AKvio8aR+e2aHVfkFSzU5dsvDykLvZodD7FlwVSjk
nZszf0rRzX3rri04JH9SmpaIvzb4925LJNO1VYB7BCjDxc3f3JSssmEQsgcMNTk7JtIsEexzqtEI
v2iZQRFISjqGHcKLWkmIKFchA3cF8sZohuWlHtk7oOkgrCAUiPPn4RLrmwuNlUk+9nh2pQnFpKHl
1EOf2fa38PCC93bidZos/6huqTYxvHN0moCF+njnYcyALKsehOAYCw6sF41BgPA2Ik/Vnfv4dB9Y
Z46p57NO5Pyt2rk1T3IcoUkJmf+9NwawBbx9/d43NyPmpRuo0mE1C9ndFt3qEWkNRZBy/twyh1RV
lKQCIsU++AeJhgSpIjqhZN2myFR07wBpM3+iIIvNifZJkPGMfAazvaPKsLxqfYxn2a7ik0z/CvZ6
hSabthH4Lfn0mRXvLC32gGOKoZyIW08HDUp9kM+1gB2Hf9SkmqJNMbWk+rb74lsF7bhqj7P0ni33
NWTtCfT4ZFPEFvBgpBW1c1CZCMtjUywvwyifzhKyJkkVwyMlH/mvxa3JeVdt8qGNK3q4zYktNRvV
D3RJfNcVDA/2/POAU6FsaCxoEZYpziGaRFCVgyjITudlzaOimTG2szzomePZ0olE5hyJfR0q6LEl
pG0Gts0DNpgXIN3qQprjNQ4lNsU/7nplVozWYFmCVrHyICNKqwTTtDLs309yjRm/kncgSRoM7AsY
8AXHoY1t2eoQ6i0Ahr0DC2qohZZH3VA4V/PXdqIM9o8ZEcsWmEl9cWkUUq/k52RhGc6I/av5MKti
ig4Wwj9X6XuPY5wKrARAzJdkAeDiG0MOILtIGzxBN+qVV48pWSyhWEzpwlcILIoHp4GZqpF/loql
KBz6Ppsmw18mcjszIjYLxDsqgQXq5wecJxa/PN9c5Bu3i28mRb5WQDZweMaqlb0jsDiZ9Wg5qPaz
noolKh3W8I5mwnssfteBRe323/IYuVbg7tcPn0BA8eR4opXsk1I5aZMEKBSkSIoaThzmQFbwfbXA
JYCg8i/l9seHq1hsGOEjUjFTtKByWguMM6MShqCVUliXg5poCwUMsMnvHEPwLHsgOH3lMArz2EWp
EDOmbSfQzLryVpobgZe/QFvuLt01a0KOJUChuKi9mrFSU9EysiGaX1WLXzVvuiiWOd08Wuzy4LmR
u+ZbYk2QrxbSFB3hfbknHWF4K8BcBAJwGNotwnjnmgQTmnKCUScPI2V9qSYrhgd7ORpPRHzMmzyw
U3NhOMocx1uLWu9kKWbykCmOiGXNrcLhhTfgKAWR4x9IuokcaG2QDgLzCL8kOs6KMxFIHxvL/fKC
T5ogrJGNnuvaQ5kEOjvnsRPBJDJZlJ2WEoORm02oHyZF0deXfjUr4HdcBB7AfXHT4zkk+FK00TYd
64TAHrEgfe8JwyCuRg2A4pB2I3xtGWtESUoX949Ty5+hIAUgXUgsS6ks6chPlVDoSBimQQNAezfB
JFg5FnqOULaX0DgbLFv9dBDCoG/IXTgkg8+W2y2Iwtzp4ID+OYrovZ43qvdaAHn7VFiVbsbN5gEF
e9ddWQVppsDoQ0YadJaSHWc4Pmlm3EMaBobRAaTFF64++RbSS28pbrLKcZYLNG24RLy/FC2YgcZM
RjGjxNyPNNaL7j4LuSQoJdhzZtWllTTNlS+QQHBRk33PMMPZ9YpGQ3n+L+o2CpUJFcJKjPTyNxyr
qbbgUVgEwZgDKqGxPo6QWauXZi2Le44ULF9hOkZpRXxamyVoVVStHg10rz83tKzVD/qkhZkJwipk
Ec2VGAgNb2wixqvQh4CUzpEI3+OTwt2VDsbckIKt5Nny6rZfEFYRO5J2OlyMAUccnzcyj6DxchDZ
zV9+122RW3wNP2vPW3+34Aa9AF9e2Rauk4Ube1TseHx+Ko0VwwcN5z5yuvXmvo/DUzxxnKdlCaCK
HdTiAKh9IHvKrGYP+bhVH16tzh/DqU4o6DP0Vcz/HKT5HRZUAJYasCmk1Et0h84MzVu8a8PIuUbg
44UegSh66BlDoKYL+bFUlq5ETbu/bw6RP0ooBxwSSjQ1Ma6+m5wztTO03Rv8uJevCO+YjgBzI7dr
0+Vrcmw4eZooKy6wOSu+gCtr9M7wU5TeeEuMXzydC5RKxMRtBiC4dqsgTOmZx89stVZVgf1kIJHo
6GJl+p7ElQtBMs8zUZspo7GOVI4mFa5zo9jHkz69WBb2jd0KCySEedQpGGjSalXHaOb9vif3k/lH
yZjkpiRb8MS2sukwLyHjgv8M5Zm3b631ciTrswP4kgGfoAWtiJ1X04At91VZFrUcWrF6gBauYRDV
rdWgraaxOOMS5dBtFRQAJjgPPGAVZyQuEEAxZkf1WXFzN6R6d+EqB5qI1z9golWN+XnmdRCc2FTl
K7FN+ZngDzEhNYaGheHwZ5Ce5Ho52BuBeqh9UerMHpHObKj/a20a54L2YBmSASmacqNxroZQ7Or2
V/i1a9GBInhqJG+ZVfNygg7ZcGW4vrvNqbJ+VBRkFITvzXngCps8by8pyiKjej/KvrUxFCAyQil+
uuMK1K1PlSnRWJiXznqf07U4leq3gYlHn01DnGNnAlfJBBENUOii00e1+zpkvVdxNPkR2nSoxBj4
Xj94ON8Qk749Lpzt4HZgggo3SVGsMoRGYTNtx+m1IpAV3NpKeCUUaI9YlFjahm3V00836/T09qaz
gP0dFH3b3SULS2acXS50qwed+cApUyDIdx+OWsO3oJICAweYC5YW0sYidOA8AdZGncbRa1xax0Er
1S+peYahgwLjdus8RgpkHlGq4DRKsKvDbRTL+B8iYbvrOIfuynWmmbaoqkpmY1Dh/4+L4vOr7NrB
m+6KIErlcjIxc4/xH6LqRLLtGCkKPDxP6BBtLT6BQG64v6ne3AsGVjNnUlctLQ8aGWYVY5+2bkKn
fzNeDjHf4/A+4vQZEqxWF43FZIkz68sYmw54WsHHTAhfF7C6ybLci/Q/eo+Ux7XOQoKETqz4jXCI
jN8fQkeUwRaA9DeThkhcrxTjHv8rOq50fhczT3W4O8FUHFGxNCoiqPKdR/rWQEnFJliV5ZBiPVnt
4BShkiKEIrK2QLT1eUFXobzrmEz2xUI/MegF7I6Z3SKp7RFIn/EruVu5I86zKYU0Y9qSClv+/+8T
fZd0/O3yPXzmBH9CbQC5cZM2VqZm0Kkdwi4Z+QJyHZ6+L3wmm0ETaOS9wnV0p+a0SnzkL06IvRzJ
6+yeR8L4l80jl1L4GCEo/c24/5SpM1LeaQo/UjNEe/4YGaG5BeVv4FoM7ymE/OqkqFkrez1d/szy
R5/8m1aKoNshlNv0Fel6iKjsa9HeYKuMIw4Lqh10JZRG3rSZx1x+pWJMKdmoqgWTPAR6oQc3Xya2
qk2l1HgT9Mc6b874rODY3VW/RkWrcqgGmfkoGbEQkC6mz2hBofqnUysSDuJca/HPi3w12Pli1fOn
OBGq8/g8jI5VO05yv5Vv9ZGl26DK87Q2rjj7qBpwT2kZv37qwdLHBPad4KfwGApdYQ6mlTPKpfB6
wkxzXhgsTmf9j/ZUCD5+244IXAiYzkAWk+lrKl1Pk27n0dZ+EMfosJP2wrl0joDzUMXIqu1s7/0G
4ANlMZzycbNZ+5DtjuJo6wUuzwoJehGug6f6jk+0IrawlcTfKU4Hwi+3YqFA5OiOCmZx73xb/127
IsPyxlWwLS+TxikePfFl5oTF4cKIVcGSAQJ+OraRq2yIDR7XR0l5TJ++89o9TLmA5KmX7keJ6hhD
Zc2adUoIwCKI9jDHzyQi/ytSFvRnWKIbOT3klxrUtfkqPCwPegH/83O7/uewY2X3XI0qDiH9wZ5N
pWeHz34GhLPk9MAbvLn6r/0qMShR3P4/gfIFm3CXG+e99sBWYtA3AIyJqVT3xyBGUD8ZtsF0md/2
l10PfvydFr46ejkrMXa+TD7L60ORl93VKmpajtvXNu+3knVWDBwM+LUWtVAFmhVHkI0qqvJrCmbs
UIfxxAN4NA9VOQoZtHwq436PHDVRKcvbL3CqRXpjYHEvU3sjAvLQJ2+Nz10nm5/C8p2YCBBhqg5K
n9lMP+Nam0vZppjIXw0YbWaVAtLA9+D7SS1vPPIxVW8EGhLEi9TEQ1U02AtNP7I7iZBAlyxt8L96
jXd1dtqp5PwsdcZFkchG5BtjiJAnjnO786eW/vG3hlXpFHCX0uA00iQvoZ6yCEIKjFav9bzZO8rr
LwuwFY4UkdqIsN94Rf6LQKuP9tj+hOt+nLWU8afnipO3XV18He+H7Nwf/odG7GRCuTiAMSt+2Sb/
PlDfGI4cqPrT+VSSw9xuhFwZnMXUPt9nWKJmBkA6GTYYTW+39/6fxQL2wfLlO/fha2IqcdzE9Rd+
6B0WxC/tmRNO8OCLpqQ/OIp0C0cPJwvQFUzhC50Bu5kkPDA3YJ1ywsYBkD2BtJP5FOCemQHTCnE2
wSEJWUAkgpXT+9LrA0NLNgdUt109WpTdLjc4vO+7cLHuCsli9lmyf1YgV81MntaaFcZOV0VcNGnt
QGgOlGSoT/6w8C/j0Ge1XcVZ0khK7X10Dy+M1UbeUu17Ht1u7kRCy5RgoEZSWl9slcCuz8WJwHow
zemTjS89tycRVNY8sSh7GjPMIFtjwAoFEvLoeJ18UXqdDzOWioNUgX4MjL7zq+/gjQ5JpH+w54dJ
g177BQiMsnm6bXcl3S9rdrk+FgjFaLib3MebgiP5GjmuRCg4cAZTW4gvW6ax9YyQs6+Zh3BeLJqX
k9IN0zlqp26hFTSbOQ+Gf0wy38WGd8ITjrd4bSTFs41niUNcBxZUxCHfrCRZST1NURVOVyy1Ls8d
yga7TrtQPYAL/PmxlxnDIuz0MWxIfnKSOoxMJRQn6SfXGKcY9gWQH4h/so8vPwsnBybcDTHHfNc6
p+V1dsT2DN+DyoZYm3cw1hyB49ZC2+kZmlNVDeQyCCAYryrMfY+rw+hiqm0IJIi2y55rJ+aBhHMC
I2X6Wol2ZNi6BTYpKFydKeGH7pfw6rWKOH/xPN29bR8f7KX5bbHdNsSYBMOH4HohUbRuj+xsWpwH
G7sYliaJzxpM1/kZPzTBZU40XV/y2upyurXE1RNQkFZu7RGFKNw393pv0DEvQs2Ag4EEtJmqMJaj
PuhSNtgJUpfkaKCOuOOFy/bAk3yL0jQ2DR/UAKhoMyOTINYaYJOgcVWaL1kShCHO2A+XUOwI3ir3
amykww/gIxwg/GwPrMvT41aOrADDIGWGcRycR8laD1Hs5rIn9YLCv9IVScPykAONF+Bp1Ct7Tmax
s25hlJ76qcyWqvOOHrZgffAm/iTYgovRFrURgHOntk7a5VpTyqH7B0kqsiGeFYH3igE39AYfBEed
aL8UQu546oXcc2LjKWdjeY5vu9Vn09ezH8WJ6BfnRmhyhjhJNvNpV4RolP18qZ2zZ/7eaKwFtv6J
jPEuwk0H9m18f+qxXgnyMbTx4qyqv6BoQwixEczc6YGrueETA+GBe3wTkjKyGkqQfL8zE6zZe6ws
1JmbGamMZeUsZG1j3RC7CWY8h6zUMIDECyt7zWRhvsw8v7aVBP4/hI60smi+mYasv7pGctBegwiC
/wWdPjhk1tMS13NGlmcPd2sv5SY2bdD3OpfXIOrVV5ygdMJ5DvlfpeLeE2MH09LUMhW9dl/sXm+h
xHY2IVbAii9LgB1vOg3QfEyc9Ul0gwEGwaAkJjsIL6tbXIgYu0HT5m82a7d7ljV9AJoua7kOgaVp
ePi+GL2doBmqhW2FtgS6GwHceQyEnvYW0OHaYnH1db+0q3bizgDnIzO+TGhgYn24/HkHJQ3HgRRh
8QwE3zpCMbw+EpZUwQyimqRMFA0NN7XZzoBGfzsAbtHd1xnTyMW4ZTQ7FhPixjD+lNI8gfy3Za4E
WE77n83HukiH/HDWPQs4EpGQjcgdzbXsbggzkwyTBcY7En/eslnxc63+lKgypaL1XjaG35SZrudW
cgXdcY53Eake1wQRGRcxaghZDtosL8DguSEI7DxGX4+1CkdQZIC+KAWsmBUdNMljWDrpuQtC9KQc
wa3iEgvPRY70h9EFnjo2CmpiZuEfgcRlKfCYNqcinQ4fUKKSoJ4eDzkyCatFpkFDaszdVdW1W8DI
CrJ4UvKy8UVGb0HC/xiGjD92ruxvflCtHFJoZ74OMCAXXJZnaNy5/hczLXepsqEr7c+lwSzqBnWP
P9RmngJLRTa+b8lGgstee+fw1oo4HHyA6TUcWKy+kaX8icIQRF69E4bM6U0b6BI/P9v3PsDP5hEO
XY65SN0vdzKwvMdt1FFZ2piymLX2WCU+R9+8ciMFCPcXUgHwjul4YrXHPOVbk878bEftVCDpCCfX
+Xpl3mxwYjpqf9hHvkpL57LK7a2S0OVcHgTnhN8rcjBN3isgO7QxmBgnBGYLNldMgaSTvhYyFuiA
/fJvca/gRevHr2CSbtko8+yJ/29r6rYaLA7j+hBviKuS0lUQ3LEWl1Sf6ob6RU9HQO4OqAdLTm1T
WbTDTu+Esof8govZ3PdAo8XluORKOXaBlKHaWf3Vu1YWI00xWstuGm7JNG8QuosXv10n3u4QYJeA
z96VCT02k+PXCp+ahh3BknwaDcIfinCWEVI+Lyx3ajnPmXz8aKKdwFvHjlSbv+9e0+PPHppIQpbe
1aWBoIPmvPrrsZLSy0ZHdXUnULk+JO4WrBzvtHRiubbXkl+M+h3IerZfa3SGMovYLnLZZv+4rXrq
blqdiRf2ipotSW1L6ZdsaZ83vwge/kb+u4tZyYXhlZ99QhrzqJFyu3E0pZPwOfhyRSn4/Z+GjlIh
OuSDHajoGZ0OIYFqG0g7G0qrH8539d1FA78Je78il4ey2e889WV2jXz2D+bw1bXBRGuaXRom+GrJ
peTjtueF4Fv4bQkTzuF6By2mmQDpqpgEA3RzgUlnQVqRvk1XUuC+XLoG/sJ1vjahEI4v9OLW0qKT
jiXsDlIWwLni6yjqyzBOxLBqhycvy1FD+oGqWAxfN2E9OHXzpZ0BLNxa0xZ/S0E2BcekeO66gIZH
6lEQQ9VSrJKvSEAJvnPB88pfUn+39bJa6+tH3LM7xzHc59MVsoH/zu1P/2vX157dLRACuTlFWgSR
6xDa8Dh+ylrJiDLzaTd8CWeOi45YTu3h1CO8D8/TWNdvM/Ar0gJ3CHow1W4dJ3dfEGZFOohtBW7N
dk83viNR+mdPv6WOazUnZcYDaSIW0ySnYw6GVAKtAKeXhoSb3WO4BZxoTgf/uhCj6kT5gwUpOczP
hRW5lK4Cjm6e6ePsKiFu0yrShyVmIn7VKJsOmzH0NZFWFrB9vSXjfals0p3nzS8ZAfyHGT/GfE9p
046fXJegbB0To+lCJKIEhE1LNAX5k8gsct+aV19V0K/V4OEA12iRTTQei+mIJ7LSnylNcvLNWMjr
gX1HwZzUzT1CEguvgd2hF9trHx545rOJ0LttglOUzLix+5KkQQw6GaCiPOUCJjFeqNvwKaZQjUWP
zrmhjx4GK+wdhy32BHnqKxEn0LmJgE2u3zOLGIgOglutAIaGABje/b4mbD+TSp80wf0Q1h0m/FM2
qiz8lMc/QpBZtwSi07qNVwsljjpcpE81pkJOdhFE+YWuPHD4US9HblhZ+Krn0KoMk3LHgw30V1Bd
+VVldb2WUH7tjOYkhdIcttPWYti6nQTZtXK3Up85BPPSyTGjBFRL0YbNSNoZAFVUHZgKRgLQptxD
sUVRLyqctXf41GbCnt12Wk4ColrTDbicbSD1nnpJQ58utWORFulbxcaWla+cFL9E9K2aWhTCVvUs
bw5gs4hL9X2BiQe/qbhfdKCTPLGo+aXQiHbMe6A5fSw1j82HPNv+mdYRAhLatypgsU0LSMz8BRrs
F2zhRM1qEDBDjWe0nJsK7dvBnCpVELqx0hq2Ziq5kAt+r/AG0Jqf10h8OULwOXsufXzJQArfwbCZ
LVzs028PhMzYzOtRuxVIg0Ifi/MEkd99gUZrG/gKBuRLaoJm5LfYtsBD8YpDzGXMiyhV++aVPEoY
/4uYuYJH8gvGJiRBr9ldyL/UyGw1KQr920gnmTBU4pprPIduP9EkwSSrSKzjC4mGDMS925lzJYKE
/THI3HfYGfV9ct6wwF/RUiauh9TYTuToUgNyaYv8M62qubcJ/pg2PDXluhzqWrQcAzJ48fQD4EHj
TFRcKLN4WKzBsoYuIET5f66nlrSon/TJ/ILJjckYJp8bsHMrUpRmOsvLdXrgp4Ypg2lHE03yOBjB
p4BedTyP/rIm9Kx6rjTourb6gDNoDZnG18WTS3+NX6ceMTe9OknOCwetXOZvNzY1X7xP817fv71j
rGsCCUpT1HXx4Vovcrd0MVBHrwTbjTzvDbgyWJICWfPCuvOtr1G/A6nSG8ab9w1x9+UIEz1UcltP
y/YR/qjsbkI59h6z/wl9hgqzP1lF2cEs2QJ3ZMUeztS6y9ynE+FrP9tIoqFc8Tt67EbWxD0tTgCj
ZS7ksVVWxrWx2dD9hRWx6IT6JThrEAYbem+BR9GX+eGAZdWy7QYXwuU0MV7FMmv3gYmrQAl2r1yn
UxY2dqIq5YJ820Tk2xbCN2Q/WW/uJknXxzftmyCYiZbMtQ3Pg9+h7mAbft50zhL6D2nj5DFoaHEk
js+eBfccdMDmbwQlCaymkjuFwPqPWCEzGfDnWkc+N+/R+gYym/rT7dEJtsmND/8ZyqU/W6Qc8sk5
4O5IO1LQKbNcSTadKy2K3DpQgSQHC3FE9UfWQh4l9PzazwCv6RzJxM5vicY+Q4MJkmf12mHm++oL
iqfkaaXc/ZsV5V6ez4UBLUjMgsanchWFd4ihXoTpmDXUTvEjWn0w65au+WqnNmL8Mmi33ljjj2Nx
eleX1m2g7AYRsC1sKcxjZSjTMKjNA7Zx78mRGEEaoBezAChSU+n7YqSVvsSQOKE4CdoZ38Ku/QJs
FrAJa1fruWRVZucRg+yfTv9+vFv5lm5QTHjNH4rk2J2vCkTJ/S2mcfyS9U5Gq/VURAdlT3+y4biU
kuvHwTKrI0c+SymxPccP+JWV0wS/zXPhidKJgA3CjKU87JbtvvYF7STzTbNPKLNBNNE9h5ai0qgy
6BkkwRq5USD2i8lD83WblNOCZd+lrfTJXkNwgwu3Xv4ciwNOENXXcmjana9JnILLwXkxcsPg7g0O
KZTXoDpdYnJpj/2SmxTJJiUtDlR7fQLKvTScB5aoWynghO2sSS1m+ZEpMz2yJX7E3YhTJ8gcz+jJ
4TFY7aIyNkgOWIEcwtH1BEZzu4U85HUqTVdXKa/x2GebaWYbZGCa9rz7dqZ7fDPuCEVSnQGGil7C
qPbo2QpI+DWiqX7UyJz2GphX/nuRaCyto7L6obO76vkLn1lLg97jatCN2QEilEd8dn8oZbyCZnQc
bZKUnxsoRLDx1eqZ54ba+fBOJVUVXUHHh9SQ023TSXEPKOkDQOcgn0RBLFr120esxA4SmTCd7y0e
KX/y269bGKvAM5tNpuYnp7hGQEh0eVnGp0iT4kFR3hsXGaO/3nnAK96+TF2sA8udOx1J3+oVUqRC
3HuQ76N7DmyTiqUg1c3njq2Xw0iqiWYnH/6cTlSgJHMAbtZCbLzSTXDd4OJETSXW7xHlHq8ybOKT
p3ZndgmbZImktlAM8JfQYJlpbTBeFchFuHGEZJCt8XCLORdBkQrEbXIYraCbkhNx4PRJD6WfMYuW
GcGpekMdBJROCNZOT4XLjax5G6lccxWb8yI1S6Bakg8AE+ELz+DslJDRKliHaDjNR9XcqpVnxFQR
XD12ECtsQBacu2VBwatDh4AD3MpkXcwqI3Y0KR8X7FSdki6aHGdDEtEztwPh8KspwIdIa/o4Tg3O
H+COpiGEuW7peleSutr15C1z4Q/KRcV0Mlxrh/K5caIM/A2NULdWFQy2r+FrufMnjsTmj9Df53S/
YhnuHKdBGXAz5kKICJpr2F4gyfzVj9xL7TNvvFSrNftd7Du/ciEOoduulqgBVxIf/GBN0WU919k3
UwFPLwsZ2N5rX1Y4f76kMQbnwem30E4VuLxPq90dOSZrRbA9odeqk7/j4XK0XzyAxEh9TKopA66b
87cEzNyRS8LipPSM9M7TzWeXb26ztk+v6haSmUZJEyeD1cpCJe60w8v4OLZY5cNAmYYliEvtF/3y
quEN24IhtjQk+7WLtIQjucqGJEFWprCPNxnKSRoaU0PHzcu2tsca6yc6REKc/v+dqmZOy0rFSvEz
sa3XKv2W7dcqm0+0o+zKJmIvEpXgs+XCQxw0X2+A7qKB5Fr96ef4hUvyjgpPZShBWGikdodo2XlD
f0u0DVXuqXrqSTXPfJXoQrodFThDgHdLXm2oOTJd6PRAiFBJy0K5mm4pPNAwhOgFuh8mRG52Aska
bjy2RRkUBLzR+CwpOjnNTL/1/Gy1KbSTLQRlNmpXwtodRPFRKfdUapaDoi3fffXuhhWBhRcV9yg+
6we7nJtkY+gGjK9aHBf7q4bb+O9/DqTPklrhwR7mgZZrm5OHdkBuLqrNqnlmr+1ejh0zvaZcxkn1
u487Vbp6r78CFPnZNVXlnyBmSfO9dnoYi7b+PnfFOmGM57oS0kgFE641yL/mvG2r+gEF+K8vUw3B
S7a5yTofIDjdSrdKNR4uNU2XDRNZn2Z26c/kY+bSHgn+25Sb3/+iL/cI8IwxGJmI9EHEFKmhUGTO
arACpLQomkQnC29SJzcoBC8oYDs/9AoKc/5YpEwCPZz/Nx+fps4p+XFAzRE2/RlUG5FW4wvSBqWQ
+nbs9DC5c7ZcCii/FTHWjGDYsjMmn+ya6lwSI396JWxaJ5GklQXmGdoaVnT+Vhi2zvE1c4eZk8kT
fA2Bj9UPphWN3xNwV0nafGLI0ccr3LukoghvHIUWNiobXBMcoK7699u0qYW8sFsyJxvB+Ca7kqe8
NobwPZoeHLpZCQXSPhVFQpVOA+e123ff1vCgRmlk0gYrlugIvNw8G6MNK+aydet16n3W1XusAxkN
lXDobX5P+scl9z70XYBJW/mEf8HvOvi56hEK7o/twBDFGjxpFdEgXdxrcW3tVCsA5VdH71FSjBv+
Zz9WuRDURv31CYwo07ObDfOKemITQKPP7OIMv2QzXJvZqU5zBntIdtpDBItswlkP2zDrXAUOLDFT
vE7XV+0P+p2cxdH0oAc4efG6aYmGn0LUZLhe1mK4v/lifCliROxmmLNayZUMh1QJ5E6CMXJA/1aA
cv9NbcDD7Z2eMsmur72K+3MYVPcQbLRhi9SKWZv6FsOPC7qWss4wr1xJK04z2vKNEf7CrGX4MrXE
zBqtVF2f312U5Ax1dbwVvSrlQqZ+XAKLCUYhwdClMT8CabDq0p+eFWHXYpxnt9I/nGbU6WilWFIu
8BXhe0mBl8Sy0QKwCfJ02R+tzMuBRekkaWA06Wswy7KWOdsApP0ML1J2gOH6ezfzFGspNthTcVRk
sW+MjJNyj7YfAw7xC5nqSTKFLx1D8cnsfrETuVQxMtdCumwInYzAtcLIRVzyYYP+9bXBAQfIvsK/
KhhgGmADp17uyvOkFRxDad2QQSTVErmEyNVAZqgdp+LW/8J8lSlOZlCUU30y8cLjAk7yqphqu1EI
zUshnDeFDFu2wMTHaEMPuz2uX1hmbFU41+BbVXs1HDapbmEC0sdv8wWdLTflah23E0/Um24swZ3K
Y6x/9asGdJpLEoRWtx7cfV1zCvFfbzR+fFIsmjONug/elS4n83275SrFeiPhW82ZFDSS/DaeoFTM
P1uii2uWcTwp2jwV6dG/g3CQ5I9pG4shxKhb5DB6aYjLbB7SD8KKz+C+38x2xUfEPXQTxXvwb984
85Q1wD0JH97S/GCfeho9Pba74dRsl+GkTh+1733wYcsntWtQYbDQvGUEWiGH+fCcsaZ647GLwMV3
HGXSV0B/x7fLa5DCDYn3q94kUL0lxioyBDHM4/s5BywsDBGcug883zd35Gs9iCEoRIbckoBcdYy8
a32jDZrVndSNqVLb/cb8SZEO1t6xCk0AQQ7Fm6U84uDGkP1UXGfN6uB7f0pfc/KRgBFQ3FJo8un+
4af7zZ0XTz7J5YnzHD0EjyV3Gsfs6ivKYZ6XoccSgYoASKbDDjcyDTa4fWSkyYPn3Mr9f7TJaZYa
tlzGaYMHCEUCUvkSSVnKdmU5dDW3mNENVEcZ5ukIfXqxOghJqGlyt65WTpBdHj1sq/MjB+mCix8H
vngAi/GkkxcQrTRjM9Xh6T1nmH0qJ+QhmPceIHNALnaIM9TcDfz6MEEtrN1p6GZH1RNfgAjibGjr
NcU6BO9qSbsvnIfiYlf70PS9tNMQNntHjvmuUySQfu8p82DFxjZCb8sO9EUy3h8WGDNb+uQaHioc
d9YJyPbIZIrBrL5sjX7SLJ64IiVg2Pc7hLswidsqxw1CmVzQlTGIO5/bA4EuQmXGBEDcJXDxkLbA
4rCMn2+G6pTqITu5TXrhvFuISxBZOPgh8FqTc37+hNjVoTIZF3cld8abTiAflAsCkpJjZ0xFPtN/
/p/93PwPxbPGtPDfWfMhY206xt6zOdqK4qqMTKeBlrXMIagqpx+gDYPSmnwPUnapkot1fSVGUEVX
MkIxpk5sP5DtQARnEipDdO7FZ84vm9PqsJT0vS6+jFE727abAGZH8eBxsJCWr0FYTlkwnwSe1mdz
kcidTd9KsDm+OfZqX0BZE02sDZPhFcu7AwDzrVWQalfIPz3BLo9NOBYoTtt7tMynZ7kz+d3dyXTa
yd4WgYx/w91D5RlzrSsJo+K6UFvputbdvVq3f0qYJDo0B1vav+mFj/3yS/tJaH58wlV54yqsfegI
T4LKr0SQEXvekjtEY1Cu6mobdQ4AIlJ2/rpfOneCMz8AySuWN0bHlHPOtN6lfX167GYF+acNu/0H
/RwHPTRBzVVcmpaFsVi4hru5foF31lINDNv7LcNibbOtPrV0C3e6Q79vWTJUXP5sX7hJTOyyfuwA
RLYYxOiknMBsQYP/JGm52hJcSR6OxpI4FtgtzS2AoPi9S+tBW5Wic7ckl1O7dmcbSWOiyXzyy/UU
JsIh6gdiM0n8kNHRMSCXU4iv/TEGw4Zd16YVMEZZa1q5+eguLa3hITX6B0UyAJRChOZ5TLI+UbVv
1Iw/UBhfdGWr5FIhyNOXP/Oj82BUy5Bixnqzmj8ovR8vd/kKvvRkoqeIkkuCuSVvMILkrZvenVmK
wHZAT9Q0Wd5uy9U1axVAhxKjNBSfET6/39pY0WWsdYEao7TWfOKoWrhIvxLyw9YYCSEZiHhvN7Je
7i7eNwKK5ftqoKz9pkC1JEinU0xLmdIAgMloWDDuvb7q4Q7/BRphEECOKxDpP5fbSoUEfvuakejN
QGh56XFxx4KI828Dl1RrEI5x8HQZC7+jBB8meYfyzOh8aCIXLkb7vLd2TG9hEm+D1I4t0A9B5QfV
akaqFX+qNfjWLq5POx6iFJhe8W8exR52wIV+a63V3jRVd+HsyXg0kjQVyhmwv3YmWYyKLITnThgT
hYVFpF84ZjJKKh+RDvek0v/YJNDxbvQrg8fRvviDHcZkTXbCnQDu9X+jWH2NCK5SFQDMW6Ko8bfN
K4Ex8PR5i4L/HcIw5Xy+U5Nuv7PRvBomAjlRxEawkQ51SmjP92OholgjcH0eNRHQYBPObs09b8lw
1fUST1JTfK7qQ+M4nBzL1o7UVJa8uOjIZxLymlsX+Aq4WtIHyH2oH8svRQEANoEi8HhE/6AmXQ/d
35sDLJmBMjNmWQY85tayUBQiWq1z5yvK1cgxcEBObp2x14W9xamK15sTbFGaXDj+8vIBWrRWVl1S
FfSm6P6QUVZtXj+KphtWxVRgBHrQGWnx8kclBcJupCUtrwy0znP+ynPBKLpIbRc0UJyHaUEL+vqH
CFDCSAStgk54++0RNGh8fN2ra+ciQhRTuanYQQYIMxQPogNz9eKlGzZ50BGROL2eX5qRCyUXM1gM
A1uG12QAilcSY1MktkkZ2E6cOAiZK/NZGqDxTS6utZS3itMv6pNQSNUj5JAHCK8/1ftfJ5G5c2D1
4LSaQ4kiK8rGoue+oca2+Rr7Z2dYWO3wnVGIDPAFtLjNtumCEExgK2i4PCfU/IAMxUjSL6ddygvy
YVl6f/bB1+sBx/5ott1aQYv/0d7n2CipaLs6HjjVvDxGh1//dlMpZ2zgX+P7+vmWgALdcyNm2Wny
GeSvvPk725BEn1U9J7C4BGSRPEZH8w5mzP/1taepJHlcSAEoGqX7s0SpscVYsWMCMLXMOSl1QFga
cIFXidlSv/U4ZpiG2NKQ0g7FPrbqipzfacsZybyQsX0PlW8SyBnsbCvvAHmDmXtay6hYB6GnSRKV
G153Dq0Qf77xWwchH1UvvKhhQRUEDI0CeP9Pzs8pGHhBOHvGbhA3bm98M6rGYLXS8WJtQq1wTaq8
E5dL+klCtrNTo3GcVcpy9XkXBXI1y3Kj+KxhjG0yI6BHOdHhMCDjoV5mJ3W3mH+QuF04U69m9/tC
DE1mEdvg7qjX62t4++51fjMtPRfOgf1kf9VUJ6e1SqINwcXd/K+A3BB/Eb31qXP/nq1IGnX1ztVp
iPCv6iTJoyXFg1Cbos2VjbdS1HUi/ro76CP6PrKivbMRmkFLG4w7eOe02Jy8yBSpC9Nq4SgMpG0v
OF9AvW9zoTQUrQbXAp9w6M7kxPOtFEIMGsgwCt/ETf5odLLIoqKaqqT0Vdsrd50DK4HSWM+oKKLH
8i0t7H9Uf+YRectjga+RYp5RG2+H0/R5a9vtQn/O1HhaSYvGYHXqW5rYXGNkbJBUP95GkwU0ZG5M
Iw5w9hgyBqEYoQvmkeFaX9sEN1uyzq0wcQ2WXAGwZPnZtxvnpmNWncXd99BaAo93DR5OHOmCynJI
FgvX12ibws+I1NRPpPxuTnvfd4IgaXXq0uCMUnV+mmLKEG3guZCSpGF8/pSSkP/KAa7NWfbYxQ0w
xL/qeQNjT5+ONqOcajSyDOfT+8+NYYRlVqE3NQhvwCzyHc9ps/W0X2sYxPt8fCX8oyi/9la9ihWx
WRtpTpV8nkFYJ3a4wh8f3ekRY6J8qTGF9lfrZ55gCAGBVto08VOjzouYgfUVXD+toJXrvk8r7TNA
5WAF3rsypaAmRB9wqHHE4UtlUYJOJPjLvMLJ6bm/Wpsa7ZIRlqW0TL0++cw+UVUK4HaA42iBsPBd
qgAA6ZehJzAlu2AkxDjg+9U6NAxhG/dj/OuDxQIHVNrd3a4yYr0r2b9FJrM0m+QhSUhebmKYfCAT
MUb3SbDA48gDtleJcMlwrMx8td9m9PqSnDkySoMhdbaXCbeKweVKRV/QVJBMd1EN/TaSdfL9c3IC
MXULSWj9/ODQwUSqI+K9KvC2HgBShmx+stE1Ez2O2Ed5BAKMK/Cg+rZj+GsVNy8y+1JqqF2MSG2K
Fh1VhiiDIUADSXowF1/VCxXPM2qc0E1wus8dO9jzWQAfoczOYR64w/S0aZYiNoJj6TbFLXAnrtsc
NeM0bpmjzKPSogcHpjO2ZNpLZBdt5Sxar69AANVn+vwP/u3Rak3Bxy+MVUxXXS4+qkpZUVD5tbpe
pW3WATYB8rQKgGsI4FI9TYPk+Z33rHj86LQ6Iq478KnpdhUSen33HyXC5lT/fHLbwcJ7mKHwj2PJ
YKapohohL5sfAHmKHwcGQBDgbTvs0gPevBsvb+fQnfCAM0X1dMIaJo98IWhByKjtBvuVhqPjshg5
md3t3U9Fc6KiUrkuy0q9PcfXxTC4ni5D7z5opLkmiXRH1xi8T3XZn2fhnnX3f7tJOAtJt3uNT81J
cxWThTKtiVnrYfAeCyJ6NTMKk6deXRqZxzgwwasP34i/Bl3GEXSm5S8V9ymDAIDCZBkhj5XXgprK
PP+NiK0pam05cil21RCIjalMnQXAh56xGrHLfa0QQyszlQq3GaA2u5Dc+0iOp7lEEo6kAP1/eddw
uvtmBjQ0Bn1mWBVP3NK0FQ/ud1LKy25I4poAVlwPxO8aGYd22QMOauuokP9gEDhRDwV5RTt8WJHC
8CahHFzC7Xn16qzs63+iSHh5RDXGxzGagE3nrh7ThqGaK5bLqCruHQhnxz1lheePwfJanVlbQ8F6
MRJ0Y+95xBrhrDNQSgLPmKgVdb+aum/zJGHnG2xdmYrw1lFrqN9ysAg5hPr61VG8JWiSZ4EUEpv/
Fm998UlZXW2Dy1es46w7ocok35xjyV/hZw8Seqcy+tONSGRcDivsF7oSAf/LCLaJkzxIhJJ42ASD
AetMo6wPt1/Tqs/OgSKMYHA/hDHrGSEzL+NhmgPObmknQpFrnbn/Vc6voF0Fas2JOrthST4clSxk
iow0YtmP+6jpfNRawsIiAebNKp8ACOiYdTAdI7Zx/A7cMGHUTtEogMeHxulDLUErIO2oED1SUD7G
91sZN+i4d8P9sisCe0N7EvY52z0o9PZVu21Leg5Bh0jrOGlZrjBvLQTtVYSFPXd+vsxS01T6Pkc5
rpfFK8vV1HJFCymM2bQUiZCGEjUgtXlCVQerS0fiGU17CwbcegcMd7tvcUcoPmeG5+rz7RkEup+g
OqvK3IIYUaRAUpOywf12zwGNtJuLOGjCigw8kLpugkLITUPfOma/TRSxjDTGgmn1wchqu4woX0SJ
MgeaVlKULJA1JAjKAW3ayXi4yda8WuZvJWXQPJpZvmZKsmxbLoW7LYgcxcd+2eiY8ZBcW6Ji7tGS
SLVXGg4pGrKn8bJFqatL67G73pC/RixaOB+bHmvnhnZTSV7N8gGODK0ZQNABViZ3EXYE2/OQGrvO
fxGvUpyEN1qSYMz137wolE/jrIMcbeES+R/WP1k81IJ99Lh5VWuHHXLy09BFgl+YkWJR6n+vvWea
T6w2Pq6UA2YthO20yox12+/TGOX4IBo7UEfN2t9zPFYM0jQHvcUFAErUbcdvb9e6IEMQpLH04Ib/
It4sMKhJA+rcdNioq/P35yei2UjfwzgNMLx8zeClEcBFScEgqI6LYIcIM+8pb04j7C+6b79k3+5y
7FZdiL+L5WHJsJCXBMPEpWLMHDBbmRuhdYEGcn/Mh5O96EXRwVLS9WjLrmciPItfJWD4JKnhWF4o
DwR9YnwJrucRhOaMXBhn0GxInPlzC6aF2ElUSnSL/vTQSt9sZ+V1c6FLzmu5CtjufDwSzBK5G/lV
/2aEqHBoK+JHfT+sdAJoHKZM7wkHV5hTYweXx0B1U5IgBzEYp1PxxBJ/uWqOljlEZ+2Hyoqegheu
3qkel917ScWuXA5Nug+Wae678dwy/rspuUZGChcZeUXi8VJHIrpRyc3jZx//OskfC+utfIHXPP5A
McSMQ5myNtmHgJdd36O1e/MhL0cPInb45lzq4qpvPqHq27rxDT3EQ2737EIc31/aCX8z84E9O6VR
mXuZGxMJ2Do1dflzC3M/L+1zVf1MoTa0RklN+jTS/+0milE9YstkdcxQ0RrameeYVCzWeIRO+TZA
xhPwg6P8KpbDvakDG5DYHuKtw+Q9m5gxmG00x58YZ0dAuHc5Z/MZXeB4ZeI3FDFz2kg6raZJQwoD
tGZxISpC+PpFYqUS+5wa0OseDzj/hNYcJhKMZVWMCVX/JGr/24SFxGHxF9ub5dYuH4lpCJk0bM0t
OvcYzHKRqN4OOpulniZBQEM7gbeI3Z4H27ek+GUS4gPCkVOLX+laj12sC4z8tFCN54WQdIhwwRpO
toh9aiYIktQQEFyz5OqoDp7y/kSAwqYIVX1ZDwwGG5VEF/8z2pPwtQ5CC4o3iIgZyPuI2YJcO7E4
CVUTK8qZFxVhvkIstomJAFWd9fkn9EDUM3ijPlit5J/NZYNpqJtb0aRVR+GrZ9lrBJrIon8wvAef
suRTLFi6EXhoxReuL/OLZ3bhyNp0jWOzmOSEDRwi87XY/VgswuF9iV1SfArVg7m9Tss/KFnKBDU2
FY7M1L55aqpBnb4QqJKwnKuT3TxFZijmPmGejzU8bEoyQleZP+T3h50EU1ZsQeTwUMc/8INU5gqx
vBFZIDrM/85osn87n+YMDLezBZs4ETUM+4FChxbNz5yOWD8q56SIrRTllC84QOnxcaKmwU3sfKpS
GgZ3Le0yVjZaB4wINbaA/9VswXewDRj4QVqc682cYF6Z7O+CUI/trPYndgRZu9cyjw8eEMSJoa7S
MCMbE5087ki+hYgxaGjfk6lrs79IyZsN83nQSI84halF9Rs3tsuK3Z6J2u3aADUskXfEMDt7inAe
oMPRpjqy5YnnBwYRn5fxWczP9o3RKVEEncnr7Ib50bhUK4MDBzKW/UflzhrCWGuCZ0xfYeaGo8Ec
QsMD3TXaNYGlXcafbLNciYU80RppbgERrlz1khla3FuB1xFopeiZqtZyJxGKHAvjfR6x8dQTGIch
obv3avpblYUc4ZTowetJCO1exQxON7bN2nn0ongTULD4we2XGt5Dbu2J88b6dT26dIgpa3y4aHbQ
RHEZlLbYr8cbshwHpuNQFPYy4A+5qDCQifCUDf5HerqrYzOMTinT4OtN4+2OzYKLFCGXSDF1CAFf
QWGn7I1ZGgHQmWWPPRfuM3SHYidqejIEaIVp3rgfnwL7/PvpF95n7KoLkhWmOHkaeRSpYJxDcncC
8IBCi2Jqeq0Ygfa6asTSL8Q8qljqRzy7RWQOz6cYK0ffsgvtUe19vveq8ksDNQxMZ2atc0NLlF1X
TKQcNX/VgU5vAhr3ORocQYJqLsRSVB1hRXQ86T28fFG+grRCEeth6FNPe3FpUb4h4XbPcj0HKERL
XNt+n6j3PnOjh8vFUWr2Y/XIfnSLMBp6momi2oZX7TcwzCa2Q5QwEziWtcV6cYG4t2fyuxF/k/tw
xAZSJd82YZ063uIw62sBada68xj7Nal5wcP//hjqMLEn8HFBh1mFO7wBUqm2E/d/avC96CH+botz
BjaCFWC9t3Y1FRA/olEQiBpv2NPu72lk12u4uJgbZ/2RWUzU9Az2cpw+kPScd5YXqzQtYxcittH9
f8Cqrku6MQoBajvCsoFTUmGhs709CVP0djYjASzh0MQkm1V3goIdPAUd2zH9I+hGPBBfqEFnkOd0
QODP+YBc/co/kSOJ+NQXkFAHimbgLwJXeBnY+J/TRx88ZbIX5PGR2lzG2Ns/c74Axunpz18yBHSX
oDKokFGPvA3IqK8HzTEa46h9LO2yx1mkX/UKq67BOrV39DbQR/yZvzmvXco+818Z8Am+1cA2H5Gs
vyz8F1QmXsyPeVrwODkYYbLunfDFFBEMrPpsGRihkbXzHlfplnGSyNXBx/nhUEFC5qYiFx4gkGQk
ZAcfVC5nJI/zexnvOLiGEkhrUlZPiXn91Wn4l3u1SCNgfQAwAyuiHSfmMiq1GL4vRXtrKN8rtxHm
Dn6XCP2j6MJ14EJqeCnvJ3Pef4khXG0b2v9CgKhIbpS3cpKQalPoHJ2GXdH7flC12L8lRJO9Sgck
KR1oNsKE1Eo39+0MaHVQ+NWhpDeezJz7URFMnkvxN7KraJkl6OLShRGwf50nYfRtjZHXcQkDSwsK
HxLGabO20MQAaxV/tkeb+m2n16C9PLLkKXngcdETKOTFQVJCkf+f81pxxKwkbida90S5ozdGh7rs
VDEc9ErtAxCer22jNhI36DJ9Adp4R79V+lWIEUJGe6ZSmhIWla5/I7Ld5dM6S+oMsKU40t9CNwiL
ChioXcG36mJw57U0AFZiKQNrDvlYVZqp4JpfuM9cSbqpEf5aPvK9zZyV5a/8cTMbh11gHsgH6Zyv
gtQKArG9psqEFB7F3Dt8T8LmRAV0zSGAdYQJhlx1IqwuMEFjL5MwZxVvsx93hPNc3Jt988TK2Coy
/7gM2S1lJsh9DiJgbGPD1EQHkPEKG25olJ+6Fmd9ztsWHSNr3QwSqGiuSxIncFeJxQruOKz3JU54
0KoDmYS2gnc//NNFx3zD8IXxiqJZ5deYDuk3p4xQ4rE8bxcapD9+zeLwZ4K/VbLuOWzn6Sj8t2kZ
umE2LqFQkn6Kpj4/waFhcy6uBqvnnTKudrtQSNpW2eA4o1nlQv/1YCMdB+rmsrwogpG32++3w92z
sR1t08t/LnQSjWKEUKvh6NMCB+w+wtzEVPPMQh9FQ0BQ2kkkaECCJo/pQ5aoBy+iAiPkEl6QEmFt
s+PtLivPKNvvyybI+k6uW8VpeMuLlqfJCMNM0c/yZXfRZ5SkSPaxG5w4SeihRM91S8gY0hkxrzNx
Bkt4ZO1h5TRftYwGvutC5U7T3TUHQKAAFEdzTJoJMULf2PMscD1N9YgAVUSGsfX8fo1r4tDIxuT1
DmuWNGJCOaWzxKysyQcdZAbmL83IAI1x4StehDXItNHwsy/o7CDjnZ9guP/fww05Xf5XY2nAcGS6
w6pwbJynVMJh7TguRJeHtw4X/vJDzc9lXcJqKjoVdwxWoaD+SLRQOimzAYOdwDZBkX//Xqe/Lql9
KXDHcmElG8ZfTqvmUTsglMoHM7hOevmRYg+0Wb6SCCWVCPvShtEqRC35A6nBLqSm34zSTjb/u7gv
PwmlsTcqdImTwzwH40GpAaT7cSrUCvcPb1VwFUE3lvPqM5tIKuM567Ax6V9KJraW9Gi1vuc3gvCo
XdKF8KMe76XrCW/UNnO6ONE2CS27gxmzMZf2p6lyDVSil7v47jU/ZHLyiB1XMh2FnXC4uc+wsltY
Oz60a0jNpOqSgbuSHl47v46CvU8WOmkGUwBHJSJ+P3870f3nqZsBt9lf3ut1NgXzSoijFXQH7S7t
qRSHCHOwe34ibje7B+HvpWI7xguZiAAaVILQzwtE1Sy5M0TDoP56G0UwjvSgOrEk4kkm1XLqbpkr
t6J74iyO6Jz/J92KnYc/gebR1Dlmw+IX5sE+fwICPB7u/GFrliGswYRJDi3LRjH4YAx7aqJgb/1J
THwRPBMXjyrk6qfij3ixeSegtdD5eKmmVAuF4JkNihWfNyA/YJ3P6sxb/bZZv0pWAOy8BqeE7K62
uPhutYWILFWXkbf3/JCAcusS54q/dEfJzMKPxSFsn/95hW3nMFCvM1JYopcc9ZRZizBuXbHDyuM7
s1mF7RSGxCd2fwt9BhOyWOHlCgtZQA9+suhyh4+lhL8IWq5fmnPKobnEgY5wmS5t84N5L6bPYM6j
ndN0FNoxtRtci+OC12/1nndur6UU+J0eQpbjQC0XpkJ8Xl6L7YxjeeoNJUsZ3feUmsFXZSJqvXrV
SqUpYK9oTa+JTJx95GYNFsPWGcvJsn3bYC9lQQyvYJutvnZFuP+XmWFy6/oKI6tiAGGhO+GmoTCG
953+EOzpX8cCNQE7ldgMK9bOvZls0CoB/uB/uK3H/dlcbpaJ6v6yuoUQQgZBUXavZwdPXRs3xaLk
PyTXjx98RQicNJNleOc6xkdYeZcNQURiHL+LhjOrtd6AgdSj+MT41JLnhLWf1kJspZMlwWvunAcd
/aOfRTsQBBGMBhyNox1h3U5rRrKBNPuxDqXhViU8BXp3jfl47avm53Xh1rPKUU8lTcTNe+HAqmtF
z81wp+1RL6vW+itnLLDvEbg4AQFgrPtyfCIipxNVj4H5kzOiIMqBhvwNe6tWI04goLcZX/SJcJ+M
zoEHU5xyr1BivO6t0tcnQSHXwvFOZmtmtb11EEQOJD/IgEOq8RSn2Q6WcprwGKSwiBpxb/3eXD3S
YtRWOXECwg7P+bzVwgSwNZbkjRW+KzAdd8ySNF3ZE5Mia2cRAp/SM6yA3c3iml/q4eIIk7sjYdEs
uxa+2wsDzPJHLMqmA54GOrn06t/GbTmCvuX68+CtVpSTI1mD2yPnuuYqoIvYgbx3tHo9zhDtctBF
QheCVuMLiF4aemyWYLyUOIqB+S8M5qv+DOKd7rwl3QEhsr+rATKIdtr+Ykd1+sl+jWDoSXzMPKb/
gzZv6xUwmRZc9jSrv0BrRy+7cIigX3uQaK5GB6Qps3fz2kXl6sBoqpfzcXj4u05ENxaT28iOAilj
CB/HaeKkEFh9rwYQ5CFpbJuA6m1wnC9Ib+kD5KTop7/kGE1F0+S/tLw/MZr0D3S4geYydE9JWEf3
FZpIo1pLWM14jqfy7KnognQosnNSfupPnRyrrMmabDigvzhVpXjhj8R7IaLywKJ5FJXSWRtY2lmP
TfDsHbR7gUMgbtP8zuHQuN4rklRTd1NUwVYGp5LTynelsT38d/lf3UWGVvvQKkU9N4ZtZ8V/9vKV
6tNXLuG7AI2F8s5D+1CZatG62YQpotccQweUPxZA21UmezI1wt6TUQLiv0DSAHwt/2U3fnoZyQvC
z3P9iAJpBtPk4HRw8ZaUdu1xFyEOO4t6sCZ1T3ii4n21rR+2UIqxi8J8V56WTNjKWGon/TOV/9yW
+rtxm5PtT0brh0qj1c9y2J24m/tLQUVGQrGlXi0fhj2OAagMyTajvgU9jvEIw2doQ0iiXPCztZ5L
gFAHz7WTUZmOcI9xfXEuFQ5G1KBOkWn/fqXGnIJg+haHmXEZwAXaeW6P5Zfv1mImkMU+xVhJQnOy
RZSb9aHaAsrJu13eNX7sjwVFo2Fv2Zqg0krKBvWCJiopRnbsIKLzDhp0WtEZVEoZotJWk6A9YUQd
wazKBCgliiAKaNuzuX48i+tILbW4JhFsUVEBMlXMwecgncxvErmtzs6XqeUSM0zlLJNcnVusC+g/
yckdAgF3aiP1JeDnrtlrbV8u1OQbHlA2rTs5OTnvCbciGom6B3/zPh+AJUKa0T8AbYt05YTEqh4z
tDtyXbMZLCdfHUChvZItRxneMTXnYeEDTgy/Y7szQ0alb4R3dJK4J945GqD52ZkcmU09tlffPGUC
tOgteXVbBdFwsFN/hxxm/42+FnfcvtLK1OJBtxxWiSzSh85djcSC/XZyhyEpHIHyBDLup2iSnc3q
9xriKafrfa+FnRoggwPhMpp7K8jAr1v/6PphdNVImYe3LIeZQXPo4abqblays2L/g7a0TYEIqI5Q
F+7U1cChR2NpS8a8fqEV9BALWbEgXzxtXmKbimiaSec6KEwQ4NKNY2Z17j/9M7VDVgjqE41qNgQp
kbMIzJYVV3iMDBn7v4OK6pwcvXb/AiOpuZqdHKAZylTZ8LSTjcW3mOTHF1tYAlxlmhxbo4Gb4SSc
gMXh0w9UGdCMMV8JnjPGlPPfNDc64RT7vnV4zatHVQFy+fvlMU358YI/6ktiojiSW1FhNlV1oY47
m4BUa4n4i/L9B5YZUPU16FYRp4auTbhAnD2phA0uLyupBa3BFecZTsbYwXog1xHGQcVoKKYQEH7N
8aWme3MAQk47+/do9In750+Q3MTec8qpd7IGKPGAUZaX8nNKcMTn9XmZzBa1+QlzHGAKQwatWWzl
Uqi8SRKrkVzTf2t3uFx6F6YlKgXxdYFxQv5HNGf+52Qos3EUiyCItEJZjr7OOHdymH2Fs37FWoxr
VGG/BzKIUYHacT2oqNJ4/T53u3BmKBOQUaPzAD4pKQ8PF8063nXUcmdAwN/VJ8Z2+1SOhHou9eo0
0oT660VDhHFSQ8WSfA8QU52bFRZucvcx5aYVZUze/d794psJpMr9iThqMy2NF5v00cEzs62qpO7c
kWhQtZGF2x1KbWcdpN/qLG3SsbNrHWae98EpW2wswlESQmqVcXbPiRj6tUyJu0isU7ZXaobXjGp6
ohl5696rqH0gCa9YcA+fNqm3jty6WWuMXy71RbLjvw8b/uhClkWiGYkxkqYAy//MMGKL7wBeizQa
VraiVRwSv99feI1FLMHukA2JsBisRjCoAjduYeaC3gqmCULyaylXROlWl6sVTE53/MVwbl1V764m
U5QfaZGwITuqaVPt0XCVNzu9QKfsd2mF3UizgJWx2MRe0JFH3Nm7x69vix2v3f9w40gfG5tKpeX1
3T8tooRYinpds7sw+ShiMePuGaid2CONFp5lMvLoNB5O6LC/W2y3cyUyPj4KcCLbezHmBXJW7htq
G3xLWj5Ak1hwlpxXtyD7mOkqkToWrzh24ymAUp51ukCfwFPjXYL/+ZGiDJ1/c6QLEZBms04ps1Jo
j0wVIL+Q5/m9bEkwm/u+Juty3DgfNixOx7P4D0DfzDMvXgI3wCFcykV2e75RMU7SogHU5BuXlYbF
dr6Cq4lyqjX2hME15vPhfb0ThgsyDHGSBxH6hyvndc98fFD7BwyDRwtbgTP+Hbojd8jzCufuwy7F
4V/i1OpcIjlFetPJ3rw19w36LL+gqnF/QqrcFDQVhmctjeUIYiyAFiXwuLUPvGac5/27yAKbOzo4
PGN8xxASx85762K3ax9cF7es9byOc+Kx7Xq5xM1JjwG3gyq0I/Cdaseg73eBuDXvx+jKFI5hBazd
sRlmbHx6bliauPMryLVyozdcKx5nIalko85WNp3G0XRQ+XxyRHTeR+XDNTEBEkdzbqig1rso4F9j
G/uB8mczMPWSSxM8+TvWRyJOSYAVh8xixs8OypWrWCE7Ixw+cn2HhMJU5GyFnjATmB3Ul+GiRFGF
NbXQPg5hDJWYwYTrM+oYVmwG3IREZzQs6tU/hBV1IIwXHwu+KP+e3+Uw36F+bLLDTcJv071BVHDV
5n5/X2T2jn+00IWqURjAqatYGPR9lmvTStZR9yCDuPN4/1/p0z/6h+obw4skw1x+Su9UojpSzfl0
3ACc8WLdlu+ZVWoLPH16oswvL+JKZxgi/0Xt/tKdIdjxef7xwY6AfV4Y23F6xpmW4MDpw/aWqeiJ
Cm1EvUJzL3206OVWvsY/Y05LDh+lo5sriPAODFj2vua2yZQi2YdKUDen0YX5udq03qMnPmX9acv2
E+Q3/8+b8J/RGCVJxRNKm4LATwJoeIlwMfRN7GiaSIvK7jUBpmFfWqpDDV8z/I7GRUQ7syqogWky
Ps8c44gtOZL1MftoJcFfH96g8S2zY4PNjYIGapravaZwFoWIBrxRy+eVCIIOC33Bb/U4iOrk83vb
ZRdOUXXKlIuARKCupOe48YnbbBUReu9k6FWz4nVSiZb+ME6rHxx2kAAyeDk2A+kytjFRXkepEqmY
opbUWt6ygYgg9Pe9BKNdhl1BBvBFfhe1Euyra9hr5JHvUgMRFTxdgWLQ92RW0k4D0Hw4meIuRSui
Z+a65xPlUr1TU84kJGJdlFUyUNnIg8wNrh9k6SU6O0b6HceXYNYVZcWgr6HCBs2PMOz8mSu4irIR
rF2Cj483+/vB5T5sQIQf+OFv4Sp4iZbHlnZ+ljtZOGXvcuR3ileHK1AxzA71s0g4NFWFSl4oTMyI
HMEHj+i8667vhiV8jzMwa2Spt4zEkkLbZOgQ2qjv2dnQR22cwgIsCq2SHwPKvcoMs8W37h03QVD+
nTE0z8IorBOjZ2vPnWpSffyIHeW+r/aDKh+aC26xSrHyKfaheVI5G6klamCmzsaSy89kppD/0l9o
jT/BGpWUOoyKqBkCdQypKU4bXreHn79NjnKOBoLZAV4GpR4trLWH6AQuy/MitwEtFV5fl0dx7hgV
QqKstUZpIH5m4hg/ufPFSD4IcejxWDBInUywsojLieyDVCPeXUCFbJktR7t02S/GCWflAkDwQFQ8
isYtBAMKjfGHdLHOlAfI9QiIaOUl5YgwCPH5YBH8gj5AzuX3cOl5Wec9izd4H8Tnf6fVHhwnC4B3
tlsMu1lSo4A6/3OCvVgmg0q71V+41RSv08ejWsmeZyxF21jn1NlU+EBnmYujCcvCyaWqG2wxoeC6
rzyRJlPaz84k9PQbcTIpq+CSS0Z9WW/76r8o/nUzepDWghhO1AmBzV0lGDclYoYDPkQmcYnnIo2w
IpC99ZLe73LAILxO8RhOjeiojIwF6AEQhNlkhwH1vy/Dt4/xFlyt8V4fP1o9WLQHEbLtHIob7q1w
WBgaLZ5eedx74vagMDH9sZhVipUbyT2ZecIbwBTdA9yf8/9PDI59mX+jfsrdo27H1KCSQZJnfEDt
BH6BMiQgJFkoI0Kb/Ld2L2dqqhTJ1Edty1sWIs+MlXdaBcDsrhmvcGEFB5ThZUUkLEIQm4ZC9qyY
hCNaKAiBcWUcij9BOlfDmiy9/fc6+CSnLJibJYG3Ac9ZKC8xtm1+nRiuWTd6+qYXov8P7yr3qkSb
R5ArALDhPm2d3Fqn3axmUp6awCMARIOLCf0biKh7odAjktJOsWVEcr3RfllFhki54NnaY2s4F6PA
Jaivr+P7DuFuCY2Fnep3ClcG1EsRuPEu0zMjui+wcllPVfQ+VVlLCUgPjmv1VaCLOqM0uswYJ0vz
kr7EFbGuQhHUoIEZVUUaufFFudWZLECv8pBVPGVx2ceFP0VXVtd+fYgUqKNJ+E7uRZ2ZV5KsGui2
pRxdOqU2SGe9M7Y1p+RGa6grmOlyeFUhbodIttnM8Gc2nF3s7Wns6RLdYfX3HpDzNQzTA6Gt9XP4
uFILbw0oaXpBCR956IBJRY77UFMpJg+sPHVC3B0n7SIgUTq3KNbcr00UCa+wvN6Et6jhIapaquee
RCamNRFd+8Y+o+mK4fpZGRyqejgm+5Dz5GTYyyaUAcOHbTXbKk78qorLcu77gqj6hPLtYgG/Mvg0
05I4rbaTl7pwQUdijwSMsKhLSoUAbtGDgH4hdiq9s2CplgpoeY83Oq6CfKMD03rnBRSAMzWyP2ls
EHF+Rx6+Fnh12Lpl1XW6D85BYJ3jCETvM8RP0zi5SDP41f1nnj7lmsHjoAalZzTXhZgPnB8jT060
EaDIC3A7VvrcdzqkSSEnb+yNsey8FlqJaIN+7Kf8YGcne9j7l6rKC59AXI2yEaEVihVdYSAeTL0c
09JPJUy7wbSehLvb9i/nC2iKya35q6s4oaRLXkgE6XKLHZvso3VMjmxAlW4eARjqN6Npr8fIHMqr
LOnL1qhTAv4J2uL2FAfMeY+uStag4HnwApZXm2jprHTt8Qcglw3VLo9o3Fp8+5GmWZKrghDUIErC
QcgChY6a9/q1wLaj4rrZykHfiYZAoQS9KLGdzsZC70CZSgOb6/nac9v04e3pCY6BEkrYQPAHvq5w
E+wnihJg4qhH/iD2i7gfc3VgN5fFPMsMS9BH5eAzB2NwTxFJoGOn7YV05iEo8NWGBo3cFRAZlTj7
YlVsZojCbrKFFzQIUMBXqtsxBOOIAarDkbpYfCzKOaTwULaBSe1nD3524BWCl5l1UTiRyxqQArAo
ewnvZK0kdwTWbKgmFl6SWr4uw84zOGPhXTaTFfmKdDUfFrizApfFDb11Cwx78R29bUWIrdvtATG4
r1CqDiNznbxJVWmjgnFp762ucXA3AAcQgMTVSE/Zr9BpDw6NP/JQkMGdmmF5EicUnawP0RaBCugw
JuCvwTaxmMkoXgyvft1FcdB1153XscllLEIdUwU89kka0Gds99/X0RrTV047mltEa6Npd3Wr1sXo
ocrWKMAAG5939ekPjZoYb07ze+h2DsaolSGUlEF209RYSInW/OWVYMtqZMv6mL+g9QdWGX/10VGb
3twk4+CfuLsjw1OQMN1Ap1dNFfvIbPOhNnLR7eo8iV3XHE+CNsnnG1wqhVqOqwDA9PpOjON3/Gz3
3MDt0H1KhX+UO0Qh3UuOFvKiVSoVSKbT83QF9/4//6iw7G/IgqGUt+jiSytXdMh1b/dmPt1PvPNA
DXfyvDwjJajQIPg/+T7yqNqbPQuZZ4Cg1nzhYttSHjZ8yKC8mlb3nAFtEW82RjETaH5fv1u+TUfk
BJ98kg3OatAu+FB5D0dYmx8durSK4J2bHXm3pJajI4AswlWxHKz9osGKd+ih/8utDoBtEux+NBCe
4NXoE1juChugYUEhQgcRZ+lnKyXVgKlEN1ZzHzIVmAaG7cvAifsWA499mzi7VmH3XPpj+2JyYoXZ
V/kOls4cvWUO8lgDi1fRnSN0gVOTw9vvedqWd21ckGWbWtJE4u0JYbV+Ib8QxAdyurHNWRMw4Su2
4oDVAr3DJRWjZ/QZ4vjA1UxEM5+4M+y7/cQA6W3XLoXsXHGfcQyE7iFbnHMvGHHWnM+xrqwec0C3
5QvohlE9WU9VVjIPs42+tZnp0U+C/DUZQ90skeDaorTaxrQDGgeBTIIoAzTE+0fkJUPOtFvRlwSA
/wvMdw3fgtEBPwpkbT2rnOyJXnsPaujGXAQ+18S1eJvffuEU3OJZMv0VLI4rZ26KEpmecf5axyVo
kK73ZxN4oWGKkCHUkSEW1pNovMAYoGACeAGQWFRpKxfPa4HDMHj+2NzSGTqSQOtPyTOR1UgW2/dF
MWmW7r3W7iCyoG3fL7SzqincJlcaeXNFz1hy9bFljqWNtkmTVZqZBemnKWm4voNvYg74RKimYAwv
wyZCJ9GnogF7dSgDT/OSe3V/cB9jxmum0SeRegavB65uH9Uht2NDYSmQpgQ2kXITQ4rPFZoFq+Ss
haUGnGaS9rXwy7L+2KD3Qlim6WQtiNNCibhKQnyCnX2ZLiPppv9MYW8mAzphz+vMiwkq7rtLNa9h
ubHUEJCapZnoubEaLdRjicy0UAq596N9XM/NwDFQ5tLh0BeTNrVija1wEiuFSCXhAtm0MYPcgsQu
kEXqLlkymJpy1jAPUh1lMpKjrF2VPeWkYwV/we5ez5oIjZFxgED/YxCgNJcLPkFIfx8RgtiZYU/j
b2Tr5C5qlzyriciJX/g4LW65u+PU1Xw7pQ/DZnDliAgm2/2LdxVk8zPuN4Rg6USVVRlPgsfElaok
/Ddb5CZg4NL2Z/DazVHM4+FZ842Z4KKNfLK2qO+wiodXkAGxF048XWqhiLVnJNwMzftEtH9kLo5K
7wR0H0AID+uvm7Y3yxIVw7/1Zr6dOUXG/wFJDRefTVCOFfxIvBPH4oxV9CWloZA5s9xUBBVn0+yV
B4E2VCgxpXfhNh45HJdhp/9QiPSuVe8mw/gGx23LSRkPZEB5ymrwX11wZBarnyReJb8M/FLSnrZA
EAvSVA3iWeD9IYAy81e/WFkJceQQxkQs8U7lctM38OLzC+O86RKEg7LOEhmEHpx5zxnfh+w24qZQ
/pmjYGSejE04jVi+r6FjMIKfX7OxGb5tj/En8MTzb09IeYDFJvOo0CBR0ZdSOpTejOkVgqP8ciTs
GSOCJcKOueb+Ebw67WVVlb/DE2CCdlGcqzjmxeCwD7K35dW2jvt2lXIgE2YYMfkQuJfYM2YDd/7y
zXKJZ0Lk3hyMpaQ86cJ1TobWyNV/E2X2n1TzRImrVy1I2fGOpumjNEHU9/g5ynY+7uNexs2wQ7oD
n1IRr55IC/IewzAsEcvb6otKbfBgJpQxfnbBMID8qOXYkWegPseZc4hiIvrqVUX4bSACjX9u2bZB
f7dWEF9pmPXKCyQ4EbteNJ4qGYvhJXWK5F6rMFfTloCuStWtvW4SX3xHscW9G394O7NiTUpcYXYT
/LLbctZ0f7fbLqr8woftxwI9aiBJPTDQcuLlqyjEI//9xARuwxM6iTY9u1/dkHPNk0CtENFgFq1K
3hvpXnGqSxQUGMkyelTxfB5DmgupDASerKV59a+qjszqBy6npQVsdDBk4G+Yk/9nzKcw/TN2hsgZ
oPWnk65oW1EHSIjlFpqYvZkZPI7KnxVdgbLRdm04U2gVz9PwevdAl8RvGNJPYGcp+TgkSPItB/cB
LsmW0N1FO1DvBBlmSTNNw89ZkEX//9MTbiSTMHdluZlyKbix2TthKtqciKuFRZti+4KJ6PnMv/ha
LP5OihjNDc49iijPgRmqzp46Uqc4wiM+xHjMxENvnfwx0I9s+wwL1DFnsA4fBASRGoWTa2ByyZXG
9AKb7uJLKtHrAFEkOXgfu4ZYwWOuf5uNeEpjFBnXohJl8oCyClbiImJdDsrSr4nHbXhIwDND9dBK
VaVAHFmbj7cDYw8BreSWQXL0vM9mtmgHSVr7pihkjQlIyvRDcQhNLm3JABKNYiaM4m/y1NRhi7XZ
CmowfZ7s8jfdkST5KJhjFD4PnuDrfbF6ta5WW76544CqfwKlN+iWmotz9NC0P4u8mVah4lBkdBUz
Agpz2eSynWGGjQXWyS+U6m86zwSnj81hYHmd+1KWzzN44yN+gHCY6zfhz0RvLAVXxr57VRIkl6/8
eOQ1WZIHKP8otofBRUjnKmFgJDwAe4Mq8jcCjPpSO1orwnET797tfWIzxGSi6lgSSLIEXdkVGWs3
Nd/9xITGXPwgLlGjMsBB+ahPw+ubLz34ziBxTAPDFbrmaTG260gzqaBcFCd9AFHeEp8je3d4EHwY
T/D53+v/QsdYO7AN3dp41UDxj48SmVi1RiR7O8xNwsxhpuOoiMPJt0KFS2O99IDP+NYqTyfvEqbe
NThdIN+T2QI/34rlSABY887IeBspy6BSqxfXZLnSHoy/Sj+urO78Vkq+W17eUY0hwCb5mdqbMCq9
Z+J9gM63+SBNheUJIFG3x1OtwNz2YJRErrwl6yjz8gfjyCBT/URdHgTom3s3Nil5dDmu2+NMfnGt
TaUo5OCMqGqRbNeSV1N0HLeQOFWFzNjOW05iMYutGdBXn9sZ96eo5vu7WlVwr2X+rCpjtLyrhDS0
ul0Og/rwh+jafH5CAFV+n/woUdHdnFJaq8rk/nrCRFJgb4m7M6CxBJa3M99yWMY9PFMsBdx05pA7
O1D6Z/gJPOWwilWohRpX0ZPbZ81MHB4DqKtnv/D/FHOasZIqsqPNzCbCs2p4dV4By9eaagiEsmNB
ZGiSHxBFT8Jm511E9Yr86tK/bT6j5VkBvR4PC7SFNUblnOyXiE3NbmLJkt/eud8sFgwJopsQtEXz
WE+7sHW6Pmc/rIeqdCKd7Sktwa6LV0+prffx9LuP5MN6oumIYG86hdB/l6naXETfNTiI3klTLKJE
p5KUva+MyIhBuR6y5wy2Y3/2BkEef+r0fG/VFswHNtqFKXckexUEBIb5iMgBTEgDLPEQq8us3B7N
cwz5f6G/0xb9dq8Aa/ABAdqL0hbR2FBd4G0e8spsCgTVMzDK6QJjHXb3w3GWH97XNDC8KftLqNpU
rgMACcMCkCVM10CNzfwF2MHbF3iAxS71t80i9I0ySNJ/WhsWjRmo0EwAq54i6FWqJ2wmsC21XJ1z
HppNjfttSQQbnAiJg+rHDaWB3Gh810Y+IVEs3G+eAYHRGzh5wrdQmH+M7ivVM5D09XL/6pWnqxnq
9IgDTRjYmia7w8C0qtD5bbLq/3R+Q/U46Q2pY7ouOiXKNjwTN3p7LZMDXpmZskrhSpv9NcPbuYyB
vQPHw/wziy9ZiYrk8mH6XdAkKx80k5Z4MTv8CfemAj8q/YGdMGftKOjsQ0WVhUbi76InXoMH4rSh
HY7QyqAfNqWakrqkM8acELEuFCMHZC4z00ppkLKC6gX6X10Ul0m5bISPEh3D95b3lZ8JxKOvDc3s
vY3qeLgKCVUgrox+aX5pWZXmsbKNWmcMzGCQCsDvy/2FthaAXBTnbPjIwJKWZnJ5bmhIfKcQem1E
m31HGcEWP2fVLKDPOIn6HqXAPErWKlCp3g/08ggR6QwYLozJQo2LhWiojvg+H5DluIyqI9qHcld+
FUBP+qOaOZ0khmKCR0wbewTra7ioTAl1zmZI17qZe/05AJ42GbGCCJIjuSePoWUIHSMQRESH2ibi
kOkfic2vhFnVrqIajxKhOii9qa8GVL8Qeg/1UBxYw9kQdNqTmYC26gtzrIf7in6PpFWZP1weWYq+
d/KJ858lZtSGkATqh/dNYKOPbUygXKAar6WwYLiCcec5ZuanJK9iMyR1/cL5RdRsES3ylsNVNw9R
WHuimR/fC57yEXjnX7Xw2Jdp2uTFSrmBzV9jAH695Gsym5io/ADt6U/iNYmH1serwpV3pVyZ1HLI
Um5le3LhzGyhb9J6JoaFFARETb0qesPkYjKFs8uAWGu7nhq/vGnnZrLyTUrCE139a84PHzuefRQ2
NTesf7qHcJbUJD09FnZSQSH7jG/u2cMsN1zdIvAhPZKYbVsaaSG/C/L0WVHqOT5RryMILQJjozLN
Db6/wLkAvtPlM45zdgMLd8QEcdteYbOOn1lOzd24Vh0elDNf4KA/NK/ztngYsVhEVFYI+W9bcR6k
bdOp6C9Re3Nt1k1hsCTAkTn+9qWDm/QEjCte2v1jf6clDGF2h/smoN81K3QXdNY1+iqKpM7ucDNZ
w9X0dq70Vx/e5nffRLbMtHEGyaXMvsHwKM9PzDuwL3beqaMoFCp0jhuvN4scnlKa1Xvs9CnO72Zp
BZW+WH/Wjs+zxgwLgQGtehTfasoGAMANWO6prIw2f2D42U/qhMGhJ44fR0nGKv21C61vVY3C4xHz
8S0rP58FB0499TdIgk+hPOp8q5jtszp8mrOqDoV4jlzkyB/VeSALZr+Ze39AGmQcdgWNOqWJ8e8Z
YNPdDSqfOqg7asf3yLrwz8Jo+tj9hsLYnsZFQjgW7FLU63C0IuzNbEZe7sWWZZcSZwjwUv43yuaL
4IAv0QML5okkoioLC5xAyjy/2FY1/+J0ztjgxqM4Er+PBE7VZy9hL/euvQsC/vuXa0zbErUiIAiF
xhekjzk7xwQnv7P0KRWoyY0rWD7G1LhU9UcG7921Swy2fK8ywfXeJzeUxdocE4xmOGFc3ZWS9Xce
Lx87Tztm9riybxNjsCEw661COldqsqZrUDNGlJCEAWTkCjxxJKasOf2piBTV+XxjCG0mDgal42Av
hUIVh7fU+4dMoLz2yfZmjvwCZGOj2K/T1YLMY+C43SKeGVDroAwedYTzj9OEcePrdkCoeTLZWHSL
MqDY/M6BMmzXcvfAMSayc2zO352Q5ALF6c75K2p5ORelae0cintGEibgA8/6HfHZpHmviaCcAICh
k+/YUwVcXz9868IxFYMHx1485mphKJmqLpOCX8yIY8hXjgEXTmDbyTxcPxLqtFLyzAlanQXvOrgI
fmlIqUheSVmnool6MTnOdg8ifpeffmUglKGtb3uQT7Ouzw6CSVed/OIoycdT6icSH/owa+0I66GL
XwHAeL8n0oA8h/mbhx/e7iiR4CxcDvZbJxSvfXxxWnxd0Ng1Qln8iZgD9CSFPCoiGkU7oVNSyFSl
amyAPGjRu762I53SYp2oa3HzqSiIUGUk5r1UHdjuc2pCPUrFMSTWFjbl2v70iwERJMu/iy+C0ga6
5ZBWAVzxZSEL93YNv9DHUavgHFtKwoyqUYshcgHLJNGDQ2YZow/OY4/KjyxRa7fQeJFAUAP4B7lJ
lC32N+NFiPZN+S9g5CFkDytDhq3RooVGvhWboIFBagP5fYUgucAN8aEGtMGHI/SvY3QjrPCYBXLl
TKC9Z1T3Y5NgJHWBvK14yWZBe/iiq8qI33GZmbFbSChFQBjzsmwBNJIRZA4uxBT9JlkUROIrGJVl
0BwW7jSlKRhlfFozkLVlg492/xKUbE9Hu710huWlZ0/O2DMn3QED8WO6hZbx44cth7ADqyJdn/1a
3XzOA6MV1rjLDCSshQ3zW/tzQQz4CMg1kdN//f8kg5NNWmbApdOuvnfnPYYH06CgtYutjKgRCk4U
RLqaRRLaERF65ZDXQxRGWWUZfWHwqwyMMc0cebMOf2cUCnuMt4Tq1nr+2F2r9Oybh8KV30++dkbh
KhtO9KG3eYODH8R4OuN8pTtZSJGyK2S6dOjkIU1tr38n8PzkkpPjLJvlzjSlODsk2DInjkkPPxRl
60uQYQldVL1UDso2Jes2gpEGHz+W2XLQnILry0H4j4RKUXR+bGbmhKTogON5e0M1P18VK4GvJ7Xi
Pv+N0V57uDD6q6Lz+v8CKnzCDM+tTM96+SZVF/eaV/NbFV70yixRNof6FFGvQI2IvsSp4EKAawyw
Ue9KpAt/JsA+h3XefBU5cA7FwhvvIxMqJM74iL0c3w+OMhHUfj62D1UNr9XeFlzz/KewCTvxvgVF
LrnCxGoOL9ic/cPDujmSAmKpoqaWl6XHDeUSaJBNYTgh4BPeOdoFNfJtAtKOT6N9jK4GaXB4wPhW
X7luyBkPjO88EzGlIHxnKEHMd+AKXmGe8UmzkMgoYbdlCuXNOI/W+5VlHOirp0UBqzJHOaYqM3k5
ocnLNFML/Xo3h/7eCl3VaeqUxDyfgFlS24q+V7rD+PV8d3wlJRhWvAjDrzbpt578qBzxAdXfIoNW
mxkElCrIPGjp1FcaUyMyrDPsEVCH11zJGrPtSJgedexb9H+A/isFyR2yXqcapn5J2HVCJL6nJ2rn
k47O894o+F+jDBjLuPvYn8cLn35zZwQx3sqzRlkh7sSMsMtP8lNbkYA6313QRUTQs++bdr5ZSkfq
tw7PD0/i2I6mPk+gdkWU2Qxwg/nFnFxZuoaLX3THkUJ5vS2/2zJfQn3ISukaOu60hzoc8mZBv8c5
KyTcqyesyyx8dtThhEPRgXN7eR9zgdHZrxiQX6uofRHD20kJ0vxH20yqhe3IaEZkWwAMC2ELrRfB
1vnMOEhX2P8tfI9TjFWX0axKLa6NadXK6/CNZYIMloomH1qwECL7/Np5xO7iqAYl3h6h0as6rf+K
65SbnfuQrsxeoKxlvMu29HXGZln4cQKB2zKig5zed2stzHWjZ1ETWpLfT7BxffYut71qSix0aydw
rdTKaML/1Cu5rjg1nHKHWpYpGMhz0gvTJDMZiJc+/o2KJTKyyDXtT1oaDRGr5ak3RXnN5d/Sd6oO
7AaMAO4l2cXKXYi9qqEQyCFVu6XLi/H6mN7zNixlkbtGLAVxKB4hiU2Qbw9a0JGl11ZH/jVYONLo
IJE4QXca/tBtSuYcjCIR26EjXeQBT6G92P28HnBt/WlmbIXR8UDjGolHeFwdllCCEHfk8Ue4X4vU
rU4Fm8hCsyUAdnFSfAdAKogZ9FnCUzWLfr2h/RflfA3Ggixu9MVQIp0MaKVdVQNkYjlZlMkYX6J5
5T0Vx72oPPd0/JxU9FHRIxjPSmEF4IN108eI+DsehQr2VpT5esremcl4G0QIJswsDZc8LOdXoG60
AAps1rb7Jfs9vkKn2AAWd8ltcmlxK/ZSuVN0NvpTHCRy/OLM/i4pJQYmGXEx+42X/zHsqYVIP3Lr
h1twGEeVI/m0U/i2Rgme67EvdZ/bXNnQ2tBscq4WB/EKnuL44RMw2i/i+h9H95U3OCfvok6k5U8a
03899//ul+lVMDoyBrKQ9pCtZ3ifNO+lfBFJQ3gwJsR1HIUerSe4+L4ce5uculhXEU1HrY/NTQgT
9bdUcNnPAOrsHTd2jUXnNxSFxTe8ky8cihpxz5G0KtRkQtgYmnM9QA91TK9T3NdmCirO+Il1sx9m
JohpIDDq//V5/ZvI237SkIoGHks/Ck0qk3Q571rm7hxDWy6b979KKbj/kXsxRsOs1zZmU2zL0L5e
PujGIyAl3u6EmofaCD26Ey3biDMGOJWiD8JwFk0TZv+0jA8yQ6tS6qeofoLY5jPW79rdwvD6H2K7
3JWI6biGmN0P4w7BX0hotvEMSXLh6JR9ZDwnTvJzMqNVXuhJMsSkEY9Qhimyq1yOKQjgTGLlgLbp
Mvmr86nnGCfeeGiJVgUALdnX5u5CcviC9oFapwZxEM3TJBYMNKAmLALBsSlAOuSSa14WrfoPchN5
2zEtM4wcShY/sCWxVyf5rPGkQMtYpEIEqfs+qQM7nzjyr1Qv30p3LkUrA/XyB6T1hyRjj8J6KhWA
1Nzh8HiyKo9IStnN6prBWyE/yne/E4l7T1HYUn+ZTPH6GlilFZUcHzlHCdynEkL1cPdAuRk+RYNi
6sq3n10aJTU4CXiYSi6sA5ocwMBvEYPx1RIXTuZGRraFiTLQ4QuJZyGXfONyx2E2P5fcZn7LLMpc
MLVnjoVO4eIb30yQRp1cVt7BP8pU29N6uo4mCxWwQkP9Zgb6qbDzfcO3pT4DTEYfNdQbKOJvtHqV
NUuWR5i4FGCu1Z8ltTbxSeBdbw6WKKtAX4ozYKeK6r+C+efig8KYWu7CuNXDceRKhbAZoU9+GP9e
NqtanZ0f70TquqSk5uK90Z+KV+MwnddvrH3jIAHr/52H0Gtwk8Njb3IKgL5qmnM1r88IVZyPIw2/
Lqmg5vmh4uyh9JZBgZ0MOqSu4WcXjhG7C62D6jsJRQbgwQ5ajXNIztzP4nZMaBBiMfmGmO5KUOLB
nPEapBYwRZHs5G7Y6BxUJV1s+9VCgzcDLkCdaLIGO72FwnybzW6p/YZCcFH9iTB5+l0Yym2Q2Dmb
QMrhlrOV/J4fej3uCm4TFO/iUqnYG5O+jwf7Vje3SXjAxkxA0cIU00AZ676g9ZUm/1L0bJoiXrhr
9U50C0JgSH2eZTBd0z8T39SCzGrmk8QNtKwUImaPCRCti9NySlZNYidwHKpjQHNr5w17U17H8dR3
vI6IBOvEf+yCpmaS2lHME3Zj4zScJnVk8lRKT7x0uvg0fIsvwr03YIZYEVYPvys64KC+nzwVjyOU
YbV5IimIUxUE8tuJGe3MbkIWIRrlVEYZrgwOImGcZ8AgLZxQs50Hgcy6I2Svt14kXTQoJSQYUxYg
6mWoZ3ZIVuC4/9V8ecwSF/+U8zYE1xJdY5c4rhoQoaf5CEef9aEw7JoYwDmJsQuGLlCrjMaqztqe
h1B3BblP3/46h6gGi4iQiV2kxQuM8h9yPSOCwRLAe8jVgk2Mh/UyL0LyJ4JcveFfZ6c2FLImHIS3
F9XaGfvF8bBvIRtYgFaIRpBsdQNLwqfU9PmqgaT3UeRkwVzAyloYW1OtBWwE+UxpEbQn9C/MmC57
lhvVAUZXO8Ct9G+C4ixHfGNHbhDQauRJBhBcb98doqa7PgP75wsRc5Oy7g2H+LHgbN0uh3Cu22Ka
5w/vvZwCe0u3V4nXeknoEVeaeiIMy6o5XF/+WPDs4VKh0l21uHH6Z+g2K5jAoXlo6RAHnn3ZYtIQ
WKg66qx6Yacif9vTW6f9Ae0CC2ZFS5f1wouTZWlaJ2ruBSjauBSU4nK38WBC70scOivdiTkx7OOR
CpQuB67S/iGDFX6KtkUpDASER5Z7O6HmY/Xo8piSs4LdrLgfgG+71do1bAh0gRTMddXY/Tv5Oylb
/nL5OxzQss2ZnVwhGUZsGc9zke1dpsFFa5CeCOUfk0od1eljnKhslHHi13HiFftzMalkIc8Crke+
MpQmdw+wWl796mt8HXBApd9Eg9ijHNKfQr78ZRVCFdBjcAsIBsoMG2M9efowUVyI2nodr7sPgS4F
SNdxIR5x5O5pKQyOH6agns3PMFdW0gPFhWgrwUXSE41Ybefw2mmNWpmiOLB3sfG8DkkNkNeUNR2r
fAm5snDHC0R1rlTwSkyX0RHST1MTYy2pRE4EN7wmUMC6GqHO5qrbaNAkKe7kh0AgJQNOWDhPfqXG
Omr6lGiRxyJnicNeNkOEhmddSgXO2qzUJpftlRXXLO50rWSaS53PEXzWKLJyhlbOX9SSMlzfFGfH
NsAbZY2jRj2tbRFkhH8Hq0HL23kyBKuuNt4VVmgNNCjeEAiMbllVrFEVv5FAp8Vo0YWTfJuBbBKQ
ETlaeIWIWlixMlq/QPwExb1MJi0IchW5Clvy/OQgK5yCasONU1eBpe2v5ovb8eQV1sNJkH25O34I
uwXYVXWSfY306/yDKhbsivWoIK88ZKTADzurSDYBxzJ0PTE47HFdAOs1pH2nZPHs1qrNBI5ahlDI
+fNZwP/YChaqLEhQgls3Yo29ViWn8fwHeWh6guqz+sCNnsMoESUdMsnrbuBuqOicN93mTFyOvm+K
nwUP2a8hVpdbaJABv1+qWdY/+W2RUotn6zQBZbsaypyDeb5+6mRgr6/SBnsosXHujCv1rXE09b4w
sfprr17s2XfRxqbUkw2+qhGLE/UJYIeJVF+OxAle8p8FKRJT9SydzH/2IPUQTyVOONAKm5+ax1OY
vc31oVtUI3I96xcGVoFm1MnQxvYUTYqScB3IwxnB6mR8RtxFy+HfxxAhok02mPn8gtKpt7Yr+N2k
P4ur/bBb7mlm/lgmjmJ1HnYk+ZR+vR31/4ZvqKITkOQ6ynSCBl7/Yy2J5HCWSvSPU/2cxwEZew8L
ODZc2WPxAEqiMkY31w9k6dWIDQA7KWY7uiMJGklBG8mpjzB62F6hefruD63ea5jaiRvp1VFvPToR
Tal7+Jzesd5Qd8MyMcTnTrM6oNydtMYdLow1fg1Ce404NAU3fTwGHL7CpKXe3DcbCod9a1pAmjbA
nh1svp3MMfGCXyUNT33UW6ohy1LCLaLsRu8iwtCAqDtFyS1kyXDz8+dajvzY9OjU6WT4nrHN9TrX
eCSnR2kWX+L+7dpOv++j0STxIRj7SFZZdZIXlZUGbn+tzcEcPUeu42TlwjVSnWjGkxsVHDPFzWxN
phvxbWR2JmbTEK+HlExgCyPXRhj47EtMcXXEJYhV0YkbTHqbafJqxZECMnv+Nbt4d9KwkaqbES5b
tDzXu5I7ad9l6BdNIZ6raoX1hnFI0ktPVvk3dtyaet82eBPbZC2VIYPnLTCgHayvSULUQBzPQxwb
qy+vZW/PldjJsFedhTdX0ZWag4Lgo+H1JotYbNnYod4PGU5tSqYarVdmNBl2tJOYmjrnoVzMyaSh
snO3CsIfuBGcD0vgjUIC+EIeG8Ww2U4h+Hfo9PIpnECxIdlswgwsYlYiY8qTFM3t0u1xFRXla2oS
d4mlDmna2zBDUGcuIpJTFwUHntYV/TUeVhcqM6asMQ8uQz6dUkJKSa0oUwfbHLyOXAKmcSCEk0dU
iest0bJbe1/BEY1clyBbxFnVaIrm0EuSyEyhNOHdPhT5p+QROCg8Ex5NBuJFYDMDNIdcSJ6Dyksp
wAit8M8cLf9487bakWT0orS5toO/y2k1gXNm6uMiJ2KEAwVfEJa8ZRPHu8il3E+bjoX0tW3LeesH
ySgGaZFF3KqwZqyytVnenjh1Zx66aa75NisDXa6s1u34F9gvK/fJVZXDd8B1omSKg9STjHav8cw5
bGqN5vHLWELY/QNDPzZlsQ979wAqOSzge95HTy62lkBNwI2z0y0HPETQ6QBzOg/wa6RQIBUg3Jkm
bcuj7QMCAgD+WzEwnZNYI0CZ9OOH6BrckqBqw2Jr4vOSBX6EVlRYVnhkdgq4OchdNUbnh48K3Lhc
ZRRGBKx/AuGAvbspWyf/o/Ib4DiesrJzvXLN+i4by/cz1nuZpVdXYFqKx8+r5dOhmjQ8qYzvhzix
QkAnIx43pKo4yQdugqWD8cextvXJ8ojcbcqaikKQAqu8lDrksL45X9O941UPFoNbOMDPKRZkdLpg
ie/Hu1KddsdN/Ga1njhueC4mOns2iQh56e3J+Zw6EmpzqwvBtQRwiBPOz2wktSQxjoptlRDwHZgc
K2M02ddvtoW9YAucRRDwB5MqCmgxKYTRmTBXYafwxjN670HGHjoQt7ix8mSTvJ1KWivB6W0NwYr1
29F7zH6ALbH+F5Cx78QL9jskZOGs3eQD0sY4whcG1gihoZw1b3Xtq0DyCyBPFKzKHJ7xLo7TckzS
VgHgVjARFNUCWUgt0FNCmJDzwmF8313iteaWVN2iuu8Q0qCd8vgoMye99Cj0YgGEE24NH1g1w9Sj
ve6MA/tUQRoNo62dfHqfpyH4ELacpC5rdVnmjtkc9MA4I9R/qslJ0kTNTud2QStD8DSLn8RybDY2
cSjcYR10FxBrD4B9JPfdAFTJfDfDBIG712QzV4uTjs/yOPcw2b24NjxmGwI0PgRXMoeVW0OoB47O
LfZkeV57VPafKLPuyf2k+tizqkQqol8i6gjL0kbJWymk4zj167JbJlwFZP0R+FrKrtNfxvfvv+Uk
CXMF9HxM+3UkWjOJ0mK3wqD9XPKaeymJPNy7Ej69MfeuE7hQeAM0fVDVnu/KHttYE/ADQn6E7WgI
MFszndWj0TAPWeL8yRna4mJ4rdZNPjrqnmSMjawJ6uYEwLnlqXvnAUYrq46tItlsOZxMtDb5rjBX
wjZZx8i1z76dl4rk9igp0WmpMQ5/NbK8TWcP6jaNcZw3wBUXA4mkSQ0VYAdOubZ1gi1flYp8POqJ
PFaA/tzLoCqniOYKoFxvavBhO+UyKJ6TM8Or4Pm03SGhCzBaX0E0f8tQ1fSQeIVVUNwoF0JSRVdI
nO8/tRG97FSne9Nd6I1OIwEeQCzsh/KDVFYL3zYp0kyafHDfKIV3Ed7rnv76kSLArPKdNmLY8Cgq
9Pjmc6Jljb7A3vjekdmPqkMMSLUV4jiDQ17+zqhGd2y0jHzVPtYIF5C9STUUjqpHffuyREHnO9A8
Rga8S0/wABBihLRwOs/YDSnIvjOOFafCUos8txnxQ6xWIfjOP9nhyPLSO3+XoY+0Qksv26YZRKOj
Qsd/4OmYCCfG9IsJl6KhN/UPYpKiF2sNfyI6ZrrvXqlzG6jSjlqOBDtDlkL/wbC4njfijaeFNvJ0
kmUmb2S3bA8vb3vPCjsNmediokCgzIheuP8aRGNYQXKWdtECAUHHVTJkp801Mn4v/GXxR6sVmXIV
dFr2yuENFoIzAd75TIbQMtt/mGwrDbjc8ZR6ztVKpToKrmykQ8vPYTejYR6b89eBi/B9X9aGbXJu
TvQ/vPdeB+MwCo25ta3lIBTxDYpP1HaAHdnVupwZ8L5s9wyx5bt9Vg0ZJ2rZ8qANKvEPjM724I2p
EM1Wn+qfNrjsnIGlxO593qKRJ/EBBaOWJe2/5p+UqQgoqJ6RCfAummYEU/Ty5Q8HcOxd+q9at6gs
7Jw1J+6LZYiY71ONkkLi63jrhUnByM3YQN5u6wmnXkRwaPNBelwGtqUO3l3W+JtoRqh1YrHdWHg6
gfOARgXugGmFKEYl1yGdLo/AqgjiZGfBQSjKzsFUdL2StfVgWJSBsFJ6mUJ2pT+4lbu69rCyETqR
y1iKvK4/Zpf6787rvAmEOpkvv7K7trlFE1O+EYlJab6SmcZAwZM8f4TR7S22juRxOrUWn7IraMZG
ZSiKas/4uC+MRUoX52TstmejAiT2ZrfanRZampLoM1B/iscgOoQ8YemHG/n6wS+6qFpI1IIsD8Dy
j7kS/HIDABw0xT3LP6T+KtA7U8ub9AuV472vWowUCoIoNMo2CT8guZnXNkVAkwo2QrBjhqteWzea
tQndQjb06HLpVIPaEPEOAiky457ZWQ2secIViQzLBmeqqKtKVLRefEoOww56/QJeAY+5udruUzfi
6CTeQP6ho6jwqzV0bbEy7dUK3E+i71W1z+DgewLGoVx6HHqDB20Y7wSYWgkR04Em2WnNKsVEqA6Z
wA79swoukNbsa3L3bSp4AA88WhcMUo5uytpJIXCGFhpd3rvg3GF7wiW/I95Q/ershzGoWW39NubP
aK7yjGDKY35/dpESImKNNoEv8hqAeU2XPVY2UEEFRBj+fokHTPTB7D90HcPXURLS+qUQMwdbsJEL
GZmsc7eQPQMt3qvePpIBwvVuhxhDxbHRGdRGLsPkUqVj9tFy9aqJ8SSeAzWsXnhFkztlWOmZOC+h
htZfVx4Lpd5pup8MkXwh0SG3wBUmJvTIkKAwPqx+ltWRY9zT3jgvYg1G17zNCUvzkuEx+IIfdQ/M
02y4SBZE9V3U7XrTJqqI3nJ6dX07ycXU2RRL0I7ExzPfX/SM9vWJrnAk3J3bpubfnxSKxdYEB8ZZ
fELm32vh5tDndqRvxjKca7uCeqx54u7+cyNWAnVbJpdAAKvgBGVUgBpWMlGs8x0mROY+Bn8+O32X
sbHDfiAy18HrCZthFGO+U8e/kUBzQtjUdx6FkJO+1rBeATirbOZZkl1d4dzoUgxRdLALTQt9kTaN
XnTxJSCARXAlLc6M0bjNk5XL16HDYcktx7K2jiSpMVgKgja7VhPFWCsWEEFs+qjf5IibNlPjk7IR
AuU3Jrksq5bxhLOPi/SVCBOehvELD4Utgb7uhxa5gsKSWwx84rpvHlaII6LqH+mFiH8bWxaXAAOj
ifCZ6/+QLWO8X1MTf5WfYmUF8LLIdWEP+iRe/2pmQNAy2E8nvQuezMVqPHCHqLlTu1JtDj6AcJJj
30fhEs7GLh/cCOFQJ7AyBAlSRRx8P3hEHkiaLtrW9XG8V/LvPgHGjpyX93yF2DYeN76RLNvxeDCt
fTcxR+o3hu8Kwx9x2LFmUPlN0nmj1/wNqw35ipAZVkUjCnxLiN/y78rlAwQWXJg9AtC5idjXeAZa
9UpVK2NMkiyhFEtw+DX0Buw77MBNqnpsya3dKD/OsyCmgDfrX3mP2tcM7Jd1vzZcW8314sHnxECo
XVRdt5K8dnYgch5s+3rWtvFQs98mmpyQ0G8J6el9UdWsJstFKgSF2A6hMWEf+pq8GdayZWKM2TWb
Yh54ZCTtqvKKQbC9lSmYJ82I/JDXz7q5fhPW/zprcvpB+1ExHzp787mowrdPg0/S3Qvseg236xsR
R13ttfyPB7cmjhWHC9BlflWBmgqEDzX0k+d+EJx8F3HWrwIfbmhUPQZDQrVujZufT2tz71UY96vh
B4gZrNdHcon6cu6M4nOXyJqL1w4wfK4soxfqdBxrw/mvDaumfQZsOLHa7qHsOjOALIh6PXuExFBH
sTEonCkTOCfye19H0zRmSuygG0My5s5IOd3nmHxkzNlTM0q3nlEc6RIJaTad5C7FYsZ6Lt2bZjo3
kgqiqmmSYHKvQkzMLs6MBskZiVnCHv6oWQH71yukEFzDo1aViQ1/STD5KtWnNTJwnIQP3/9y8aU6
o7bDEi8GAX9lE6qzBU277OE16s1f5mSu/UHGkk99bh5XB5kcyjlq9q5oMZnv82QODnRlB08+pAMT
d707UPjmkYq0QuELOE7pJABdtEVl9J5Y1xhM4zeqR1K9f7MLgOcbUPv4RVLBHRfvQ+f0611FttKk
6PpBudWtkZSRJt3p13A3BS6IRRKdNmRXv6TX2kfpy4+n+qhgJtEKFMbO76oD0jR9Huqnv1NVYd1N
BSEMF8VorU5aghO0bqyy0tiDoc16jtPB5DQwby18ntmfkmDf31WmRK9DXh3gmXFhxwmAXu7xEpNd
43V0pXehIwfmn9RghoB3Y9fpJd41SAGXyuTIbhNM2I7Z6JF1hq4INsdYFefF1pRtZ3Fbbp24NWw3
PGSGOSQmJfxYKa9kygjBrPkR6V3E2/Pmmwe0067HPjbFdpaOiKt4f7OQsIyw9x2DUZW0onWWKjWT
pJ61mHvQiHGUKLejaxGhyPFx9ohw0IMzK7EAeaQNnHys5P72doFbBULo54JykhJ0mr0MMG7Kz6Ao
NXB9sFwQIu/1lQrQ2W3a54CznyPS57+ApY1BtIFEQzdGtn3P1Twgosma9xXSFCX+axIpfIS9FdRr
raZCeXSH0Tayhwu5+FepmcO/VKfIgRFMnBNMVXj0qNfxMLkLMISveLAfPpFyXn+C2zkqN+3BxoZ/
9SIA9nSl8y+bcqMs3J6K/yfOPWKbBjgalD04wGnKNwn3xOAEwmszpfgf+yq0FtloMNcIeeLnW5za
RRW/WS5aVbH64uW3eQjfIz/PfMKbqcHLmR1FcSCeQwDtzUXn0ysUd5fjmoyG76xcb384HEwpr7Zk
1/kC/G8rHcFbRUl1wcIma51IzDbksq/Y+sJlxFv7eV80th4YkSAmtBhULCkdB21swrbmm2F1TbIz
53EDgqHeUOEaejQncuB2XE1vr3Yd79oO4Li40KCfHuU68pzIy/UfiRcfny/EoO6BzuC4+c0eodH/
3yYiotC8Nb46He6YjMJarq5oMtAm7PwIP4miD3MxK7/3DWgHg8PGNi0HVHkR5wTTf3GCEbvTN8Yg
OkTSrJMzX/1TFOqqmZKT6tfTh+UbBQSfRA8+J3MCP4szVLjzFut7l5iBrwYDl6k0+dmMtO5MmPAZ
91o8GPnYOEC6Uv9YViemwdmAurd/Vpq1l5x3ruNmcITZiMehpof8+VREPS3W43tXLcXyz6iaCqwR
hPO33HjHVITU8xzPgnGytbjRO+Lo7z7AH2Sv/Tqoq7E/jAe5HiueMdrlxgjzC82iuEtMBw4dKIkH
PCdLKeJ/cBq5upM/YkUDVO82EvWpQVDrQyshy7wmuXW1XtY29lP4WDhk5UqmsMYHHfvQ1/jerasu
JWS5NzUBQLMi5OFlyie2x6YBCWZjT4sK9kpGvf2LQihS7Dv65yz52Ea4UUXjJ8ftvFHBxm6Oy7Co
sZwEJ3xrgN+bFaNgIlECdVk3Tv9hny6J/Th9sVpDiiUoUTjehhKhWgEZ5bDKmbj8+llfL2AExDCF
FsZeMOTEqPUatLoqcDddo5B6lm8kUOBXVzGwxgSuK6dWMpskcId+mdtd9pfU6cc3rEW1NVUH06mL
WEged14I9vCvJGZbFa3UHMdFPFtrzI+yy0VAiRvh9ux9y9JeFjzVODTfF/qy/ZTXby9dlBh4Ob0L
LgilJgPGPNLQ26W7eGLkNXvyvx1eLfZByB5w9M6ZB8SpLJJJs10/9xb2LxH1uWthEBECn1PSuhic
FS384NOeZIM24Hqvaj+982B8XX2QDST1sqOf/QhYRmxmZaWOCbHJTN87YgsasSFXkLQ6slAgbeXG
Cbc2od2RqfLM02fJEGy902A5/w1ink9Xn7dJl4KRX01/B3sxx99P/sh3ON4RcWCLj32QTvv2WZdQ
YdYIgfKdgqWsCrqqEnflflabQ9e0CY9W3CZsQjrUVXJ4w6BiR1Nqsdc1BLeu8Vkz19lLrtcRnG5N
rlPHxD5B/rNEDJOCR8soi4/idMuTnoEca0/8Q10CaYXHu54SX0f13TvObcy9ZlIlINNYMhdltE/v
LX5V7GVRgjUv6I6LZKeZ4NmYKlOMeGxW/fI0Mxh6GL2dKNiPZGOZW83HcKsvNxr3EP0fTKL8m64C
ThX5UJjT51AmurqAPwW6GHMt5v96NEa0sn8X+ihIFS35ky7FNpy6OuXgYLGQu3GlF41AMFLUBqDj
odN/xkbaZ+TCMuhn5QytMQzGsypBK+rleexB/I9BFvFvrSIhgmz4M4E4Sd6FVuCBvtU7BvMf+/Ou
J2WtM3V5KfTaR+4diOjdRzDsqW3PcuUlZrggkD6P9BZwUGNqFlSp2qKQdp0GwJJ4+0nfulzh/4P+
36CuqPKDrDqqISfOdMV85pw13fq1u6LCiV0h8JWTyoz2v/0QwdmNc2GW2gRfdbkF/EU/Q04XGXVU
v+gDAxdlVfVhGT4z4/XoqSI7/dXqYh1n7BBAz3s7oUtaasl4PvLfYbqmaR4wvnwIsf/WmCHvRXxH
J1fNP5E2k3IYxxCP1zERaUVNVxXflTR3Adr5xV5+KfON24RFnP+1TdUKfNMdC7KeQt6nw3CC6pw8
OyItxu+oZT30xBftIosld5mZ+k3i5Soi6QO9HL+ftTv1DKi5Ku0INv7ArYJU6xYQJ4cl9Cz1I8ZD
d0NVsH13OeMKIuf+KzbMEglCUAUFOqZlJIybonv/REnZ3rajVPI4QtSIE1hZL9LRUxYxElvzjt9D
9K/IOtQ9jdGS+rUY5UpOg06chYDo+ZUBjSw6Sd4uIZrJprWJhd5lSyb4Q3To3Cym+E+AxoYGcNb8
umW3V2VwDQ8MKtUufWXTXFVjlt17OWWj4ubR/A/t8LgnAClpIHZXxzc3HXMIDVdHcFRnXXuoBlfI
msHdTQq+QzBDKyR4DSY7Hg+G0E6HEjg1OhXGWba2iTjJor97BUo4JOL4HxXh4xCb0WZNOfsO9GI0
312WQQpSunIc/5avhoyrXlzB3p/qT7XQUU+VPjo9Ug9dRyxpLn1mfD1y59XhXfRhVaAM4Cbpf4iu
lhTWfXAoTSFrOKE6l/HfcMk+e2Iu3AwVoVFpFW/Y7yqmP7YO9netbOFD0nDmkQlMGa78ShmXxpwa
NHrIuA+7oqobGbIi/0yBXQGRc6rYebVBvLJ7LPDA3DRpr8YzBLCCX5iQ/9/DrVqORfzj4nl+jQ/Y
y/6LjJIGllbQ08pEio7oTE4LDoN5Ga3lGHhC/52sLut/UdUgUryNwNfKo6m9r/o2dT1OdhtWKhPC
gCldwY6uCtxTPDqEsS8c/fc47hc4Qx9H+Bso88SENyHTmRfsD52D2VFtdhpzCAohgd/PXzg6FTBb
OqE+DbsltUMRAZBSKGttdn/Gj37q6j/JMC086fxogA4qFUHKuhD3XrNZ482qZ1Lcmmsk1ETN5e+A
QPjv5n2ob0iGRx2IP/KckkAn7XpoBbfpVp2x8gR60ZVoT0gO4W3VOur16CCG//8Kne8tmQm4qcGU
0W66iIZdJVa9RM3pp71RNFIKc6sR1rhENt59eHyUsdAPhJEtb3V4A1VJGMc3+JW1cuNJIfXdm+61
ROA6/niRp1yCsddX0d0HjM8EzXSodJa66nh5ZqiH4Wm7CyIwkkFWiA2ot09FTe/62ECsdNwdD0bD
wPHDpFmjcxq/bRLlZNV8EQtSid6BOquePqfkXCPQ06kknyFceKvoT8KpIJSZRloc53+wgbBWp3jh
fFJnn4dp4S+5s/WrwKm00dCCn2B6USEoBlphuXvk2kywbwwzVF9N9yLXlPli0TAr66UaM+IwKaNc
f5dcTNlfmhYX7Sj3QsTqiHEFMvJuSB2M/c6TyRDNS5vf/dVSC/3XO5Ojt65CINRAh+1AeyPOq0BF
Cm96/lYADkoha5rQJKTdQfNpwQV/Ev1U6nP6zWo07VGvxUgYUspig8A0QMk1x0+ZKSNrcAay3kZq
JyZuoxLFF3hn8k4IPAvl/jrXcGJFc5L8sNN4oHa7314Hq3ou0e2NYeMhjtm/CRxGU3zkEaVJdEh2
R3Mcgd8PQij41oHuZi9brOOsUHWX0xkuIq9yRN1FcqMSYPNbol7lY74sMKR74/dJei9GvEhwdqsX
teRWePb/PFtEjJxVFglRlSM/OWHJrfh4f/QhpzNd1iPBoxy+RUjAeHh50hVwYLVtKK5AP81+yPa+
PdekeiKzpsxtFwoRpf9aIcGuwYzY6Id57/hzfASlrU+kjtEO0fxkoIqk5rF9IIRZpNgKI1vkCP8r
xje9+QV9mNNpl6U+6kdHTKIQ/tEq5sm8ZkoWUYdI1sK0YvKwrXH6C4SVjp/dvu8pDfPOgHdSt4bs
K8Xlz9Vdme+x596+cjJXpZtU+BsU0h/C0a2TNFc1XK4QMBCKi0jFM8T4oYGnkYO+QfWlQpv81TQ4
ue2lVOt+ipbY87UPwbevc4vO/wIcbyvbG5lebpenke/hkdIgAgjeTC5xeFNkQgBXZmqTrFK+67gy
Gl1nHNjh6LcJCwJQCkdS4fIzFHIHC4GdWsjGpVMMnSRHhlLLHbdAvFFyjBk1lHx2Rr7fMLzkjb9C
C+WJu021IL1n/Tb2WAGM1VJU4Q3rIbAF6EV/fDyhn94vbARQQN+xwMToz2VDVBMS+v78CXjSA7OQ
oLrPexB3YNAs1Y2kJpHOny5xUiJtQiJZ2j7wxOgJ+oiuDx4DQH0nC319BUyEHyz7fu15a242jjtL
jKLKPEXB8leVpXeQ+i0KxPB/ECctFUiEKXDbexXfulkupajwTyOQucdVshp8EzjIIwEpb4XvelkE
rzbVHXSeQq0P7KZGViYpE74ICgZzyah7IiYtL4uJe1hkBM8yIGqEUe++UCbUM9nKewNnlLHGDzwA
MDhvOkbsYevJ210uwT3wmiTYW0ZVjRa5/0ETlm7fDsIP4IdA66+eZ0yUleZuvl2RWV16IwEqELqv
gA3Bsi55d5y5lPGnXcdy4bldO7Q2YG6cnTDBotA3feJqlfbZw4y2Ygeni4rfRUQRcwy5oe8PjnCL
+RiOC6Yw97hhmU/mWka7uPxajuT8ow1dmGyMOLO0HwMy8yTPrHmTOOhNcIcaOK6Kr46Tb1brNsE9
HrXDUyQ+Z1iEM1YNL2Re1gx3eaP7TF0mXT2bdRJzkkKeSsin57J3yZHrxIqbDnXcY3I05rqEwP14
s/bXI9oUL+XiowaZwL1mb1Oj6t+2kuNEHBX6l9IM0eL237aoFU5M5ucOE2LjH0WWP6VENM5JCb1f
4WTyobtLBDSFN5gjLfbvXDi7Crv6Fa/0+wA9+9Uk7DkRSQefLQk0bsVeAEFqDRPdcIF21Dz2+Mti
bwBHrDHNJetcvnaEa2QvTrr4gbVpS7gnHPEtP9CiBnaLTHsyL4+Lkeau9eq2PPAxz10RFj7KjX3R
WIitWacMf6lNFDjRNk8pnf5ofTxDw/dXyM02cATVMZK6e0eqL6Jy3brIoWCQadVjGqMskKXCNn+F
2JNuTPVLSHOLKydEOeR46MKRvsv3EW72xbuy/aMjPIcGtsaBra5Z8eG5i50JZhIGeZuRls7jvv2i
XIoFLT8mVZH1Ef/VxM0QfpcNF5KueaRZtNwYgWqwWjrysVSIVavNW4WPK1zpUljAYYzHSEj3zueJ
dUz5aH2pzeZtJjv8DItsET/RmsMcfgcIIJBzI7jRRYsuAWWEW4MbHRNN2yBLu/N347Fwtdfx4gX4
1vKJ4i3PCzG563dhlcEaXtps4Ym5tTzpKaIWCv8zg/YwscN4gct11x3tJqgWMEYrpDmEbiGnmzD4
5mtf+5/0KKAUbBoQYstHyI8nHA1ZMmQJIOO2QW1A3Agh38cZjbzmVM0bFQGcG4i6y2m9LLM8Ok+s
MaJNFMKn818G0swK4nm42gZTXXVD7mAR+KNTqJCpE6dzQcUvaMHGCaqFq2/g9MQ1ufs5wBGU053i
juNmz/1KuCwJ22zlKwDZFKoGt8df/AmQnMlLmpjT7o7GJ7aRtkoCXq9cVMZsXC6tiNFcBkUmFHnm
QkJISPp/DVJb0zUf4o3w48D0JdBo8oD7zkRIZLyCE81jZ9IJtvNzrwMe4CgXAt/h+8gtFOLUPSuv
OJMbrYSmlL9JuPh0H+tRxWQYxpP3eSF5ZNMKo5G+sHpaywqRPoTjB+Kpi3tTnXbM344AhbmoIe5j
BqArxIU3pWA78U5UNnzI61MvBXx+V1dtx10AQG1mxLtrM5h+1rdu/g6h2T7OJ43oknBKTAXRPmuL
QjBYzlVAnrDLKWEYog50lYyEHZMTI7GGLzz4s52PmmHOdg9Lxe1Siv5Iw+QFiOaYxV4/KxGVd14X
eyWVWQYEHvjBtkrGGJ60gGpjx6mzqB7rnqs4MNUe0D3iLAL61X1y3l7mamKitqOCnnR0+ec1Psdx
ggCZanX5FqFNAs04dkVwfzX9jWMWaB3RBDJDWqU7BlkySGHmn4C8+97OmumtfoKuB6dFet9iBBZ3
efNPBEMIBFnsDG/VtSNEAHtix025HttTslD4YZOQWOwElhEznQ5B8Zs28OmRz1uXPkdmqZD3RXEe
HL4jJ7Me+lpABTTmI3mNZv8yDUztu4FNLd9bsRZNBryGlNk3sFOzjn54mAZoB/7aff7a2Ht4uEvL
Q0V99xw8we/fCLDyUa2z1oqlyTK4AN8Hzs3z3k93PgnJw4+zap56WeuttnaT1oSqAYZM3JwQETzG
7sBUQYfZboR4hYlPRzUl/z9eaAt6PjpcZV03QWbS9pgAYzRv1gKSO/52Qlbi0I+JcCm7GB/9q9hg
zVrxG2MuGP992/PkPDxRgUzpyrK64JNiDtExyYXqhsalf69srYNV+q6xVIsxa6qm03/Q9W8N/7gb
eV9sY61onOrncEF/Eueq0CfASBVaakrsaJ9ilUA1OjYD4gUEFLopPtJnYQBY4sUtV/ps3y3ds/0M
DZ5H4eCOF3poDhjz0bKXMSz6MwY0uNs/qenY7fxHFPowIGc/c/78FpAR53lgJpont7+7lY165akO
C4ctlVqATOWTfES1vU+JuyqAwjP+MpfjQCamEii/r+9lJAl1uBlh09X+kMgGq6cFdtNNUn37DvL7
uh05k3CW43G/tejShuU17xwS0LFDNOk1rk2bDYg1iV61Vj9jhzY2wafzyObCi+BkbJkVM4jC+vdn
G4B0rG3oCeCpQhZa4Y4Zn/dx6Har25nisC7B7HQMtSlHtWv3bxnWusYjtAm2t0q1Fb7+y60uNs31
6ebB+Ce7dDO+GAj9VfU+oTQ//hazzUh8oLQMZrp+giEV2227n7UaS+iUBEy5dcIeZoQ0O0sHl6sA
vEQGUJboG4G4MwlzIOFG/Hzuk27IFI2ZrapK8L+x4xPfQFirSIomgN3aEvnfK9cVdHGV2gbCqsCN
kZwysAydRfq/RkEBso5ScqILBQhGLr8DaI8soqCVNQ0FDcODSUQqyYkS+7la2UYmrQsVaPJFvw9m
pBxPdlJDOSVuGaa2h/R96uKS4XVUJ6cXcmQwso7yfAiTplNtxfPvkaNeWEqTxYxcgIi4hYZ9tvk5
4v1Cu5n7LIYSPFB5/ipPb23opMn1RQXZE7JVwGvFXuGsvuk+7wuCUZ9scnkRc2GXuvuRL93gLwrF
aSUiMQipxbjQzYbYbft/fVWw/xe2x3LnFE+uvXMVmAKreezNd1D3rTKZ0AKisUA9EA7DRbog7qne
Mu/l4AJRww0BRujh/qxvqfXCIYBNRtyjbzZyTLm8oYQYw+Iuc/nQPyouLywiA7dHeBMd/rmUId7L
YT4hbe9asxY6d0I8BtEyFaImf7pcF9j2SSxrnqDCF1wIP1YOfjxMk3BTBljxfLOKoUYoD5CkAELe
dat2dZWAC38c3j3/oUp9ImcJlkHobA4StgB75w1hk4kRgPLFbyAov6kc/okE8n+KltKkAR/jPdlP
FvUyr03C9zO8IDYMBRs5R4WVd+6GbHBtVO+9f4eOIFTAc6geTbeyOr6Bgnnt2x0AA0TduqUrQr5d
witsoxG/+9tznAqgqQx3L4Z8VrHgVrvki0VlxRlNGJE6ZSQ0CSsZ0P/tPQ7UKdI03ZzyKs2UvGXn
JVgmINqKrLPxO+5KMePBms4EoVzoPJBTpC97D7o6HqklwdPbxbQhLI3jcuMpRKrPPhE7cXKsVOyQ
Y7WTpfO1yeP99Ql1Ou2ncjBX9HK/sZlS2mHzHpZHnnFADXXj/jGrNX8497baNIvBLMvoqQWp+8lF
j6BYxLFevpeeFJc/+TQil4/xTMGQQj4fbjrIOUzThYP7jr58Vx6ClyhrLXYawOru+n6GaCtP9qME
GWgYtOt2jxkfCelq5aEdZABC8hI3/dVQgMlvhVT4gRS1+yRY7KtFPSVBRZNO+Z/alOIrNI8MRokQ
vo5OuEJ6h7Bni3rw7rHx1A08mvdlG0fvNYtxbKuI8jQ9969VAonbF7RE4InHIjeNROWRqSRMWNOp
OF2NHzd+1B1qfhb69nKEwzslHsA1lmykNvu5DcDW+qn/Xb1jVizCBerzWxRxtk3cTgs/mOQuU0SF
2qYGo3RXQ7suKGyXLcl5EqW852/TTCvCdi8O/8fXnqOLDYifZEpVL9C8i2FH41/rFOdu925ibq6g
8iPvTh1X+aBUcn8UAFZyggbY8FUHH7oylMJmOKXwyRxEHLajWNy3RgtJKON9GU+FuneOGzRnK3Dl
s+k9Kygsz7NcejbN2qzwOo2Bas+5+qs53pg4SLIzqInB4J2FlJPCX+lrr+Bz47mn1WXVY5/yGRx9
NQeKhgSGNk8iPqcHwvz1MZT1xgxu4FaTP7y62cQ2lnuWI5y2Z+DROfgZK8r9oVZPiOJJv8Bk3elN
JMdDYNVWCooQbXu7xf2gXGfPEcF+qp/4nJHv4/2jWOOqwOyGtkqDBfj43t5xmlXE/BCuIWayvDwV
pXaVVORYYzIjlxejEcWthHXwjQEIgQhIR4HPT141cBA4Q7sTJM1sQNFVRuZO2on3OOfQy7NruSdz
2NTIxcOnk9CtqxrVnUM5aprxbS7+F3szzolDwF7Rry6dmsvSaCzBhwQXWFsOfnL4WHa/P+1YWmSh
7oiakkCFyZx5BLE2U1tjp/U1DmG7Hv8x+6UHzVdCE4a2O5rYHL713ZOSzULh9cbOOys4/ze89ai9
SDJeIS9wz3fzdgWhnBtjLfl3z4wzGoYIz1kziWkxfJ/T4xPgkEkDwzmJKvlL14jq/yHu6VIhZL2Z
OiNZq/nWUN35/Ywk105jwhl6NT6VxuJ7E93uOIvsjAqjy74D5AmxSyUn+UvSxQ1hL9PD+BJFbn4+
4VZlXx7Jcsz2MV7tG9ETDZ2seYu30HWbOrdIgMdYrO9YxeEyT5BWGn6X8a8UbuoRqW23PEkYWfmc
kuQfWeKJ8OoXASpx/QvDmkVmVudIY96eliSk/0k2gk4uBNm47Xk7lz/YjBBMY6MT/BkjPrLk9GVI
R2RIKavq8y9Abw6t/NbJor0ae47u0hvvlSO2gyWMrVWoJM+eHs1eeUaHhDNV5FhITfcOen3KzY9R
5lXVuVGyD8yavwKr0kLapawahnq/1Lv3dGzBtIMwKybYXAwnusiMg9z1rV3Ew1clUpc6BH5IobmP
hosY/3+2A2a7EPLscnzLjj5rGiOwxumU4xlwjTRzkIR9m9Yb7RI/icgkBgiwQpFkPhH5idsD8MDH
1Yq+Ih6cOFSp+UM7x9v8BdyE81y/7aikI2Ykf+MrR8pYUOGLzw4JufHkg/Ajonbbqps8uP7gYSDD
SgHzzhxkZSncq3T7C9615x7NY1PGN42opFwPxtu9VwGWaCFo1sG6lxPjMtAZG2HdSFIgdCT52STk
qi+MBdD8uuwdOEF9yo1fRDwtBabZCFnBIAGDOxVBXhXgtYxqPs6FoX/008ywbvDijT21avhZMUN2
T3GFHkrTuCDV/ufPLCWoDeJCL04EKFDhKI8EG69Ce4NYZ2cgnIDdQWZMZMI9q7ewZRDYi8QuT7Zj
89xI6Z6pTZfUFukpIKeQh6UbQMrIMhxsRAwunAJs9euyBvYQppFWAiF7D9zi1h0xYp24826ppRiX
G/ETbH2BtA0xbzz15YDIwpaxwLCEQyhGKPSDG0OzwBMn1q+6aRvrOQu+biES7DhJniQL62L7KDyw
VEQOQsmGUG/GIls/lwCPtOreLn6BGwapUrpthVZVwnG2PC031fjYfo4F9mwdDb/27K7lW+qupKzB
q4ADnYTbebQDKCryNvclClUThpFzcMysyDcgu321r/V7ZKEhL1JCLfHfY63NOICsNf3PCnWF+Zp8
2zRzFBDTlaFeNjUKgKgyJ15lOepNe130+c19u9pS4XiS5HNor7h5o1nAxtq43NvZRaqv2o9B+e7h
7/OuxhVueKAtZKvfp3tlFc+cWVzOIj9AiOCr8xw+IJ1v+M1/eiQyLH4xZHkYgu8z4vWKDS7B+m51
mButaRYS9ZWkkLWPbsF59betIlQ2MK6ytSpXtgMuUX0rb+mw7AxZuGadvWa1MgB6vN76mMBvyWcm
de9IlejPWEt90wehan/uaQrcg95OpwlyPckYb+Mpub/avdvH3iS2u6SMvTwJQFN2RgCO+3dayps8
l9RYK3x70CHJFz/BouSwwljgqAOnphgQ4WIuux5kFMJrUvNaD6aSq95axlC99ENpGc8VT4cPXscw
UI5v1q/vbRcJOmAGvIJPdtippi2LI8Us5osfKrICgkGSUHk/fTrzs1ZZ0uQjCH2wXKz/sKFROpRi
kvNkzzt0o46J93xBtrEZ+CT8z6TEsM+kGo9yj7Nzj6uHqjdzN22RJaSX44abjIZqvWoD026Z3V0g
VhclBT6BvAsje+nxDdwc0CgluHS71AUK3StJm/kZ/I1J5bYZSYa1BpBb+MfwgcNwTThqjztjvjLH
uOcLT8bXs4W82oPnoHwcSv0srcebXogtmIyYTNY5MjdpsFDVxtbQl5g4PSD88ljN+rKGNYg939Gv
U9YBwrbiuElnREHyh50OcAQ71VtRetbWXhMO0JOlp8Bss0CT0VH3shjz7wZpSFMTYzI5E5hiUJNs
TWp1rHzw/Bqyw/kK1nFqpvCdoZhXYuzvVrkWfpGdMd5/r7jZALxk+3YUzrgQTNsCNWkrosoLFFLp
baQ9NgfG+uzcYxwme+s7O+IqRwO23GCYmAR5OsegMTVUbZYcvjeIDpmEY4XDNHGpWd6dy1qAiUXN
XC6cJT4arX20WaNOdrs3NB3I+cJ4AxmVL9kFFYlNSxGa+p/CsqV2NfHfbxt8YkiUkrP0fOiYGoXx
p1nRPzx1HP6rnNOMm54dFCtnty2Cr9SAwLjWUzpkUQ5czYuuSovGGl98KnV7HpU9pzOyiuMp92PK
QLNghAXEyLhMpDuMYtRnGKG4RNJdFAbEIahj6F5FhbL1KALQJfOq0x8GTE4AlaBAx+zTdrGiBPQO
FUwWD/OgD8d6KJw1ljWh5i/30JHTIx68f3VOZn65MtNgQKJ5G5I9/w6J8ilIbVMKTE8q0Q8cD68S
7tjTx/OsHAsuxszxJxo7yfZZIK4f6nPQ0o0lKgXe0q1OgoYEp4xX5GWeSL41EsTAl28yoU87l6w7
0f7lYSzhekJWKOWjoUwG654rO356Den51bko7t7SnY+PQd5X712A0nMPEgjcdHH06mALGCtPnzDb
KOmTq7fBvTXXdpUdNQk+WrM7Id434Jjm7VxYFtP6vTAN5aZtbQb5XmQ28iclmU49c+8bLSK3zy13
Mst8Q0MZGrpoRza9tLQyxm0XWgG93MrjwtPc4xz7qidLilUXq0vySTkbPEWqVelHXUm4i2EHhdaz
z3Z5rpaHdu0Yrqby6YtrhOwxtgVSe3A2IUU0dYZwq06Fhx2GXLLF0tPQ7QnowurXl3qwC1kI89Ej
T7FolXJ06X3SgFkT/ZIhss/3eSYzyIWYYbvajV/SG0Et5tjOlERZx+Di5/LGd/IvFmc5h+Y8oith
X5zkbsupoEmM8d2zDFEfYs9L9Lss93/LJ0a5nAqQ4Egv1jMN1LIx3B2DxEX3PB+Nj8mqHsRp0ycy
xzyEoMc4VNUR+g1us/kDv0QjCVhetovcBPTJFwaO/JpJNeigW8STzh13G6V5KnvvzLq/H/AZDpx2
AEsZ/HiDBK5tjPOMCTInANvC5le3UvYjnIVVZW0eKOq1IU9HFbI3vnaXUIH9+8kQkz9ApMYjUSpj
NkA1U2CFJbsda8pp1L5Z4bRN2vqG5IwRw2lZsHmOV0roUv88h5rh4cAl8DE/HI6ow+COowqw7rKf
FWxr8wAZ+kjorg6iQGfbKRT4pbmxN74gtftjCCKjS97AW3MQ6+JQYOSexd0LNBONF9+BgNyCMUAF
Q2aQYHz+/AfpT9xJgERbJkFPYGSwW7Ep8IpktMy3p16O55Fp0i7TAaJ0JysUeSUbd3KBjJTf4EH9
2qP/5SH4T+NQxeCay4UNrTz8eb8f2jCs/E+jIJLDoQNPDVBez/txQVp3DHco9EOuQcXDkn24QFl6
lub+iuvU5HrtfGC4zqct8ZoUqn/5xzkV/i+1xoCXSK2mTrSF1t1AvlGihKJy1TqukUh5y5Ft3rIV
GcLkaf0I/wLmVFjhpegmbtLXiXAkAHTJ4pupgaxrw36YLASlxYI1km5Yu2KvIciVAB2ZB3YgOHOA
gzmiT7NuMstDt3pbtEeVQK5xyddrTs8rkAgWa7OzplchLClxaTQM7sfAN1P1mog05KLNmAcqSpnV
tORTgpJBPRbmthhROJeBkMafBmkx86ziqy3B9xuGJpS2HhEph6D4+ywGh3yCJa7OwLEYsBMy2Phi
T+ExVpTamEENeATeoIVdaE1qioRIC2LDnnxiYUXOlxddG9uM1Tg4edKEeKXQapDLvEEfvrcVpi+0
Lnwmr2MBhzS7F6xtvj/sFWitsYtFVnGcVHxrOClPApBx00T5vI6nVFg2s/mg2G5MH88bpa7scAs7
/fcLf2y+REHdcihF8/qAkhigo6xDtDhRPfy/k4Ip/msXq81IPMyZFZX47oujKcLlpRpXA5cGKJYY
TIHG+/5G6Nx1I6HP5Iq+LjT1kYpB7frVAipD4GaFK6w2qsgWkbK/bjx0Thq0RoVzrNE8l5PYEopA
l+gc/yUocd8kg4M8Gsp4/HxaF6Qpy/C/XGClJyNbY/SoAqZpOyFZgmk2qGceWnhZidbL+f6S/rie
6IRE0hl3sxYXDz+5v4ziyGA2n5vPSbgpgJjDt7Tue9tPDBUWsdL9uGD8WyTHha7ClmnzCv2IIKVH
H2dKjAcaoVQ7udmQlH29K9MRH6rFbZUGrwXviqrXYvlRA2O2y5LFBSFvlpCPQy6rWuT5ozgxvcDJ
S4RoYk1gF25BrF94BAu6ubpbsArFfqKsZHG5maaD4pvMKLUsYxmymSGNjT4ftLN5XROVIlJXsru9
V0RCUGAKRZwVB7CX9MRjssDy3jonZISv7A5XBoJD3zOYr0Ez84Ap+OAUpxp39sUWsEskhAl5VhR4
Rwcs3TMdoapICgo1sSFLhAhRrp1gUKwDP5C8PwMRlmmkWF2thADPfvKX6bdUZtRVcCT6APhOCRUY
qDeM3fHN2iB1vazseN5PYcR4Kf0a73p9/FFrLosjGANzHHcdHkV2Mn8XDYXbmRyw9tkjPVrhTCek
KxCgQVEc2yI7eCebIZbvd/boM4XLDcnHWdvtYTMJOVQs7dJp0y+7ZPflzhgzX2hTP2xWY1RkyZYa
FzOKf5igzMSiRRvYNOYTZ+B4+mhMIWmmEmt6+v4joKXciaO3smNCecUsWVesRxQg3udeds7Zkly4
3sAvYJhEBmDcma4xXynjKK2QYUu3GbYfusy1I6t2/hlNO2QcIipwlvXSGVCuCE0lmbhSG62XMLtp
J/cdxG5jLcau6A3X6dwbt3Qowe8+ZT2OzXIkzTTu8kxYco8gZTB3dRvjpwJ5+PRty8oFSkZi2vXI
Lyi5G/B5BUTF7y2s/NBTj7I3txMjOZ18oLhWQ1uHQvLIWW2cKv35Wx9WPzEp32dhsdhZJMYVFbd3
yODSdCIvrZaI0XnQHc+MqXXdusBlxJR8Eev5BZ3RWgGB/LMkk6R+Vvu6OMJkIw4ExoCW8ner6wyJ
SmbFSBvgUI020KqHftnXls4W/MFxaUqo1BTgLEGxf13l+g17TlA3RVeRRtnpG0mdx5+x3mszqCCM
VDoTjWgPE9bEuMELA+tBLA06AaK3UPJ5K6N2Q2eLHY4StR+YpOilgpJH/xdQYlr7NMCuJbAWtJTC
I/xcZNZyUrkuJya9s7CwHeNtiLmHgKKd9twmdR9KvfuqH43a5Ems/uXyDneQ8IRTpgrRv9DRxAJS
e6Nmg1Xpfnf1uk6xqOAItTVTc6BQcABVE9P/OsCTHeoH/cW8awlITMcgr0NRmPiySKlGfD0yougU
qb+I8dSX1IiIGALGC1T1xkSIiG3JiW+AXJ3FCNiFDA1Knfq2DeP2qPxl3daGPU1usRC+QzEOTYLm
ieaCCWYQ6tDCcMY24mUQ5Oem5bLat4INKu4vvnOqo9qANZW/NW1Tmfzx6qRsfg5U8wG4AeiELzpt
SlAw9JRd8/ApXkSqvAHgY3H/NJxJS8l4B1XwnF+opmSakPnPqP6a17kZ0WxXLqkzSKDdr+cpzvZd
ifOtk9npYWwMm+ze9XLsjqMrvDPOd+DpTkb4aoST9MaaWBqCU8+8sLXJcLV9A48b8qhnjVMa7eb1
NUDCWRxB/VI00oA0OwElX2RtOKiv4b2JCnmf9og/f+A/cJTuCeSA5NlfMnodbP8QfTDlTUesdkgM
qZ74Mpf2ns7kzFNlDyWGcx8Lu5yH0sveO2dCs97/o8ELA39U69/AI5nHqmrBdZ/B5nTI9rgKGiAn
q9PXRvYZzvc3cxc5q+nprIYY1WfzfoOBfpx7QuuvS/ZL+aC/SaLDjw+c74WxiHe5gQkUNz2fU/3v
qYgApnU7BZ5lvLiH3e5kDUQAdPlsRz6MHfZVPCjJ6UbATm7vtaUTvFJmp/tzPikxC4ZX/h/VfobG
VkSGPl4ficMhd9X0LKzuZC2oKc4CVoKnCfkwCK1kBZU1WpJnFunvc+/0RXID/NOfLWozes6OOSEo
k5mB2vpsORWdMMJghNrEb89BE1P6Vo/k1940iz6nGR2klRXyzPpuVf4jaR08JXnYalJ6rFB0DvkQ
MRY1Wwx69OgoforAa93RivdlvQmFLQiyw8MLeCJCqyNQQ9WZlOIXKJGhb5APKMzL4lWoRkrpVqUC
T9GXp4Vh1nN9NO8Utlf2MwbV6D10naaOpxq9kLWBBEWI5ZV9XrIsAmcqTM2vDlrfqWltJTjM1uvk
udL9XyO3rDiRqntjP8kihtO+wzEibco83QksIPMO8iWGjqmDm3oTEV5fKta/5/De+l+cEvf/UKwM
9SfmcFQLUyPGmB8FrBaiaUE/O0WuzL5OF2DEiCntU/KQneBrLKNrGTTXmapuN2WDRS8YLi+4Nfaq
iv5e/EXyNHib14GRRCRhwKtExg1elJRMek3sV3eiB4sQXK27USA+uk+vPYeKaQD2U2y7gVTbBSKQ
k8oHxqbZrzhAcN/ko7atL2KJRRE638zvJwM/OPnoHhvClhWIu1hDXLmMwNd+Xf+gVF92WEFODa9B
MAGo8GY69YWvpCNt9aBeKgqDKAGaCqPly89/x/xTLJXiRzxYjB1IOHAz/tFaGw1Hu2cBZxcBdJJo
Wp4MV4WLVt3fCJhaWrqzlpAe7JHniloMFS7bTz6IuXDvTG7Z+lyAkkHD0lW62QP5RnVz7EppukrX
lI8ZmDP/QfqOyPZ74k+c3ViFlwOLgDVunS0g8XQPOyxlujbmRYFChe9FjMIr/vVnA/TWgyYDdhAS
jmPQx3AhIeYrsjJlKrIe7NOThyVC1VkaCQsxI5FFW1gCZZM3FYKk41TXLK9b91KTvsDF92dHFatc
ctU5DrUbYZ11gxHttAivvvl0Q7RLdLsx0S2cJp2by//NyzSIwxUAjsAn2k3Dbyn4I0qOuqfb5POd
6S3xgT2xp8IBhJOxCdEjm94saH6D23CDagI5Wm/A6Tox/uRbb1LRZDlRd2qo1OxRed4OblPLNrc/
nsK0gESyY/G6B5MJEzZtAVT63mKNkLdkPhL2YbUkvwO415QXvPH7X+Ezr6rbolSPQ8KPCXKrAm3y
a4XHkNRyW/yMdaXo4oxMHUcYQc/frHjcAyEJ8xghiB0ernjWdPfuxT/73JmquAymb/PdVz50hvLm
wUfGUvP3TFdmBVHHk/LB/we6OAxcdXJ3a6vdqclppb8W4jdKF3VM1oUKLd1YrDJNPWqPePlFj/nw
tZvGFBHOgwfIJUSdJroQNgNe9JakQVGslGpDIrZ3+bvHnd69xVchs1bKtqh4O8O9LXep7Ed2LRPh
13nvDJPG5+I9UVrG7xu+9Ev6aJ2yrp5Xq2XwvNH9mafEYZMXqR6VVMKJKt8U/ak7mXRAHDC3b3fj
2vR6IqmS5xGKThV3G+NuP/LGBZ844dNEKUVx/NBO19Yo8C+C+VBW6SB1vqcBoU+/tGjH5m4Yx17B
AyfsrX8sT2M/CGGSAbQi4FGZYtcHsZK/OKqYHFvViaBetwBHTRhp+ArbH6OpYxHwDK/BYQcql5YV
XYOwjmfL8cGziTiZZo1M8QUrEdwb5sBXFDRBqiUfpptMg+zXnRyAjnNsoe2SzOLYZr05543Vk/Fw
3YaDZ/hlkq/itgMWcPMxbqayAXCpvwO9tu/XoUCJTzUK0guXL6EE89+dvMV2MpKg7X6E6aQzbhlw
LYig7mw93M3fKYLoecVwAWyQ9AVNZF/T3IJ+CuMCufm8um/rTwlfnvUy0vz0vyS0FeMj+zzvmeeJ
ch5jN0ezl+Lsxq5/nVljcuH4+gDe+mBzEfGDY9cyFnFAmsDzuZAitjxMXfayLc5kmz4z7pziE4uJ
3gXBk2woWo/noRnw+6HO8/dxIew/8kKQj68LYiWUx0dDjBAlOBdc6bvRwTd0z93cSRyXaIR0CsCD
iQI9V6UedAnQ4xG4s22DMAXj5omC2R7u93ljQckdiYW555l1yaRScjemNrw5qPjp52FKbpiklauQ
JML0SouR9QOtRSA5fGqSIOdqxgJrRhr0Vj2KL1sDJyDJBI+Xqt5tElNsQukDwPmxwCzmb9KmZqNo
G/3a2wk/5Fc7FYYhxPk1iQI+u0RY6jgxFR3Wbabntr9TGDWplN4bz9UylYzZEc/pMBpnqcxRXeDV
GDMrR/YEbkpKlEoTsPO2DDnzmkldwdDzptXrMgYPDMGTtFZyQY1PhgNIUd6By6mrEnTl9X1XEFOl
/rWphByMHxgr4NlXLM9vtfGm1k4mCrzI4XsuXSmGrwH2wqMJEDBPn40MuLLOSAJUMR0dEBH+BvE/
EQyibDn5tIgsfDSW27T4jhY5NZsD60hJMEdqphWuszjYRRqFNTpmuqpXyGKtPEjo1K0GzKOb3CnS
hPGlaFJGHCvTt/q/jKlzTKGC3K7qGDxyMRyVfuVO2ZV9IMoVALlBBvSCdtrdGeN4ym8srnq8RR0J
aBWg68MX0uk9WefUSqKRMK2QMlEtyiOrLdKLhkaX1rgN703EiHBC3YS4ioG2Y+lh/gpRQIFXKgtl
tAb0D7YdGFqKXGPl23hvF3W4tRmi0GDM1yolTFJ5hFm4asZX5p7uJm7dMWjtNgm3ikwOeQddNZUq
xTjZXHVbS4nw3MUYftlOOgJ8c1KoAicpsL/q/2Ne3KfxzwPytoZpx9g7wbsFVNE8QwvjIXJHYPpE
PI70QMTPemCGsWhxZ2ENGFVCxahmqZnINCO0oSUtLY6ehyvh448vR8tgPg8VwGy7jlsKzkKkfsk5
uGH6l1ulEq6wKahR8Wb4/UqAZy2lp54j0qTIJ11yZsf0Sqv90e6E/2Q3N4QUDHdRI0iUTHnwVVSb
MfWNh0uDBbEmNZ/acn6DUeVi6bZIdmDRXyjevZbL2LF7c/iVO4NXnFwfoPy69N684RGTqE+b5ygf
sfojdQGhPFRCKChBiTTH4yfBhioRO4IVdIbj/Nmdqylzds+OAr+m8m3EiSBaEQUWz5wAmZ/q7OBu
NaaYbp2CBp13fQIgBxb9QO3MzI1werV0GP/mqU7m7rzYeAnoTSWrEu2SPu40SKVRpIufmG58WabP
j9ahNdYv6kuyTSHJSBwoG0PGm0O+WaV6jGIIkxNNSbbxK6lEPQpBcvAvCfPDJGLqOEyZNQIMEBOw
Jite71Ox5xKhrYOXtj6U4RLP2I8dpdupbL9qH4yE5yIEzma+NZDSx2NQn21o64QXPnGbi4EFkOXp
0JaEIFLLgq7dvhSWvYYVx6jCSlp0ojAC35ahDyCV81gknApN0KlvmZZ6jZ0lhtL5flobm4F33yMq
SQXce0jny3YSp/GEBqXLb1X5xGS/vzJLPOv5Lrn/+vVgf4AVMmky3h2DUV1eezB1OvA2a59Gaf0w
maKBByRwpWfTCzjTfyucNvukKhNjy9+G9EdCAqLMWXSRdiSfoPOKSyaBo/OwEihul8dVXm57APw3
9+Xx2tah6Rc3IBsD7MuA6+x5E1+ntqlZiq42mcB4T92zLLNvEG0kE6yR2JgzUQQOkaS2yJ+kpB4Y
aOHq+gMz/ShRsIwte4TOMBdhLQyFBZEE4v/29eUQR9ZvJZmSZ2pIVC1Olo91TVhpxJp7In8tH1WR
VN//f1XJokK3N7FDfTgpU9VIVA+q+UdqT6ZZgw8n3CsP29Ywdp6M1pkmBdNysN9N3mR0sgejxRE9
w5XrXQX+GnQz4/Hf+puyzlO4qSqgLrpegzZicdwD93ucLRJ8lMc6xpqDQvNaOEohlcJtu4AFERkc
QmRWv1miaH0O6oEeVKiA9Qw1BXTsXCQ7LBQwCCjKbVG7YnBDSstvSHs0Wue/xB4r+mwTg+zHzQdf
5prlIPko6gfzXoGdusGUbawDNqjSVkKfqL2EfStLcDALgyMOf+UvCiQU45WzZTc92OlNuAyUrrAp
z5GPa99OKFWLk+0dRmGtzvn/ZNWJqIGMv6V+bTmnKv177+AULteQwKlORmjsuGEgsza6zgkJnUKY
TJruqrCeA/Vnv8LMIvTp6+SBR8lbGVL/7C5tVGAtb7YtRRxxySSxtAGo8IHNw/BEYLZDZ4UTJqhY
V74XdeyQaNDIm5xwPL2ZWUAItiJPCFeh7Bq7/2+3EniijIfa2uaT7PjeerAYeQdHGIGLaFAnguqk
O+3k30Qohnzsphz66CBY8uBdXWeq1qSe6PSfme76/TcGIE9LCa8wr1HKuAeJR8ATgWiZvPna0tCA
CFxkoLifq+rREVdf5YHfCwokd5UogSOKSM/vBJ8do774C8UuWPKeOKOZwavnh2DRuC3IKyW8G3dk
vZa5FAWpEO2QfU8F8RFiN7X/FN+o5uZ29xn5ZdXbDVW3gnEF4eCUvcp3b0qX3AHvcMHRV38WGA7/
n6E9U+KNPkL7dSOKHNAncNOTH+3lT2zh06pffwglRQ5dDNqcJuzIP8W6V/tfjaMJA518F1jvjKKO
r9SS91qlRU1XB2sp/KHAH8oZP3Cx2HMi67kmfJdcyAvG6wWsT8GpPSTTRK4w5cdnTb6HMjA1zTmx
LQD9HGGA6E4dvjt8XhAG+MS+e8b/QrFSH5hUcCGUhciYQw/AEO8WzsQOMt826fmJF/X272XgqXs1
7bXPMU0cecopdaoaJdw2wgY06rtIhDZC6J74KROR3DUFfMKTM8E1zUzrnXPN3SOSTVeKQgPigQbE
CfROTdtwuukTq67YMJ6gUwVfKhmvT7A+O9HV9aaurpQMIJ925CPQrK1hVMw/0kASd+sbL+XoGZIi
VwvHXkLUnEqjtdBbjFlikJ4g38EoMql4Cz8QwF9dnyNuIeGDuEek8+ve2McLiM59VvmLGDgfIxyO
VOtX88Mo2YwSkd+uNUt6QCM7z8bb8cOnp1rtL99ZUBRe5LF+Pp/j3TeWH7bENve9JWBdYVwS/KrA
eWO29zqnAGKscpljByjiQ75zFQNOk871+77W8y/I2wPUllVd2boPtdOCLNqCQ9rHEKN/t0YhTGZa
gZcfVxqoNpTSktaFnb6er3bvvXmbYBOjRKNwpD6QGuZ3RT2D86+T7YkT8SoWgEST90E0wIA/aylx
Md315La4nvpxfomrsPDGEVeNg7i8C5q98K9KOJsNQONoyyWd6R9SxS+HH0fECcbedBbHN47ZFDvo
jpbYK0TgVWwYMk8jtaVUYfEp6SMoVJoXcT58ClJQhej3gZV4USwUqHX3wGF24ZLYk4yTNeIJlzjL
A6OpTKl+Kx48FQttVjhv+Ct4syPAkVPCzdExWuz3bcaGYYHZfd7wTPEZMOPtOwFmrQcOgqiVI0fn
puQB+7gcllfw9rkD0dnYr57yObOw+Wtquq6Er/Dlk4cNtmq0oZHoSYm02ZTcV+L+OiOXTRECdBNk
kGlw1bmSXJeDDJBMyUk40lCdtWuRU726b5KDsLEX+qGEuN2W4aZfhOJfDa+LLjZnh4yEUHpXvxKG
/JYRxQQnWCv7MdECxQnQJ+91uXGHrVNoM4P7BVDOx00PpE0qHbxG+ZgX5YM9ejepgAQKcTrzgBU0
aLe0/6Ss47YxzszBzimffBSsMWvlQEcBSphW3kk+vMUMpqNLeOrU+UNwBDETUjrslGS7q5WCqiTt
mqU/2Zf9p8SHCIOOPDjcblNmXNdH+6Lz3okz5pmeH2slzRz9fQa6Ff4fYMVB618lmPU2jeV1XwXm
wTMbKD1YMnP4uSjGp49I732DwmRR6PMmbd18KP+yl50U865em/d4Fkf4sjUp/1NNuxii1HixbTNP
jTyWBxYYn/tOXnLpDRqLG5ffJ+raMlZkh+wot2Z2koVVsm8OgVWa2p5duP8XrdzHSPu+mFII7C/Q
6REiDJgHhfN/RTn64PuxqP5dBzbLY4tcClrDS8uCodR+Zi7hS/Wb2lYXw5ZdjX7eBkiRGYZeQgqj
Qf4XLNMfLb4uI27g7nukB9L4sVj/XOQLgu7y+MnSE3lnulQz8tXWNWIQEAYDOKauccL14oP+3tTS
6rckmjcu2rHXJ7ZBh0+r77q6G/VXpc5SYNhUG5VrQoCbJNHAyyAma1i1d9sBmg873PqFfk107+0Q
iNRe72yyd03NJg0LGkLZwZ/xIwS5JVA0GrPZwpbp9Y4yRcsxep2tIzGtqdgkEENuceRi9FK5QFfT
id42HzY3lWdgjprXYC5yJEJKMOenGxbYFjoHNe6pdvXNNt+PeeBf2t6YXi3r8YwSQxUjvbIeeUmC
NKC4CSfWDNmko73j9EITVHUMZQeS1y9wcwCSrUUY/8mpfMvBAxKrwdG6qIqsfRUsGWm+0GursuF+
J3XOLpkxQDkiRWBBEZ4g9fSWAnqqz8AEp+U6GIpstAEGHWytv003Sptp55SDrp5Iv/ugg0HugudM
Olvs3Oo6yjMUsenLua8VdyGtm/B5KyZrLEIwONVIPiXhp5kXDIFhpLyYWR6Z2uYsVpuM4jjCxXtG
nwTjNsAvjnmkDgqTyd4keXFDMO3QlmxEUJ1M9CVTp8jKz0on/T72KegE+/Nh/3w7HXkyWY/uU+dE
2NmNLv4+eNNTLxNgG/lbA2/0+hoOgeeDp67gwfv+nhkzZROYtVJmGzhGUq41DIuPsw1PLFHb9UYZ
wMYTJT2AFWcVAYdEFK7J6dFTKbwqrXunasPDxg1YZGPG8IyT1yffWRbDwBTpFyJ0A8Fj00RYxSD3
mc5jah9Y4JwWeqWAJ+JmQoQX8YHsG6mLcaSUtCexwBOWYo+ABNJ8GwYfkmSsuL5XJBXzF+8UcTiV
gmiP+p2n2fTjfo0DTGVMABZknbct8frXtV/+T8d21zeDKmTnBOXRdlUQPjxMUUOeZf3FBZI/YJtw
KL6nNMuO5Oa3HdOdD+uXrBwDqYJmHZbjZtFkTmaHOOwZ9KAwGEhBZN5+SC8+/fvlr1SlThO2sti6
Efyn6lSoAYO5kb7l2MhFmJ684Jd3rpfjyQsdnkPImdI5QVL6nP2DZSeH4zWN379V1xFKiV+F5WJ5
I3iCbZ5F3QD70PBgAPeh07yxR/ZJDLW5Jex5TyQi8q755M9GjGr3mBAZo7VBQ9Hg+lPZeTIvq+Qc
KPoJ7NL/cONy5hnZEt1BEVDGZjy1lgJHM9LpWTZenxCPum/P9IS1IrobtXUrHR5GZpgr7LQVwRqP
iFUgiFltHjtoSiR1WyVCVvAg58BBx16qdwJk2vw40fSeJ4MwtsQWUpUafXe2Vv1C2OZdi+KqYVy5
sNgyLyQEorNLIO6hCG1zgbAI1doGBknkVIHvkQdnK700J6R3qhZn2LbZ1eQqextkAwaKOb9Bs2zX
OjXO2FDHODxbt6iWBhwaoVrIZ7vQzYGPFw7ORLU9ftO4rpnMZ/Eej9aA3kw/1s5EyT78kqoDk2fl
RPskHTkCkSlS8N2lIAMg4mwbgcz4RvZvgl4iijZuTAncQynzdKQohPNkNS5jdwzKDIT2lkuRrc8F
nVyN4ofw1/DY1uEZZQRucEvXsVl7EJLvVk83vCB+oEdmkoQXOtd4VVFJMFVMp74xprtQOQdobVju
wfBpRZTBcENdFSmv2UMtsSD2XPLpckhJ+egWtEn9i4qm5XPZqt25vAIi6mSR70+SM5Mxu/mlCA7B
SGWSGk4CcC8YSyYZ/vvmWZY8GdVlwWrxf4PBkNL3uqMfUFEmQ9aV0WajAp4jmg6moue2+Ruxt3mY
psQuSUi8x2p+pemzvZXr5MDvZqi0uSdjik3fFGBGUXgCEs/O6WRJxVexozHtH5E0WXsa/qkX2pME
mT5jEpcmbHLgDpW6do3fL5fYe3Qp0fdx5oRRHsmOALbvaA0/U9fRzfjYhRrD/hIv0ahgRM9+8UTh
mMlCcRa1wHb6wCUNrRz6VxN+RMcBswiHhfGcHk5lWrDoFNbmpQC9qYeMF63lY62Y3M7GNe3NfZjM
LLfYKolTj9Hryz7dVT7t21G3Q6lhWD8GQh9l/NeKwLtCIFcqEVC9pOcCbik35au+fFREWwdzKphu
/UopYdQQQlyjSaw83lCeHDiRmnmXEELXzjuHuUPP01M1bH5+mdM4sCoEmigcCql+xtteCHmXol3p
13hlW/Ie3JXvIIGc6aNLRBqmrusc4kcaSXiwLV7Pj8LXs0OPwTv+ruKXyp5vviZexkhXJba1Gc5T
YkgWSQUevniXmKFdDxgzhTuP2ShuMh+tRm7H7Jqj/4aIJOGAWYD5J8RdGU/xKdo+HYL0QHOEzmi6
SPqMON9mIUGqNKcWIavOsrOE7+4gjDtTf8zDmcGLR9p+xw3BHvsUIpxgulrZumdCqp+K3/Kblz/c
095r718lVTgFNbSYzmTjHmFClyiEZLIlxeXHIXFw645c2NH+REe9EkGDZnvK18Y2K49MOVD/oAJL
gX+XVvXS5FMNUoQHNPXgbF4cErYLOy1MUa4Wg6Fhy9kMmeBPBkrUEA4r7MVNLXUFLwNTiRNqX9pg
HppzOi3kCg2BrH+rk+Jk3Pq7ZFULxdwm82AdPDYHn6F+jmZonHiY1oKxhopWpqYppLlRdJ4cnXBp
oQFysJXPGcekVwT4LCf3fzMjCyREIJKjQsDv4KokmNdVhHVFVyeBdT8qwzz4Y5beQRoQpF+1cgJP
46/omwoR3FQfGbSW03K5ILHAYW70kgb+xcCFmNUfxy/y6TK3msOlGT1CesOho3mmn8X5EpMq13fv
OayfJ/4uuRhQtscRvZZTIOFh+45iYAWU1ulgBSCC8yHqf3OgyIU5ibpOodnzLkHZFrIU0PcaYknH
vSfpbhHZaftn17gMlzVJl5mYmk54YPuUQ0usYKND01ZBe+5BCFThMto7NXjJfvl65ibqywdefWG1
Q6tnAj7w9ou7SSVLKPsLS60orSlDIzkZacssjJQzGzaE0ec6kZkyD71Ve0ODKNug9hCB88Ey1/+v
JQ/rekgy20TTwSEFxKObwLoBMbb0ouIY7OCa3cZ8Xc6ZIWI6rZXku2lvlmzEhXMm5T6BZW9EFI+m
SBrbHUpwp2sNfovegIj7usmUZ9X2be3TJ3IPFiK4Lqr0uSFcL7vl9Qcbeb56ifk7oiS6gJOmMCY6
60WKWhlZE6IhpEPnbSptounhckfgU8cUobY+Y8qP46BUNChoWCSz/OYtWCgGb5FiMnoLYpR9dPGy
dNBzHY7Pn4nh3QWa7aIpUKa8cEA9pU9GIsQkJbkOZ5BoxzXXIBQyPOaaRGTbxFu2JRx085NY6Jy7
0IXpisknNI0si+l8A5iqtkI/5oxHwzHdHkJeOStpEpgjtbOSzaFShHOPJJAkyTeH75G9DN78ra/P
kP3MjX5JvJrPbGZyWqb11C7LwffdxfmEc/s0hRNOMm/oSxMsxiEG731jhF/jlxHwS/+KAMt+ONqy
nLH4XRkfJBk298JCCgey6oR3kK2O23uzzx9WDVkCS416UvwsoYppSpkoEHTAHtgJZuXoQjC9j/mi
xbe8sOjU+JkaJ8EINen6TWmmDrKTYPoE+iv58+HT3mfg2LgAjeXX23yX5rBsGjrnFHZkasDxlxn7
G2bBoz78cbWefIvw9qTxjnI2CWieYqDHGOAtiJEN6FGuMv1I3HsAhNkylD1SWZTcvgj96ETMl4ja
kJprShFxR5/8mzGx0IGbp8rDIiwzfAMAwxgl20M1NrbzT3wfmNj8UDgXrZcGJGENV50hnGFgWUHK
uo6E1JWAwAayMDa5H2rn/futrKyupnitbxvZFICTSTyj2QfTWGAEoWv6+33BQUKJVlwoC3pEgbO9
enUMP3AwDjUMd0xELqei7v72vpFmH3Sh+cJ7fsmVWApDvDSnJbZdAKtzIG33HVFaZEMc+nvGHjJQ
GtSPzyn1oltSHxedNMCpG1eirYxOvcQnJorB+33z6+O6PviGytpt9eUgBrlmKv1jkJ8mYtwL0tAp
AgVlATfMkuFMKqIWUNvHm1PvU8xThxZpJ1Xh6OpCkoE6uIM80e59annH+umvhUnNuYgAh0BTbGPh
iC4MBpOvNbDq9pHUWquR+4N1YBX6l08+qahXzrtPSCy5l1NE2n3CBzqq7ZkavnDJcnXflp434fr8
JPPjU7PfIwcgAV/kS1Cx1y35RPXxWZPe6OldFx8Di6KKyMtvdfNL22bw5Cdbt0COJZs5V9TXzYOI
9zeuuUdzCb9zkqeFebBU0mszVQhKz+LR1kXzYBwzNapCp/HZIdvLzZXs+6wH0DZP9vaQjDOqh19w
n+OQNeKcyGbw87NKonVwvajxwiStPAagidozaK5KaJ4rLLfIAqaEmqCBLKMkxj/O2IPHzgVEKcfb
g+4/hwRvMm25FCeOYxDHxqebxvvoqOKBjuwDWAwKw1hyeFd0DgJaZft5aF9kgPnY5t3HPyNz0xru
CoNRXJkzCDwAzCvX9zkZsLVZCNoUzTuLav3Gq64KNpp75kzTHTbq5w5JveWumF8TqtrwbE6bKYYL
c6y+iZV/768arFhMPR+5xSpcp7BmEsNFno3BcxiOWUISiZkBnD74sOE2V7w3cpnXVU8R6dzGSGuu
FblvjoEDTlJKV1dpLtCdCq0SX6onzm3Stp6S06fbrXHNkAanHoD43UPaGMwDI50mqa6MSlN2a/Wz
cfftvuqczbdMbbOXf+6gd9zCbatxiHc4hqPfa/4MGxuXZpcwCEntP/FRKM2WeFEcCPK7dIR7qMUT
yqWeeJTM0tCpL0iYyI3HSfIWCdA3sXV/IPCBrCF+9rW1802DVWXpPqT0nOJqZPx55D/rrUbzSwNl
fe7Tap9ewpyPrJK2L2hdTR7B+8OnyHwkrmPPQrbtdK7f0b2wTkOGLQfD/CW7zvohf7Kyy9QZ8C+3
lQTUMJxY4oR8c7e15K9v+M33KhYLP7iAxIWpITgfqzezAOtTOX1CZgTh6H8xmQ8Z2JNJXmZBjeAQ
tYdsl5fm3d9RUI3hzjvdXvte7BA6C0qPXGQDiDUrD31i26BH5OSzk8qpfHV4aqLaunNuK/jxXVPa
ENyWWH9CQqfgTnCWtVf80siRKJAgjaBFIFYhyAkXo8UnaijxNSZogjgnOJpxO3zXOi7gNwnG2d/9
sYcV+yByV5XjIAXTmeGbqM+nqQkru3XsCWgJBrtvS0pZWBFyEFD3KrxkFGwnPfGEIVzgqhLy3Ewb
xESwK0W9U1DtIfXdg7TWHYNGQvjQG+kNGtj/tQVYQFPn2vTOZ+emlLMrtQ6a1NyCDjAJstT6l6SZ
+5LNycnrUklkf3nkze5VoGKKT0bffMDWMB5bjwi6uIpsZ8VyL4Rp7OOKOLyG4Ot0dizIa/kKHqlQ
ECUkxLeQOxY+iAifPDWcrMXg+e016S1noDTrywHGASX2XHRqB9+4xb0Ew05qkamsCh7wqY5q61DW
+s/y+C0SepNg4ALwQvv5q9bsGtTwWE1BFrWUF39DG7Veo2xkN3LP0GFvmM7Sh83qLgCLVN2lo/75
JKwbXI9JmHgvjm5/c7Uredj00uTCLErt/CHcNEbDncSPodvdXr3RI3f/xIlwdw5FeRGZGyXiGZNy
2Zq16Jb7APPXRjNPxnLTUF8Eq/LHxWbLS9JNf8o2pPiR/1nI2gTEHsS9KKLif5LTzwZ6wUy5K/Jm
UiydigEKBnGWFgvMMaK3DjG6myRpJX2qjlHdyjhPIFLlzC9l4U4zKvaQlv56SAC5tuBOUm+a+WGf
rvCFxMxVpxoJZ0rPFPis4BggJSL0FBKygBZNzubSvOKl0B/0rHJamj366wozy+Kung3QfTwgwReG
dgXH4vhBfBBOtmTGhq819SEHIX6zLwVhoziH/H/JYW9oawT3l7gN1y6GOXZbI9Kt7dFiQd0G5+kA
OQ2+20MaXXAye08uiDPIlqQGtBiQB1H1zuBVeW/xMfcSNPZHxvNR91IvwqbOxmYC+QSekOkheon+
GXoW9nKeenTrkWsdSF3sCTsnrVb/WmMG3dTRn+PuZCsJYj1t5eLbDif9o3K7CynBVB7IL6ZZBIBE
fT9KnB9rMkmPyLSVLheI/if8NOPj6u2gvijYGSh2I6sA0y1nWbzxGqKVsJMhUBnRu1p149I2DTMY
M0GGo1+K0P3rLeV4ztaf6es3XSIZA5E29Xxmk/WVwbLno0lW1OtwI9bCtMm+EtDsEIove1a3E0jx
loAWQ+mr5+LU8RdID0VPrSiogiy02nArv4Yt88XL2/YtqYBJkRxk14fZmKbeJZQFT0hLHsXtlu5j
m8/LkH7VLTupNpa+29OgLehCn4991LfjsF/1uixuy6w5aQPaECASyCdMJ22QW9bA/KHgX5jMS/Ui
mQ323sXBADtGwHu/j+RumTfjyM/oU4ddH5CZYDh6vMd6QVKaMJT6JkJxrWfLi+nPTCtnSDtCFtK1
KoaIj0OSe5fZxD4R9FjT7v91J0sARamXbos0Q3OfVhG3H2CQXp4wkQlYd1hoXFHXpT0mrLr9yO8/
apQqyN2ECvbALBADsKBNRTuHFcR6CF2HbdvG45lDyCyoS2M4WmGDHv+LOtshDPSdNhhhalWm64JL
Rw5OJ14MMrG17hYwg0BUxFrsmtMI3s6nVy5AuITBAHG6SvZkIqDntKZ9aLHLZ8bKusbB7khZaaaL
dcZwLt7PFH3gpsPxzSEsXnBn6BRRMFhKh8DNKge1SvPJNVoEcq8276dyFoLRT734njcH2D0LOSTA
wiqDClvvMDrSsmygbVNp+beUYey1G+DAJYIUaEsSIUlzbO4zywenoRxE2UZ3gNyxSgeseLjLKcCy
nXgTnY8BEqfwdxhVYy7trVyYiOU6q/0vTR/hypNEpTA38KqXJF/I70VEgYIVuIOzz3ah1eR6nmLR
1fJHXtcQKCAyWbKt+MiHgFNhQxc1xeZUpNfsZN5xS7kR+IxYwRw9cG9RUTqwr/ETBsY4ke4Ek3U3
O4kwR+CK0xpPiF/MkfIM5T4dI8soYirEiJXGMnvuOlTdEL/LqD3r8pVyI+HpVpimAdqcNbU1wYtV
GIIfD3NyLB/ib6fCS4W1c+Hu0JUM7HQeoOjeMyY2OoSqgFK6H5IUuJ5inC3ezUk/Y77wZWpXjx5/
d3sxJN4cuhMiT4nd7UFNDrHBfz5zKZZuq9B55i/GoCcZugoIz2TDMsHo4BcgJoFFpxALGSVwm613
y2qzAe0FfPpLjL6gIB2ZFofGU3nbRyWPMZgeUMOzFX9AuJPS91FyiX5r0xohvoppxwMl2MBaTKLO
WcH4lfNs2bPzPnRiN7qayTIwRNn5RJpxsbQOX3Iii+74HIA9QNvIKejcptlZEg7nVZlBwZu/+DdF
L5GyNZynheilsZv5lIBGiG56LWKR8IEwZz+3rkyDNrd5JZnEvoz7qArpeT5++GlNuZ36dbEF2m1T
QN4WaHyx1fq2gdFMKDfotrhTi6HIL14+DYtmMdsRFbieSt6Ya17gQSWOJYlW9V84YomigQcEHEKT
3/qQclv1m1OKZB2u6K7sdIKgvQAZYTWyoS94j9skdFf/gam7DW10cEOdcIVa8yz75eiSieVNWhnp
EwwZ8aiSRvxksU+MjOVFGvLq/SOaqfuVK5OaYk/BYEb2np6uZLDeFTh/7LQt40xEXnjsjZLaInZG
C8QUkX1YTrsP2qkXAhoEQvNcRA0b3eS/iTwPb+WWSh7MmhCBS9LK43acqnaVghKiVbqRJaCitAQr
Tgj0YzwDW2mPc3hnRgNYn7XebqBYVLiPq/bkJVDs5A14zVnXi7MqjGFED2irnr0elWHUvH46WX1i
PgDCMD/KXJbggyYHMz976aNKS0rqxt2qbRL4EZOsCWOiPIIyQUvWh3o7mTK9qrgGx6RKWRxDM/q/
Xit1kEeS1UpCgNPA7tx6d5Iq7sRVmvNgQzC2+A8qZzB3zPPAN71f63pE28nHM4rZHqmW2odEPDSt
yBudAEinXxRrw6eLCA+FVbUJHuKhxzLbQYfSKni55jsq65rsYB6JE2f8Ar2WZ+4ZqFri6l8uEvpW
KQEEvpy3qpW/eWBGsTneWm3latJtKtSOJ5DfONOWC7FOE0w6Yjz0sAyGbHhtYVtvBQbOJ593Qfzl
DJJdDCcKW1AVqCI1mm6YimESsJuHkw8i5MewchBxgAtPxb+1XBfxWV7yonLnqx3HE/BNJDPDvxx7
ZptIsZt74AXj+NF4ubqMOKP8xlFhIy7zAUj/A+tqf6Obglwr+p+0pTDX8vgX0lgwCM5C+bqjWCg2
HtD885sQQUcXXtMsH5Uj2TmLb8ck3fBm7anYg9ywJiusfUcSUd0/tUZAk6Vufnu6CcYhljuPLE3P
wQ11vT+Y7p0JdHXOvwTKDl9jqIoE+zQcRZshka5DMG/q3pjEDd4wMjre5y941QVSQRzYQvf2LukK
Vot+86Ddobe1SCHVTU30OIsmEIBUnofUw44PeLbAVe11pO5xyuBuTIEpc1ilNxFJ6BN5ORY5WGxg
kkksbOAE90FRv4LgD1u74NaJtcVXdmsyXbhtbM7qviuOwJdV2HN+QlQozF/PWN24mkhKWWaywvd/
RmtZjyJ3Vj5A1CTHAXQ/CGmi20c4o1PaJn/oSU7NOIZGkZ3TBZOFdrKElr9tC007e8ux+Im5cr9M
EWkcB95MnbNgE85tHcnp+VMz3xZ+LpUuMLrmonIpSmNK2Y1+s0MJoMJTjbDeUf3uPC672OzUSwK7
zsDCljthBTx7uSj0i/fmnGA9W/f2fpQDJk6p+8fyRKAm19VJhLSoCcasimlRZzDQ0pwHK8zmaSXc
rQbrtJQHsO+6m/8fkEiBakg6Aq/h7vDgQvPuk2L1c/ONJnTbsLXUuR/WPm/uDEMkjBiLMpURLvG1
jWVCqwx5bGGipxFZ3f+hHUOxYqU9uwiD/DvqQ6K7Rxv3n4ZtH7CTCcoHs1ZYQ6EQBcs3dDuMiRtL
82S+NyrkoVuCqVNmAodpe1mKEJ2KBl1dQTHI+xHS/vcj717msFJ7169QRhQQErG0DgEfRGvL1IVC
hGDhYpBXIi20UzJxYqn/7HHxdu0gR9tk+CHF8uNCJcDGqz05puwioXXx8jmTZrropwRq3sA5/rLX
AyJqrHohCyQCqRvH70BF7ZIWnFGMyKrVK6uvkcthst4pMvtdU5AU3HnmJX9v6/XsHB9jrM5nnJBm
vobGcpzrUYTGbc7df7tGyalPX5R5qaRVj5KnC5Cprs5bpnApsfo32wgmi2IAooOlTyd6/H5pvZkF
mxLdX9loaTsEW1jZPXF2CvMW5m4HAPTqCmHqQ7PUWSmeSbvz5QZHuBEearQdqARTYdMMJW5B2b4N
G39QkNCgb+fYcgL7X/a9x/nXEbINbgXmVuyISr+aj+dEOZkIg5jpedaiY1A6erjGDC4dUoAGBnFg
SomyxtJIOfjzYdVqnLJj892y5X3vyitRKIbimgE//x3BfwXRKun2h9RWOAOG+dG2mUw/nXR7Gbox
eL7yH0EomUWGS7IALfGNlMmeHftFiWrloYMBI8Nd/s1wxGt9phFUf6xBQWdcRxQtEheGOT2+qppt
bc+HUADIhxs9llL6s7SaIoW1Z4CNitrzeNtDmes+0RUY6FVMlV0Bz4+wA6URlVAW82FHUgcuhvsi
K3tfboExm7oX86FFOLHnIooOJh298eOLAPQFDlmXxOYJhTHsguZX+3Xrgu2TgRbjRFgK77YBmZ2w
5gk2kzigcL3Z29wjCJtTssnOCp7sX7z8I5GfYINtZcj6J7uPkVZ+MJEU4Qi6Gg+YJ7WoBVLclZUB
Vst4ujUrGtrA3sFBNpaZCwLz4rtBASsw+Grvq7xpjHu21OwW19RjFzkNAu3s0aTh8srra84DwL1f
/SkegI7z1Rv6dFe4pwAi667rpa+qbZPaxcQs2ktsz94E3ZAshgDexfw0MV1NvTYMi0uyvSZ0mm8m
kaTfxXFh/YVrlZfy3aE3215FZ9yL2/jzF7Y3B4bNAXT72t2AFNsuiEorblzS1YuQVllmLeNLVZFh
GZTfWXxEnq+4g7hfY07jNneQt7ZmKoqN/gA5phzHqd+jAfJfejqVg7VRJpFv8mjmmjAYUZCznNkp
TCkA/h5OTTHOqt9svemL9qh5/FGJ1KxNyThVT+Y77MgbQL0HcdFx1B4rJTlfifFTa1BZY5STzGdo
+s2edMOHwHq+ECwwzfU4xcvyPiOTWfLgK5vqcLosXYbS/g1JS9A9edk/BjIF4nPkEns228iOAUTT
jI1SCFVhIP/oQ6uyvAjowXcORS7Vt8CjuW3nOfVlZ8RU01TIiywTbAixajkcKeUePS39ZfbkzFV1
PAhRlhuKKlyI4iuDjePGF/Bg4+9FKe0AMYXl/RFm2/wOqE8zvnvlSkTSqj83S3bhBo4UvHq+7vMo
0VI3NuQkp8rAEiYe2KW259Yxzi52cIctW/NsJCw4IngtHFLM3ZKF1hZgiVse91c7v3+j3xH0Ka9G
XJ0xpz90M0Llw/2RlRQgDhPuJYOCfjOh7zQUs4rdbIoEv3J+LeqLXZhddn9E+t5mma3JCzjzDhMs
APdLNm5goE10ij3X02f8ofui9PvnWoqSl7yYdzO3Vj3O8CsrOULUSt8OrcOXlUVtIwnBJo6FFO32
aEqElgzpWLJqS4kdkDcOHKI/WjZky881OrApAGoeGXC9nnjsEgOseR1ACtlpJO9ZVNt+tOso1YeB
A0IToG9sreheCL0CT2aQfZ5wnOBGrAC5c/5Zgfv91zg+AcDSvEG1Q1BKdr3aK/7Myh2QIx0uUrL+
GU91qK1r/yJMKlxLO5dgw71QCpd10pXfvVYQ7v7NXxozfhrcbVGAqBr6yG737oibrUEb/79mGbDV
iC2o4fZQwFt3BQhbaCEZT4OCk/gdH7iu/pDI31c7asaiBDfMA3fr22G7xAciChG0d9u3GBWejIY2
EUeeimXK/+i/TLGbGFqwf/cm3cIiaExnvwybIAneWvDSB07pPFKP8YtayOZBxkIdLjoCnYiAuQRI
w7Bx6UGqQQWIqVMP2ym8Xm7hUvkZq/H+7lkl6eAcR2WUKLQhErczCO2GH3Oi5pPP88NECbLob/sR
uGFk+GsXF8potMUOC9WSuuoZ/Zqff6rHiyFNE1Q4fBGV26ZNfDKXrXLkO2efnPZcF6Ww3478ywnH
u1ZSA7YQvPFDFJM/akhDNHm2Ckby/H+kJBIe/XAEhurDIB5zA9ZzTWQnVYCNKKNTgZXcccSvSJ7G
uNdp76+Sx1Mv59krpLirQpaynMwgJk2lpr3i//xGyEM+WDozbZVdKNs/a+U8g/hhsebIU67fC7Cf
3DeRab8I8ipaHv5Oeh+OO/MpFGSemT+t/SJFcdezZ9FFztS+YBFz9Bej3HCXqqRFnFwKWqWjVIhF
x4BJ/Aso9ZCLS1r+pN/30yBIsOtq//3YOH74hZEGOw1JQjHTSn6BF2BcjZmK9YFaC59RNu+KN69s
jngQEEvzSJlZvPWEkm4jYj01POfNyuh5plbUnUyVpvssnEv3nRFXVjQ2WLTp25Vtcq5Abj/WIk60
omXJ1/tyyJa1ZGLJkxA0qoXhJX1QH+TPqhkfGiccQIn36e970O40cToA30dN90kRvwiHRLH2hMIE
pOll3yGMVLwBCVjG8sfCUqBr+FI7J/8yaNVx/pMDyJ72/O+HKfB0Xt79OsyPQx4PlDNlITBuYyFn
45St3XjvpovTSkMcpsoXO+BuRUyD/F8zFyIf608h0F/kcdbXwiWIaaxRTb28V8rpH41HvxGIKPCR
Avtwas/GvbOV0FanZBYdlYVo2xSI8VuursI0D8zJ8Uz9czHSw8pPLOxEsB5d3vYBh5Vpj4lIGv7a
TAJ9z8uDh8MJ2yZqRM2rBQbIZtJcuW49vmCh9auxK9j54bFgOAj1QSGERJgz5NcTtJCKZKsvY21e
2nsu7JIlFobwHqMZrTD8BytBBnI7+wfb+wqdM6c60In2mb9PksXqQtqC0Bqpr/aXzzXX8PsMrjKA
fiC8jW9pmLLzZchDwv5rCGJ9UxuNVK9x1AdsnHjRa+CdtP+BRrEQ72ryoFyZj35wrtNRvcpVoCzp
S8fU3ivYGDLrPRex4GSvRWIxtRCw7peC8bzydn7X+2r7lo3hO/wF9sCxjSBADot2P558iHO6rb7/
DNemRxeeOdCVZpRrqwhpxtNHcJ8Y1Lq27lYoUAGddxL2+Qa5pv32HXLRuyZmQAha/pux9Vg2bKOb
Vj23KmHR/fS/TUMgRwV/hrRsDKLYvasjd0RaDtcq6K8AQkwymg6lIyvecl6mkQo9ch/485wpD5dQ
EMLY4zWMnIQsi5Vzbiy0/dwsnddWtg5Gl7fAUwS5ZdyrpyfuA7zh/X6nlD6pznr9CIKBzPZrgk+7
2VGur3n76YTay2vLnMoe/rFrO2k8bbUW6jSIqxPRtFcAwvAw4CAAJeUKgp/l7WybEbqqJkvUGbYn
P0dgm5HjFirap9sI7gEXZ28dcj11mWM4qFyI1GmNuQq2E8nkwHYf/F4vRBedVlBAUPe7BvCVTqo+
Wj2mbXCpQ5DzJx95Ay5EU9JeFZj+nnrnC1oB1nKEOV2QTs47dskybKVbAL4sSTAiqK7K1L/4kp1Z
agzG6C5DIfRqwlz5dzyl38F/LG2Gn2u9M2101hSuc7YeOovHdSqyT5MOXo+pjoS0MhsYKog69IGO
WQYZKbs7idMzM45litVNW7wwOcBLt6YJ/Ggl+dAxiLXw5vVYFsQM6QppgMtptAuawdDA/kLOQ5p1
s8KhM/+az3FZPi3ZczNoElDCCfmdeKavc2pzb/bB7MGTGkqFMsd601B9rxhLItKbCUktaXsAFUxO
xPh3ah44DCX+eKhI9l3nMJdnxOA3fuKwEU0EOIdUFjtn8XuJ0cIMYGwHmdFAKi7d5glbnPUSTT6H
hWVYAofdprb5oiYB6M9EIpFwiTuBZOUQRb2b1uYxO/ZyBoQBRuCvVmhDiHmRWJjU64+CeJ00yzTz
y9IKWAVBABTfwp5kbw+ibeuMY1iHBY82cMoLYH7i+uXDXLn/uHp3D/tlkhEpvU+fHbi5PRQnh5aL
cezba8v7e6ZdsiMTbND6fEiVhqtamnMulZrd4a+yOpi0zZ94fiWzHHfbqU7iiDr/EY8VyLXN+8TT
G6yPBAwqT6Ba2O4BDqF0Sdo/Yh1YTfF+0Puh+F8HaIQ5lHo5Lra07bRUMCoym+d2ueSxm9bPBl02
prFLB5Kb/dvRH8lt65Dq7s1w7gt4xgSMEu+c7Wp8uR+5pMS1NmhPGXWOOa5sJpUvILWtBtcnMg/E
kZaqV/16DukcOCrhfX/hSC80W8NSiLAPk60FNK8L1DhFrkGZicilri3SkNG8Fvx5tnupQpCq96k1
nfYEr1qJYYa6V+wLHdPjqnb0xXPq9oYSS9vO4ygaxk+lbQ10OBzGiVHbo2+0sFvxt+OkQ80A68Up
BtZSi3fpt5npo5NGjVGk4EH+Sz1R2GJ02TMK3RzfKMd9rsMThAt8GBRRXLe13gt0odCnfzsZSW1H
y+lVZG0jUBehLlIH/NT6lQLf8ZdwfKOCV20TWzYyN1PVpEX1JVfsWgThyI7O8ES9dbQdNV+qKrj+
KjBcEl8dDugsEuOMXx4GktJqCj3sYSvzmZZHRzz91eGDLqLho7CkeCuJG67GfurBtsvrXIultGwd
5WS5DMOuIuaq0d1YOoLdS/r/VSPlrHew1SaTJVDwq9lNVDQkseemWGvEoRTawQT10v3ngCnbcosf
Sr+BumMfMG9bPIyTbZzDSP57zgIOwy6qavc2OVY+nnW9TxCu1USIkN/2UqcJn4LMGUiw+ZZLd2wS
/s/qP1cIRhxAScldZwsoH7f4FYSQKjT2gDVd1J6J/jOBtNM8RV1AnQ+E4ZQWJ4XyLDZZi3HwjgNJ
MzOBvPbXok8XUn03Z9niepMD02IPLt9nthm/X+wJMlyqeM9wiTegnDb43LIfL/uPH2yjs8GEg6OS
5p1Y/JWMPeV8h82Ly5LHwvupid96FpGrSBtBueRDNA8Ngw+1LdynNeg/JMVyWmNFxRPUmVICbgaN
QVhIH259FbUJNNWz/6hScscfmPjY1iNgfUnew81pKEMMoht5jERurS3qIyYOSLgVm1mF0ke+lHuj
ID6UsUeTdGWKnUCzcd8flxXIP/4gJLnsAwfnGFU7y19q7vDrxvmirokElFBKDiagklIP38lkoKyn
wdYLDEfJpwoQnQrzg6qUbNXqjS7Uh0rVKku6xPp0yyZMuB+YOjDlNxE/feetBs0CAMKNF5E4aQvr
VXAtVJdW1ZzL+0y9CFdFxthalWuo2PoXwrhGq6p3UdGAlEv9v6dmY1RC5civJetlDvQpW3uRBxbw
vFC5wMBoXpX9Y8b57G1yiHoJyVzj+QemnilyPV4qi/mxk1+pWLDuv1cz3dNiji4AOS6LMsNaA+V8
ODjlrP22CoLLlNk1PN/pQoU0s8/gM/Eu+a5JmGSfuP20SLcz3L4bbws+uFpWo80tZojdbxTz/1nL
MxMdq9dr7iNfbCFxd/LXGkBBQKbAORsPdn+NCgzOZCdIkCqfLYOCgiHh1VXzgvsHY4M4Xemh9BLD
1woaShi7YJG2ira3Jjj50Rg7pyBQmMi6lNebLWPXyxXuhjDZpYxDHAhV9peXWGr2PrwuS+2B5cNy
gDFrRluIEpzXUNGfdIrhq7E19QuPwSz9RobxkRzDp2LCWDWVMQdT5GkicjxQtRkkfQUevu3Z+REl
WadmsIp+hZMBox0pV4+ExMxB94+1GpSeoSyhcUGYvFflDXskXU0ime2SYOBt0DSgiU+d6VOXt5lF
X7RZXqoJwSXrSjCbgZzOIzFwBpet1FfoQT4W1erh1LpJXm+5AFznwpeyc3gcKj2PjNfiOAN9876U
cUSyLqN2qHN0tFoceaddFB7utTMB0cSxDEoW4teZm49CdFfbsqrfcUztJhpbMlrxVzCae+dBM2We
KKkG5CuEjwtC/A2Vvt+No4gaB6wC2rwxbD4eB7jdwiZptkwqR++uVj/3G+ODYL1ykMPYa93Ccmnt
Mp8P2S1u3Ru7LKVE31DOxePEMUhjEwcm9ZG6MABtAbfrIVPshnPkyqK+nPcmw9jB8eGT3C5UWizc
1AGorhuCZQ4pdpCOZSI53GpK3TeRGDFVjHryVKvErRY7deguN8zRORXd70d1AbLidmCx5K0nJkYw
P4hyQFMO1f8UCVEiN6SfDWjVDDHzxuzVxUAUJ6cBxbg2YzzaAsQFsSHOa75hpz1iVjtPpR20hpaM
NC1/5ewqcYKmFlEtsieNf7JMiqhdPVTZRURHIq6XIz9Z3/f1HFf1daTsva9KSQf/3UPNwQkX5mPR
8rKa2Zb91Ax3xXzgOsHihBjvATILkxMkHXmk3IACenQqFUKj7g0OQyp4mIS7zqlwH8Buq9TDzrSY
lmHahXRdtvN8DGVnDtCslysHUmUEZJaprOGJHVmQql5J+sxoKtGf8bnKnlin2ZcasxFvXlt6GGYV
qC3C0Fpgln8/0VeRuWZdUuaYtk0GBycrQOtgymsYt/Op5sOThrndt7rnpNnvmAQxh6CII+qDzdKE
9sjJEBFr51iXYj67ZlEi989BoaqzGahdn5deiOC8J3F6LRbgOIB9D/DXyJZLAw8c/SJQwnTOYVbR
rHIWNewmdYaUXB9h+76CxXoLU8kz0iEbPSNrIpjK3kOiNIXqK8P2zVe0DRfdgWc8HxHNA76CZlmE
2SBgGmfTkju1j60ZKgDq1bliHA6VsEAKJjqpc1LagqjBnq5ci70SoRmJUrUZxYwqoHYRuTFX9hAM
+9kcxcs01VdLUoByT8ZE65KZQWb817XwL+AKybhhT1VLADWVU/60xI20rGqmfHJMaejc2mqS7WK2
xDb5L5PbTctHhMdXLbD+DEeFUvQHTOedXbP2+8mkNsK+t74fngLMAghKoVQ60eVbVP6nw3tALneD
Z8x1PS9T69tmAzFmU1ih6BjK9RjoXlDM7ARhPH61exX+d1xNn9b2mJhRT9g/aOueSe7OLwut7TVI
eZbqdqrnrb/oH9ZjocDeqgvGdEabY/D2XEcYZ/PG3pM5z7XRwSyb7RDnKxnnmqmyOlupbKhCgIQR
2m+WrcrBP13Z3NVVBBjYlcrQmTxnw95TWtPE5oXKGYlLpEXI0Qc4BnuiBZBRbUeOWRIx2Jft3yik
Op+Ryg6juds72p18CZoFDS+99bN41m506nxitx/fG0Xk64EBriGhZxD8UINOohdilVUf/GSDRaS0
kFxSALV+6FYQKqJcqg5jwwWRmroIcW78zJK9r+DoWmGqrNSwhBaPmwKhBa7fxeYjz3CB673QQ5qz
fDEV8/TlXgwXpfKdI2wILzo/gGGD1MW8VQ6uZG5yJWgW4Wy3YTn1MJcDnJd165dandwINStpcJM8
tVwDWKObWcXJoEmCMTBEuiZbtOGVMFRYYeAiH2EXxiUA7511YvCuksVBn5azNFaV0fkBnVmyIm17
YloiIpvuY0legK8CPDTLl3DRBQTt80I42V4TexryUJ6l08dj+frsnpcOtYZuyneI4XwRsSXHdP/g
ajNUKH+Qawn3zpida6MVwusARbH1Wc2VjupW86zzTs8OeVozgOhHA3bxx/nXKK1FQ36xl9C8aAWM
Dgkc6NzAR2AqAij8gMlEtsO1GF8Q3XQG9cBmmd9ogLcDyTFtVaO+LhIaee949wHT6vPkNS2vXfL7
wVEMe/YX5FNebSaNaJ7GSMTh7GrSjfzNuB+O/bipziCgbgo6455MQk4ldRwVo57m2sQxPSFrhNn4
YBEuDFSGyi2OOXTWvP3bHnKYrrvxpnhdqcAbDK6DN2M94lrDNMChiTiq0s+r/hzQHeV4j6RZAEL7
Eeu2AVdk913xT+cbUtJHO8t9oAmB2NM4Cw2G9uamK2KXj99UOOOF2nq1CBSNbVGuqCFIHxWvbgBc
tNhMFFpja7YJRlTFGHzuwlmWlu+yVDFU3EFJkkdjRGp2ST7Aszh1eZk6/wNh2vw+1e4RZSdA2AgO
OgRZHaUYn+01RBp5oKFfGlrPiNiTdn7RVPnpGPdLgdRcvKAGTeWDvvUP83N1tc2X7td04svKBHZo
wOlYrqxzp3E/5zpo+a5P+zPkdnqpRO2d7yzCCm7GzAoBzswSPawRZqkUEYBfSJ3FKhGbwWVLyoKR
IJpZwN86rRhHC+/a7aiGeXRycUzg1Zq/iZuCEJbnHjUUmTt4mDdbdDvKu85eDaWO/3BFIfv7ok28
Z49BWReGRV94WAyfKeTNORnjQ5CnSJOjbZzIyW6BK/pTfe+i5nOi+hSa8sT2DZCDdV2sPsIPMpGu
hKWmfGBrnU5xutDk0OeaTUdtt8wXZnDBRE2cOGAgXR3mu9MAq2sR8mAFFrX/9mcQPVzEGPV2cDrt
onT6OPoxHVvmcch76IbnDg6zCBDoSE65fCrRNqu80JpL0ivKjBIxaaNVQAigxTU/UaCIGIi1xigz
3QYjSqoAArepCtKk3XdoGAr0Px4LG2NOYeWbbDlg00ehTtyv58v1Ksw5Zze3f+yQtfnje5q+4ILc
voXMsgEepLLtgJdUuY9/8PXUqRYIDQR7wEawvYuu8qYfhXd/8ga8zTyfZzAoAobkj5iI79kYrzxm
y4f9a2pn/5eGE5t9TOF3cEpxkXsgNModXFfVPEk3yscvgVEtIe/Sf/SbEpKonNJmLAGHYPnYk262
Pfj889EK34JB5xOVoszcSeN/CdE0qR8XcVeUiBoqnFMhWTGT+kxgSJpvXEfN10HHMSzamCxjGWXo
nFHfEXIU8Wa697BtpN0MHdKcsuhRDaOXmNZd03SaFFE4QX+xit7+NvLR6djpWqSlDuXcrcy1K/Fl
J0U1oUMWPS9gKlAjUJbzPvcl1BqwThQ66dtM6/6Ix0Bc6vi5w0I0I+2GvqwwxDFX0MGXSo+6KNws
B0PTQZZAiwI6Ly3B/RAbd/NE4qYi25OA6dRIa3wjm86ZR5ndQF0M/vd2HRGD7aIiFHmOk6savWvw
uA/OtnumBuDnRxmxXsC0WGDLC6WwzslZ3kzUbM3M84V6HMT5om7uuDp9iMYhx5d9AVVwF3aI8leX
lpVTGm2M8UF/H9oz2cH4VVKl/JAxV/YlnKtKH+PT8IgPznVdn1ifjzIi/7RaX/vg6U+Hqb2Zy98n
grq6wZZko1bYhw4P0wU1yZcO6YAF83goFFTlOzxshN5BH4WF324C20yOCEhYGAWoAiAT7vgxMw82
O7I9KL+HIp3BZdoMJqw0X1K/PPF6ecfUn70szcjXlQgn6ANzPGqsGJ32a8tu6BuzTIjNtvVM99iK
H237Aiiam27OL7RcJcZ/GlNnr2kalJEzxjMcBLowFWc6b241LVREFCfHiuFszNp9OSFyNlAAtfKZ
Rvt3u9kbuBwDLTf3BdCvxMrgSyCy8DyDzQSCVDJrrkkk6xuoA80p/s7J/lXKqF+gELGnTkVkwjk7
J7zxqSy8q7dyFl3vIwYxgQIja06Nw2E9VtLXer3GmSeTvvqqzSLl+5AWckmnkFdq6D4/3yH5k0Vu
3fotyvLWYgW9dJ6Beo1jLE4RRRoQbyvAZh5fkd7odvkvMEycAqdKOz7K3Z+zRX04PGpUlEwNJQhI
AFeBH8ivoYMUJbW8ufKVTs4R/p3r/x2U4u+I8otPDLkOpSptA01zRgBe8Ik23WY4bPaL/Zn/xrWZ
vMfSbAU8OjbW3+Lj2StPQ5uTgcsUjvqZQ6t/xeIWjsmrbTQRwZkgXuv1NVtgDBPp8YuFgVNnN9XZ
wDGOt+wQAclOY7WAfExVO/JPT+NDmwtSotrv9FLqBD1GfGInbPLNPrLHeiNwvE0L6fUfnKG89E3d
dCAuv1shNm6UysTEBnCYdrcaREfLPzQ6QGMjJ7V/iE0sTiqFwEW3oB1t/8hkjx1MTUWkXkEXYtKf
kd4TtlMZwoONCzEFdzxJWvjnWOt0ByKbKB0aGgm0vRrz478Oo5ySFyjQGmhBhyGmHTKZHhuD0PqL
yzpnl/sIQnmEu7YXt5+3JqZgFzqtSdGr5ZdKR2g8hKiEUdW2s3zDStKyVhf6OTcFiUArYmHW2Vm6
nacC6JIrKVrgi1K6E6sdpWzIsq0WvEp/dNeZn9LBq0/D7XzT/ApGSTDj8yfKdJaXYK+Yb7X7MCl9
WQ6z/3fGR54pmI5Xl0aXkZaGCRT9IBQ5k1sX5U5OioKWOD1bjlPSYV5d8sdZxMxeX87JCbZy+39M
rji7z7kBRlPKCf5G8nDg+C/erY4+uSj9+yDYbVklJRHRn39AtfYCxK1i4lYEPTbQ6bDM8YSMP7zd
VLOSWSQUvkzJHs8gwaVvF4OWOBUKiRMR0zvpjjTF8SxuEccA/SgP5WhkWEG03Ym66zUVd0o9ZR4W
NMtwnw5yw2KPbEd7ZNVy9iRUQzgugR80q6ta+U1+K+W61sw6DtmVWOY8AMpqJ9/S8Sc8zczFAK7p
VJZMYoczPIANw/RX4bgZiJs29un53d9tOhCaYOZr1FzYVxfesVG8/hohxA7qWC0pO+ER5mSUo1E2
ULFcV4Mdh7/B4Iqvi1A6nGdn5uHKtfEDsFYP9fYfOMyonCSk8V4f4XkV4Y5iZPiB7rpYxWn2W+z1
DdQA3EomfvOfuYovoYwF8SE8AQ42bX+wfd1+cDL6USlJ9Q0Fp+R4jQjp3UIWS6e5XiU/T3PpEXRx
P9fQ1h8UinGvRXjKbmoXQgCuFnFlQsmU3JcaKLxHF7pxiu5kXZEIaTGHWgwYQsnqvcB4123mLL+o
X8vcTkvR6AhaMw+nJ+e1dC7ILyHg39VH4uMjpC8/VB79n+GGpqaYjKlBfc1uitrottvROTWt1zjf
BK+AvhXrT9wL8E0u5b4QfFGF76QQqBoVyMM/wL/rt2meCcFqf/yeP1lCSzCLueU6WSZfErPj7Tiv
O/jt3g7XLwU+bAPekBzapBsyqFfUy1p8sgeRGTjR9dTNeTgJ5kNQmmpYHzghFt6/PGDCc6Vdk9Lu
Y4fqpJsbOza83Ty5IRcWISkhFjbfBVxgJ1CV1reyJcHxKtSjL8WplDPUxFHknI2UGC5u0szeDnwD
7//gZDojgjMyA0hoFU5VOuiSbbevA7Ev/3SxVaAYStlaB0UwOm5kIdjpP01e5KuUEiwpLt2jz3k+
gtKbSouEfP5+8aGdV0nGGNA5Tt0NPfVR6ObEVEnP4/UFLQPPzv7VvgVp79ulckL+32bnOG6K1xjv
ovt9jnmjfAlyvOpUsNrh3ALndO1XKWNUyLBmVQQylw3cPKiOe9tmi1sLb60kHPdYEkzr9CZye3JL
mSN9/0IPlb+RxO2dsltK9vjvnK4UIsS1AzTrBhjzrQTAUlUQCLpAQTjM8kqmHEtZ4hBi7PE2w673
ca5DMejNnnKmk/bsNxklqdZIcyiqQIqciHaM/R91+ekFSvFcW3Ed3QSVXb6zMZz5HKtfg1ngAo1b
7qApHpb1U0mtd7yi9c+fHoe4BFsJz4Jjk2S1YpyoDJY+6/Xum43Ok2re+1JPQPMiWy+kUQsHaNRa
LTfgxqXFq+gjDIiVTEd4wDA6+xFyLU0TkHIN3EyXd7DjCPQA9aCxLlx3HvIzJrmTC0nTG+/DCkNO
iqOXoE1LeEV7Kw6Nrkf0N19/0fWa3m6an7JI0lTIkBcldLcbgGY5dLTDtZVqorEt4WZM5Dj/kQrW
xin7EE3DNT+bCdSH6ew5goyZKYwNJpCVYnXPtMELAJ7/PvkI6k7cZxR5UIIzqpxs+63Q9nPcXsdl
nMkhrvAJNtr5N125ZY0tzmpzwKZqUQnxbn7MCffAolrBQ4+peAhpQxGaehpPqxODMKADfiJYURm7
9Jry+ro/DxR6PhbHNzt0/J3LdOc5mdGZ3mVkz20DXrCWqneoACDwuwYYKQW970XYoAGAcCTiXUEM
wZa50rt1u7VkVQ2HthuZUkgCL3avGopBgsCnI2OVLBR3IzJY9lNOsvVZBrEqPEGEzxNg8iuRzkm/
J0Chbn/RafVRx3zVP6omVC3yD96H4pqizQ3YWlAOqystvjH02mN5yhIQBdlLSgdC522buIVJ4dIc
IES8abPc0Md9mFbA+8FTBMvAWAzCBKg+QkaqtTs+eJsZMSixy+PQv4Le0Hl4SJcMsZ+3PJsTQ3nq
36gA2vVXG4k2euWp+XPivnT6fBbHdcwbkblgHLzcrA5BEAdt5VU4jDOy4oh8veYE38YPx8en6/Cq
CiphVxiJaKOuBGzvp7QQ1YMxbo00+WGPNQDNOmJVE/gltxR0vJkM7SMa4yImjjfzKKkfPQwfE6C4
Joo7vw9x0DVb8GU3xkkdDqp6qlYBKsd6RCCIvrJoUybn1NZ5+IKo+/VdEGN4EU5NArOqpy0M7RBb
VurOSj219pVm6LHIanonGcQvRakcXhZINPAVIL/+Y+3YKcRYumWNw+GXk9cVSIP9X3mtLGIfL+9B
8G1c9vBiDc8RWcWg5nzh41JYkLvOa16eP51FZY5R/AGgGL0MK6cTNzxBEJ2i4cFV07UqpvqO55fy
rFLlu9d9rFgqqjoVLtgv9OjDMcD8Ssv4sJLRXhTdFeARIjtkvu9D3+DStPf3UmcXjH4hSqUbgd7S
XsOn9l0QfoskNzyvSxO7itxytxYyG5KsVcp/DtUOtAzzTIM0+hJ6sC8oNIcirZveczIfTu9/trr3
Gduir8fjhOShjKjLWd8veKEg1pV9+TgSnScoXKM78GEGhJmBqDX0nwquyC/N6rZNfy1hwdSbuNV1
MNO2WwZQXtIlvI/Wyz1pgiKfwmnvN0g3r+7TITclGEcXIMsfWSPRe66IPHz/cyjTFyFVWQgcyB6Q
kKhsQUzO4xTHOy8rF+ZYhoSJlfGbA+vday+XOp+M6ljOzXaBgAf/49JW8XZsKz9k55hUXJ9T38KJ
xCxKsdxi3IeL+k/+Rgm4EKaB6d/m86GPOhoiVVZxOeCAHq48tqVaHpwCejWh69k8XGdmfyTP1Gqu
wOLyzvhqB+ojjYlDyz/QEudWw0zHJwjwMhnrnnAtk/4SqWpvggGSl8ByJU2tClQPMGtTR1fSBjjt
8K6LHw3SC9Ojb5sFjJs09p9MzsgLX4EMfZU08JKUDeZaV9ahcg0Z7O3cFYiXpgMgYwhIvF3jFDwN
k/ZGp6F0sUwImYEaf4Vla5aPfpdXbtq9woZpr4jJGYZinEB2OHyYfagA0SltP65EOaEYsMEj7Ovy
ndkqcGBsbOjARhDsVMnxMSSWBaqsn2fyAQKIIdxOFXuXwSASWDo+Ng6BZKbfUjELakAyctidCTMT
SYnySsLQrms7L+ET5uGlt8DNhc2anWYKoP3C6B59qAag6xrnwLhdSa3d5ew5maNkxXXbg+eY1l76
nwRCBhmMeJKLZo2BCVOBxeXVbzC/5tqwwOs4rEpKVjyvJM6HiU6gmYyfRYf/J4nkpe84dbfltpal
JJ9LPWW2IPAaSnKdiDZrF57mRvENJ5ppIfsu9eb2WhYej87jhcDrpvtLZu0TUjHXZBY7joaXCh76
n/vZRCtZcEjLkd89BBg99faM5gWcHe3FIdtaDyRGVwxt5pikXa1CaATGHKoMrkaTmJEDYvUwo9Cj
XlgFITvkCK8zFHRX8SbhCv2d2L18l5SN8piFmLD1h7nnLpAaoQKT3D9eXoHZ1LOSiZpeNm4ehJAc
1H/vJPr3Ptj1aRKIWlGsxxTxrgpNLQKG8VDrQbiqPqrno69a6mpfIwdjTRQRoFIBO3hQMkJcaXe9
OwGNpcszjWjSns1IbYR8Llb0THxcaA+YE/hrpidv4oaDFbpWs/U76XAQCl85FegHkw+NxDjouz1w
Ut/rTdTLv6q2p9d/voSpB89mYC2vLlDTmqi1lwmgLGCj50zer6RsdSItWnSTeU8gIq3A5ud8CEom
F8lUlWYK8W9PM33THkXsOW8/Z4mwkEAeCyhozng2i7OrgGx+2rmemSnAsCrQgcgigduLpsW1d8F9
y4/woRWvpM1xqGiu6xmpOSfim05JczduzezR5orPylsNQsjX4W4HsiqEPLlh5HL6tZne71wdT2FX
6UNlIbIgl0yaKPLP92KQL/lpfCGkLQfi/Hh9/rKTvIFeAqtgMRyTwmLz+cEF9s6K+kpBi6KfsazO
8cD1le4X24FKFGtjpFfDjq3Ux2vGog27WvbgfzEweccgW4jrNUlNoioNChTmptajd6sC79y45Zl7
dQKtNGh5NBAVYiqkI7qF7C70KEvnD7w6rbDgxXH0mtaY3siaDKHTN5RuOi+jmzGDAgSZa0YRiBSo
Tb+85dadb07aeP7/MDeqU7JlmV8+w9sVEVbIK2ZElj5V3FlP+fbItbPCPmfvzc4sSx8CQvOGkL8M
lrIqIREQoQd0iKTahzMB94V8nFEtpKiQdIPp5YQN0OBhmT745GHvLAuyE1mdJWzKJqzwzibDmFlQ
hY+0caxBD0v+Lzh6DWNikYTs2OOAEdZ8fDVNtDYihb24YCN2Fbto3+wrn4dMb9eZLMRKOsgq+Wzt
g3wf6bTFlquECsRVqj5NV4Rs8/viVaU+AkFZdM4v4PF2cGh6/AiS9SWBLLZSCirFfs6nAxbZ/eaJ
+uFXt6/yIa0kozBNhNuh2E+5UxuWdWHJacNyn5NByTC2deDPLGqZlLT8nvq5Fc0TDnIwotH/k0Gn
u1SMqySfAE0FSZ87YQrNl9gOhOPX4XiCknOhmUVk6MLuuQszxo4YRNszIJznZbwyGC7UutgfE62V
HFOuKjxVkMp8YYAkl/Y6IQw5EarPx+zk64iVIWb8JJL+/14D1uqU14OPbblZAfoG1dCRvPwYK5wV
ScUTEVI7q7AVfyX1jStKZoGbKkz/ugn8jd2W0/t6v0KRUo5twkzGMYpHp1aYSgRSnByGZbuVwgwm
YNE7b43XPDb4n1A+grXHBE4FVYtgK287wI+Frbpk3x7XymILaQDy3jnC3Gt70oVub+U4fmDrC0Wq
NVPUGLHK5HMIn5kkQc1/3gqTEv7WZK5OHEGWWXL7Z4+rHv6CuSSngLDsAdzlvALDb2Bgceyv3j+a
XgOcgw1OD+FHtVvYRNHrRf44QGuZr33hnqgTluA0nXy3yp69QQMSkaT3u4O+p/7XE5yoWWR75ftp
AgMIIorwLdeLbp7dQDCDONN+fcPLuSolX0LhmgopOB74O1gPVVr19sx5hVZgj+Z6Ieoc5g2Gq/Dg
yyjCnLkGq7MiFu7lMPtGq5n6ZGTETSEZMD7PZNbawdC+IHSmnr+NubusZydVdejNGsdKxIbv5uUK
iB73kiu9a1H2BQvm4zw7GUzFH/CfrOQvBGaX6TL/bekAaV70db9mOpP8CXNBw+CcNLlS9VMscbJ3
5qItw31/6+hbNC680wh6gR8evAKmgAgXb0rNPX9IhnMvtbwrzhoqEVZ+T/rrCR18V9kMcqDe5FO5
9aAh1VjgDaXlFcDpvHwVE4WHMxHqvhTWy3CG15e9qEPm4EtsG+yMsrDfGDLU3E973reZSskIg2f+
KSCN5hKCyfQibJupO3BnvAX1G1t9/2YJGp9wJaoD8OdP4Y8qVqmR2XK9+JJLmgZfJ8E+mLmUWANv
RrrmXWHmr4RwtZkUak6+5tuaswhAP7w3Mrh91mo0wlLscpuoAE/MgSLuz6x+8TRAtUon46IYTD88
HFFJyotSz3tv064Noq9BtkJkEqS7+qYl9In6YQh5NotQWRt7c2MJYCJPkMPYxlMQVFai7P7gH1s9
XbjCrn3ES3wDNPydchXoR0LvWgN2eOvlCUy9P3URbMx2ndwO0PjV2KJr9dGz2jLGJyhn9yceZiGr
IQegRxvfPfIdjV7IxNZSU2qViFMUmyJoKOOhjbbXIsmvIgxJ2X7B2rKkEpxLGUvxvYjwqukp4cHN
c+AsPYs0bfPxNH0SpIP4jrRmxRfaC83VbLFNb7LcHo0Qde7XvX35gGjmRdz+GAmxqsg8zBlaMmzz
b13yfCZE0e1lGnrkH8+QBkMB33iepAaD/3DtImSziw9zKEDEbYFlEuf36l98+HtEr+JS8gH8wdDp
6d5A4BKCshvEKtVok1endUOhXclwcexWGgiAm/mr0MxecMcnULw2qV4FM3/veMxcoi7vpz4B9vgy
ox0DQA9ayvXGoZ+uQ3SH20O87s/tZ8odREF1CoOIOuDepU6jiP0i/558QR7kg8OH2rNufw5bRDXe
lKLAO8D9ytBCOUgaDbG0qzBvCew/klVkeqjhDTmRcgU7mK0ip8+o712U1A4aKWBBlutGjqV5Zh2I
UBiobZ33N+C/EyaVng5jjoJe1KHdfgtkgeGx02x37rmvGwFcqBWhrsZPtr9MB4BRkcOy+gz/WtoE
RPAiOgXY/KYFoQc5c536rYM9Xi8BFh9896zsdTLsjizAREpK646exYwCMjsHwmdLDspsg0aiakbh
+sguZhFSy5R5SZtHQO2kbiMtew6ZvjkgFrc9MIdMjXWcCu6TiJW67FasIPD10DmQgiY6CM/lwzs6
8mEgJeguDI9OHC4AjhXmePiv6MKWkgtwhD29qQ0Z8d9Nq8Euc/Z/sqmrbSUqQoXKdog3qgwxasxy
Qay6rAkAmaJlwlo3mI2eDzUs4C9dWY+XPn1Rqb0nCaMiFMqt3vOG7ylH/IhuF0lXhtLv34vcFmg2
OpVqXqXjfIYGO6OyIFsTWmXOxxw1nplgb68Y5oM42dbxnTcHLekdl0VpuGNdTaK5IYG4GU+8on+a
YXbvcY0cyjY4PGSpC/lYukigZWQBfF/Zo1nZXkBPYVa6jt8O5NQhWwLvnNgzfhEUYp/VwUcvZmvC
UgMilU6dqsoZuluU0CtZ8QeEzNuZkBwMJaoIXcynfBY8/uvcLDrRcHxUZeBqaK7/axZr8kmm56Kh
z8GenjZ7lnz2TSYUk/Vq/BG+eflu9/lhXpEQEOqZuhaWqWTVxGjWCqU1+mGYXuBfUb2etZy0BhHT
XwN8IWfhninI/WtyXAixfqsuf8SXuQOrmxhkaYx45ZvsIPmddQXV+ihGrtmcqQJ02dq4zXa3g7iB
SdQh7IumVJm2MynvIu9S/A34s7YpODExM3gwF45DZXY253yd/d57ZW4HPddKAKUYf9g56Tlwd5Kx
W7aLb7Bwiduw+uJKeL3sq00pZ7OEo07RsbGClOqV4H+uleWAfGy9svD4xYZ6u8S1bfCjWiZCbNee
+50kagvEf7utYXehFt5J5aD1BDzmyhRJrPkb+SIECWZDEl6K277bAUlpZ4G7BY92u9FRD/jbejck
yq+zoLsSJntn2YJGei3sLTFBvjfeNHSk9MOC+c6CGcisBc1+lmyRqlAMq+0FYXGJkPGdNQbza+KW
0HZOjCcJURHO0WixGVrmrtayz36tMRzNaDXj/VDT1+IRhT/WGc7Qmnkc7OzmIft3on/R+q4vgbRg
L246RQvKNXWV2uSNLt+VKdGp/f3bPMV5VwX89A9JPW+HJHPE1Mba5IlumHiRp4KLKUu4gtwk5nej
CldiSrrP2EugVFSyMVYcgRap7SPrhe6ahjtrv+0E8iC+GsPN0g97RSB7oAF2ffsLr3qiKrcYiwyF
c2K0dBsXqLTLzK3msqlFP2mcjwanHUIhIRTjN+tu2G/HJFTU5siKYcz7ANGIVALWBCyncQrDdlWf
KwnREJI2GemM6Io/NHoCg/Cb0K1m7hR2kWt69Dnxs2ZY/fkFUdQWCunJoySWrATe87Z+GMHICKQH
ZbdfyZ09gjApZ2wASO/Y1qOKJmubvNsgscwllTrMp7VKKbDw6MUYGgOo9DnTxwonqwZZuEAo0D1B
/JgD/H2oNOeXC4CJfEdgBdbUO3GVE+wJrSw5duPe8nDUAl9ESBhikECMTgoRUqeN3NiGKDRNYgQF
8fNrFBopdHb2C6cBZML5hEASy/IBvUU2JvuWcr8uLUboPShPgFMMVvIXC4DDKV54rMzKoNIHDstH
oB3w9WOx+y0mnR46rNkuphVltnQZL8GZK+ynla/vx7SZM919VrO1VQHhkEyHqOdK+JpdLMDYTl52
nc/g4BxQC8rj9g7xzx8Gu3kjWNEpFs62lQPPil3Khn1HdxLpmNCRh396DGjbyVCUbouFha7u6edn
BH20fgwnFarkdLuS7x/OrFSc47MN1LgzkhjtfLLNnBhDJO2X2MvPFP4qB3EeKW8rv/qWWKJDUx3W
ICr4kLtOkX1jgm+mrlORQXFdjLUZcoIbanI3QzwXxP+COGTn9CQ1sDvKpuI+JckAJIldDFGEe7ld
WWHb/LnQykJMUo+8CpTJ+tTMOaRBORxe1Pec6kgUSOy91DjATCAC/oaDCnBHYWQMFTmY2/ROxhGb
fwWXvInxT9Ih843ojFlUBEQfdA8anmZKmFqiBCsvEzUv/xvT/NVoi1BxYDVoQiwyjEq70ffUsxhX
+39D9WQleuWybFQ0jJn7/KOisjbe3jhcq/Y7vMtyvqF6N/yWx3CUIv2hhG+25btS+Z9hc5ISyGGl
Jes2xslxfaTVEbdxuJkh4x/SVZLA1XkgJ9iZme+RFLkItnUgdGrQE6xDkeQ2JKCgA0mg50CyivS2
K2dGOoYswv0HGlOpK7sXbW+eZ9sadUOxQO50DjXbJLPZWq+0lDI5Bg+JQqy5seFoDrE9RfB5f6px
1pYJS+BP4A/yRQfRm5OcwzJ/39arx9BXUCAqJ/c9VKgTQP0aLDebcp27Q2b6XH9omWdl+Y5VXxT4
k8AtpFN7km29l9FU9LzFdMmtkZDwJUmKKrAn9v/jyjfF/yu43mHohM1MUHGV45Y9D5u/hS9VhZf4
61y/N99zIQqqyx1gl//jV9APgtDzKuS7zcRNsDxm1NnSh0b/5qMHP+6DL4taAFMUXVMquNUp6bdx
xXEgj1k80CSXLZJvouWyXnWojE8x6zdzzq1cwvQxXtvJUrdCE+A9yfdJnPugyraOaMsgpeO3DTMb
S5zcXGXwajIIG5GYZTZCP0ayg3Xrl9H9OutBAmbDiJO6pG6nnauJ28b/H8DwIHKMg59OX7TaI+FO
kBUXTW5Zq5uXPDGy8DwMhMpkxg9o8huLjTF/YYFVQFEW8P0s1ewj8lHzbNwKl0UaW8mkr+IciGUi
PyKIteh5zx958oFNvIXRAVyYYdP0w37E5LIEQ6IzKLdb9Qk+HJ9rgNz431UNIXe5u2l4et2MlEzz
OWMjKBmQdBmknKv69IVS4Wd7fbzk4Bb8Aqf/2WzeYAySeJq+/typOE9jnnVT4Vb6Rd90aRGyfk4J
uyIqre54FASLf63i5dam74bYCUBrX2rV6qxZxcCpQSpvA9UoFRAPt7XZJuB3IbIu05e0CIT3RvX4
sYaW4CjNDS0lpYj6SdMIJNAyrcQsi+vyIzliSOk07mC4O+cYSfcbRWck+f+s9STpa5xc3iUilciL
RIn3JjSivDekRYX+yMnGNipekA85OJ/Wx0bON3beAHCgwX9aZ+a4GsTrR/So5tNARc7Eg2zQubr8
dHf7jcVZGv64v/8kA6ccby1y0hrXSnyYdHwZg0Av3cbojN+/WZfZoYD13g3d1PDNShYbyO7xI0ad
gsdws/3lHMb8L4tV7Yyt6jfbOoLw7P9dqVivVbn6qjGWo5+RfOgy7TRWwxpFrncbH8e4yZzuy9ln
8q2EjRvvKyw4gYIPN5RBqyUDrHZWN+emQtO45SMewz5uRz3naX39Tv9Uk2G28YRY0gg1DVGnIXYz
Epd8ykzbQ9tLo1DQM6GBXih6HxU0kPss8H30PWNSrEuKWFq99+rFN5tC4zSjeGvkYDJ6wyNllK9Y
Fv/nVFPzSWJGQMuXsL1N1FWjML4R8SUyUHpoBwdjHxVoT4X4lpe7kbDVgK2HMSlv6LYa9HuQAv5M
zaLDNRPHlz2/Y205K65HX81YM3CVmXxOys+UrbRHK6Cfe9ldD0+HzqSxVPlwVgg6m/jz9B/29TGG
06DJdmcjq3lrTUTtLj53Hr8HhNLxjmDVOGOhDWabOhozZGZkg5pWXyBW9tF6sMIt7wxwPmOS5mK1
3uzQ7l9yTQVxNgO1JukTAd+JwBynDvFAutE9MuFX/BOi4pm1ORXfte88PVltElU68QF2Z8uvVoXd
nbntZmCG91U6aUCbHjdrF0AumLTnL9tLTrrCMH1P9YE/+EGpefO3zbQ+xmcATbttjR8iKpMtSm0E
sDjczmCaZqMY2k0WKmLRz5CpW+ox2LXeIFPtTUaSvDRC8KqIpmQjnA/uhRUJVQ2a93ZC8MIswVQE
j4U9STnP3VUjsDUzsopE7sEClaWXm+vU0X3KeOXc6xCQj8NvVu8IDuh7lp1XTun7ziYXQBczd7kN
lvjU7Ug8JR5QCuDgalVmmi7KlKpo1IwWVVTfNHixfy4xrbUl2IVmc3AzQHW+93M6gr7mTdDpae2P
YaDTTkod0saVmP18gHvB1+/quvkuczPeYm8d5BxGe5LuB4BojXa4S0dF/N3x6dPJal0Jxw+acqVW
wQWwcqW89KgvU6gPMoN30HFlb2iCabmN7NpSlMuZK/dErN2cKz6WCcjavH2E1fC6JqoknURPRPl2
kw4sC8rd1OTmOLIV6QUkkpOoww74+2a3SwUTjZ2aOlM3ljT67BDYkvrYbt6HtbpK+BPI4iTmCbNT
u9xDZFaOIsKMb0tMTaEJkxFIhS6QKzQ1nHGKerz/ZSFthQV7YKbQdyd+DExuZooYYY6m5gRpT7zM
PI5rzdkJ+AtW8MKSmPhxAszVNpmLl0t2i/ArUwdzYX0aGDvLKkf5S6ThJzMsJada7Ip757p1IspH
sYxhktOuPMtsE5lbG1nVWuPIj5F5iiSculrineCAiVL6zrUNHx/pT+3Bd2FU81AQ7OaigYw2UTPU
OSBYiNNBpzosx4LfWoWOVVx+aq46lE4HLl3unwWvNdlALWDGAcI1qsPJOUhinoIYMjhkUbCK+ELb
6u9wOokpdnVc31WA5k/XFaF2cWfcFGaVVdON+OxqQua6dR+fBB4yYtb9kdMCmhKLkESAPzBhrS/I
NIZujNuBPoZTLlqOTEt785KIA0cJA/3SO5MWEX1HqUKWEvb4434aA6z4Y/RfY7eGLZVLYKvgjdOZ
3J5zthbUXh85MW5t3ppyzM4O20C42RAuSBBMBPufQcJycwNNlKJdwtwGvFL45hwOZHb3I6iM+Iv8
C/D58dC5ERBpiiX5xKMEO0nDVy5AvpE2TO/r69qzQXdOwMrGJ4/ZPhPULgy//nI7E1QXdxgUWLmi
WjiOxF2TPbtusuo0h6nQVFOSRHxdUCyUQHn4vrl9SbyYkDU0sOIq4HwdxlDf88xicRCvu42wNaLX
eNDyvT/2cSnctKDjhDYR1SHvrwkt9iCRyzvs8phvcr1RlAFvRzu8VjagVuJAcHzUhoVEuC5s8Ct+
jPn1L2TQ5RMDN/8ZGIIv5Y3ZEIPHmhLohgIlo8bZt9EV3FTcFHS3WC1/Sr2yAh79XKw+GxmEtIkE
72OvCtxi+scJpPWGq2LHpVuNUv2jtns5wk505mp2/IMnEB1gYhSV2OQTwFNFmCTbbGeUnNGOA+U8
4WhAQ+srCIVMsWMlYbUM+/3EtW2CWLGaI5mMSZ0/A9GqKuusAkJjF4IEavf45wE3Gz5OpIDgFN9V
1jwNHT3kDa5C54kX+xefBCvB5sNx6HPwuGGIf8LXkYS6CZqGuni9jUq/K/7XweX99BIZ2rIt25Av
7bUY1coXXQXCiekhh6NlMNtYxTzh/8x4Z8dekY/D8PUNgZ8Xmq6MmBJE/HXhYWn5QURLUE/fI9XH
IICysWj2wdGZMtvE33QuwcRl05Flgahd0v1ASYM+9OIOCPUIS4KWYq6Ii39Lb1Up04UZzHWPCZ2l
mWY4mxPKofp7pcUGUTgjeC3z+0FmEPvJMezqb4YH6y+h+WCYUptHYDYtm2rFCcV6/PwmJXAIzsk7
fc7+epV6jGV0CQGns1fVZoeSJjD6PA/wIjMlXzbCl9vm6nhiJSudCMFcSfxZfL2DT+AnkxIBR8Yt
69P0ZfJwb9JlwTm6zKZdvJiHAHqsw91JGpjRgj3hHKMQyO3HAB7yjqvJlWXF/s2pQJRWtWvE3JZi
hFJzeveMEyEnd1bolCISfeyzciYw7I5qv8RloQRF3/IsPZvaeMuuG7fwSUd123sStamskwkBCQ45
BKTd5qK6Yl8HjZXPmzEB6OshEsDfhKNOwdBjk4uNHEWnwPn7i1Hj9I8YqxiE+KbBSL5N9A8o+klV
zeJO4QBoibUAEr6dfLuXOZCbBrXuJQo0TFc1hYqnVQja65eWuN7aDSSxCgP3V9rkreR/4L6HS0YX
ktFnqc5J38xOVvydguo4DGqQGhTFYVkDjcloCSg2mJS3XBWL/gE7p2Hfvc5Ii6EmzY/RwdRycZ3q
lx53vDJp76hGgTKtMO/8XM/EprSB610XHh986Too6G7uoeE73oMZAX4wcCh0qIDRIiAmg7J9GKPX
En2m0a7+H0nZ0kgLyjk2uMHpwMgfbmQ7/8LMIyM/H2MlA7MsK+VlGdYnwxU1V6Lk6yNQGtMTnIyM
ZYH339CH3Dp1wvjrghoOqX5kvU/Mz1ZRVIQo7v/0PFoOzGDKHy9Swn9lVpncFEryJSOaAOQIU2AJ
QbOIwhDES/PxEPOYQ8mhQcxqMmp7l97sTTYbQfWrtccUq0FgwI4CohYE4Ok2z6RUl7aA4wuAUi8/
zQDFk9TmL3nyVvWR1p+6ahU11qga+3kDnRCkQdus4DfnDhYvK1RXE80iKna2ejhUdcgvzYvO1Car
X65CnIS5OviJdTux9gyTPYmlhTX2UYG/8tND5Ia4Scsz1VsgZ6YvkFmlsT66yFrs6lcGxJZ3yY5X
+bgJNrxDY8r2ifID5FuLiOKI7KoedN02PpRYtCf4LEAJkJH+oL3FNRKLG4DTC1dUdEkGmAKsIMvG
5TIcZGvpH9HBXpO3gs65oW2xOo0BtImmWBVpRmLvM0oTvYY8l23p+yuzwmAW6UscJ9CkqFQl2H7y
l4HDE7OrOZfJ+T/ZyZkMPqw22ZD6sk68hPb6p8EHmtZbkkYO72X6KaUgLau/GL10/x0iLuWk2eg8
fJbR+LsbpRoVS6mW7KN8g5LpIlhYPgJr+fTyudDH/B+cPUZwqa0KS7to3W4e6wgfetqVX2BPhLGd
220u+HPAtqABrCBmo7za8/eqPJef6WCPKj472sQOpWDpltZ1Uoh2HFkfnUP4c6c/oAfWmu2tZr2q
fQJo7541s3QqNr6E81rrhujHl3P1qm0eo+tAoVGG3B/oDEVO5e2VT3Luypm4DxuNmsGBdC53xBt5
CCxj6a1UOYsgqOzaZ6FZ7kcs3KdLMt7aKNvLaw6MNHvqvjDAm2xdWXP2SioznJKaVKvwzUetB+Ip
XuvnOviWqOnKcZbTo1/8UzftThLSAFVTudA3MQIqyrcWVZV5bahx8PfUetKsShrdK6gZeoL92weQ
385JQu5tjHykngeVShA4Pq9XdRkYpsglOWZBzK2YrymINkAPnZDJq4NVNT0YN+TKXF9ijd0yfOJj
t8dN/KN/dzQrb2YymthJBUtYidiwvkzRtJG3kNocgPIgVNzrfuQqApLVPJTp9V8LeDrSlIAg2Do6
oW6zeywuTJGk1D5l3ZffEgj3sBlc/iQ9C/pYvI8Ndm7Oce95XYuTjT+TJJK5SiCKJsAGLlW4lwIg
j7xzDA3kWwqY6OJ4k0XXmeHnkSKgOMKvMswKTxLXY33912Z4ieg8i/wP44kvZfMX8jhQdOOM8RJy
t6ee9A1leYBfg3MMwz3hyFWS1yInpombhDDi5i2UsI4pY9FZp4h34nmy68+f+BK3Gli7gBZ36LNw
2hS6VOy9FHsuedSwKBJT07T77UbWreS78u4FCW3GgjT69lAstGO4GQNIqy1QaHNQcYyiTYZY1/uD
f/QR3p6WbKxfDKO6EOO0T57CSZ3HV3c5PCmfq7yjxvrLkVY1ScOr85YkoD14HjDg5TRXuZm8408E
fARoTYnVnVjP9GiIChbJ8hprKEXbWS0AY0Zg/vyMQrsSBSIWMREaS75dMA4+Vv8pEnGT5W1xVic8
NHAdTT00UlQ630mwEFwOj7tPGVBAvT3mi1+myGB1vdxtpxc0lVdVlZfNFq66LoRubDwNFw5b45uz
gjlFX/rxV8AQ4P/JsEwDh1eeijcr+Md42o+Xp5Y/9ruPZut00s+yIYUqJgiB5bYjGx8DMbr1pAF6
nxgwHiKP6d1TA6FlxlTFMGluYjVWbJ+3idwh3Jlq+NNzq6ZARVMtZHu4Pm1tEsB/9rBqLgSroVIu
4rBpTr3lxKDhPu963i3vGET1yIzONi4D6ZBqY3C0sCNSCUicQLFNvEJoWu1g6F/36Y2uAYUGnrdg
zMciE10Qf1tlsl1/2LUZV9we2n9Y4LVJB1+nA1gOAQfSwdKDhwEZnpaeEm3k6YiEcB0jX2AECbDS
dHONh4eWeA/gYdfT0qDhBOxnlSuJcJYI4ivZMkhlfi8veSdOlFdp+drFSHif1IvbMTBcqzbfVb81
cHhp/SomFP79DSH0AXqag9SxaUMBaJTM3Xv48FdwzuX4IbUtEWnHSlRxIXKwIy+SOIz3khsHSUwT
Ctv3OqsZumdjitSFWVJlsCvPkiY3TDEvl214BD1ZNkjMPyuiT2RTFuRofLIb9yw0u4Jfq5SJy5+9
o0mykZ2cIbc1P5RMF/0gaCpWRUweTYQvufcJzHSOrmJL+EtExdQZKbGsP/a8ndHonbUjrVj+xDkj
qQN+PhKDwLuql5Eh5ayXJxU9GVOB5oTSsbs1sRqIZi1BkJGs6/b3uenBXDOM4FS779gMsCfMGZ1X
6csnACjkbL5zOZB3ydvYZ5N7wrYCC6z/86MdMMR9DjbdagkQ24byU9PLnNptAXpQUm3AUE83E6FQ
7XV00zOxDhsyhos210wNUy9Y1GExcsUqS5rUKvbkcDKwaZVE7d2Z6B1VqQAALoa/FG2s2w3I6Pin
wGLbWF/acsCrskSaKcpmo/q9DZAaTcc23JtEWTVblTILk/uWjQDF+aGJ7clrQtLmM3VXYF6PdFWl
i/UStE0AbAFoiskAZxV8lgq9v8EBCMziaoYNgEp1sGDGnHKc3Q4hm2Cp9WsMXu/XbOyFBeDcsizF
ojeNGPhvHWVonhl/omqHEuFG9H0min5ty3xvKdOTRcYKciOd03b8C6wbaa4zHJ+i8lHdDklweBbC
L/UY+ki+h5L7QOSk9H14ZdXgUeVAydC6K+UY+oL/PjQt2bBOLJtSGKi4L35Gi/2ahBxfCzWLaVfq
wMnKiim0451wFf9EYDdQhQ1AnUJklU2tklnYz8U20xvFHhPfBDJqeKoJ8q8Jb7SO7IIOvNPw9AF+
VZatkudUA+IWaP0eLUotzvqIMoCuksrU6uoKRPXCCjnX7V7DOq3LXps0eHu5D8UjrvVNGXSiyy+f
a5kNwCiSDB5v2PsWgOrFXcv7k+wOwfyPZ/OZ5YzKXxX78qF0Gva7lmo0+CjVJVPx1tzYkjR7OqKi
zyz5zVk+cwKz44umKwneBdaYSg07cY/u5TtgwPAk2t3iHgEbE+lxzNEqY49p9aad3UEzxJgZ1FE5
dsrwOWjjdCRuj4p7yc2XRXztNE0CX0A5u4iwkEp5sxzU7AJEcv8UsZWDQEMuyvQ8XruVSNpfwSwJ
6areWgoBofSQFwqCR2sypeBGlzHd0Jtwy9vQSpCZ3RLbjQ38tgRSJHxbHmwtImT7Tq3mVYyOlyBI
PKs/3IVIK1YowIxXZsnBhq+RKXZF39OeavEMFUyj2mxb9tXT1IEuRl2prNIuDgppPt4jCuy+vskd
M3CUECCWSR7H1WQwfe0GfjB2I5uW3hVJl4E9bM46npF0zWnJSnfmhu+5OXXueHOcIhEaNtrqRjj5
8guJA2qL3lMLJtwlQpPSxeg0sWM3VWjzCITUGASX5tdjtmux6K18nUWjKLfzyVhShWbrGQuy90OA
g2oHibk+MwxiNMkOKoi8Q5Q/+1R/gaaz+FaSS58s0rVed6kDaKx94Huf19pgx37Jxmpfl/7I4diV
Haonu2GrnsorYMRoaswxVBMu6u7EWnNYQXPArqXoLHo4vkOO2yqWHDQ5XCL1d84XFKZ/Dpb9JQkp
VEXCLYkcJ2296PbAYs+qhlIueOsUzu/ZLQNejqSCWwrtwpIx+rR25B/SGeZp/pnbIT/lq7JEXU/j
JRhnTta3Rs9ds/q6sspHMNHaajOToHeoDV5ElfohdWFREUMA6sbH8KseTU91fXkd8haQ7ULv/RYG
E6BMNH662SkTCVF+S3rMOn+oO2SzIz55aS5wAoQBojZto8lVIZBdX61W/rMHaCSnDMRvk2y369fW
5WNZLi7CGFKuMFrXER1U250L5JeLeVLPb3KTL+dZDI7lxMOoPIwbABxInFFktYFiAQM4Rm4dejAy
+C3rMiVJaRRRjTwlooZnXNw0sqiw48v7sMeDwTfnu9BhXUS8RqhopueVTsdanl7eUixOhr1VbNG4
FQT3GHoPeTq0IjGD9Wofzqj3/5wqdtrUS9YSwf2YOnTPNawN8GdzeIxbaeETxiGzfVwohn+eUZlt
fmKIFLbnsxl2RV3HDQD0V9h2iYmYTR5q8jJD4lfsCbZAt1PNFo3OYrnhNAZTmDK7JJHsVZgVbDu+
owwIuLzqBWXjqccA+RuUl4Fw2WzRA7gBRVx4/eyGM8UdaXTbO9v1TMOxagWkKdAK8+NfPGZIyhwZ
NAhGaNcpqvIS/vap7o6QE/hLzxo8iF4hBsKqrG9nBew14rnm0ZFf0UQRViTvjR5CTNSu+0TmoL93
5YdSW0vubWjHNsjhzoJcnNA7IaRa0J4/7p8SrLw9qRXWuTYS/IWy1gWJhbIQufEfxzvmusZaSiQj
pkImX53tjDaivM0f0yr8d7XKID8o+uBC4012SmwpwnicLDpfR92cMdr9RG7uyrFtaUpia8yMCRXp
nRYiRnGcZ+yXB1qNSlk4mqE44+vR2DqEnubi0vCeBIRWLMbdxf5TOOpjY8afslFlMR+RpSZ+iSUy
+ex3XkJ8N3cktD7ruocbcrAGDOR7jEGZKxNC9dO9uYGoODavvTGLUQXJHV6MqRJWZCVv681pnHSS
/bpiy+HeQ6RfkOWZY2MDU44PpFwT25r5TDKYINEBOMEDOgFEs2rsShSxJ5WQNXgVpVFI0OHQLnZl
OAw9wVcRxCDKoXZaKdwc3DadPzXoVP0jvRgxy0zaY+c3gxj+hUcCH7hd+q71kLyEpAcVeACh0BRv
6qcDybxdU3JZjG8CUmQQaPBEH87YO2bcCF7N+ULCCTF3FC9FGtQm/mhJHSQIAmXf5h+4uKgY+GqL
tAtVcg2cxbQOqkcFUKs6pdixGHjJLSTI3xRr20PpPlZQjxQCRX0i0TIst9t/2K8b8kPiPvJKX1ak
Z8qZTYL+HcZAuI2Ckfez9PNOFRXru559IhQYnOZbff5ZgWTObER3u/L+npLW2ktuhia7S8x+WfD2
runit2JPNxH5xvznZxCE7qt56halrp249mT3Tkhy+K9ObzYBUBmoOIpJOUwCaACsXtGKHdjs247d
Zd8MpBXmD4NNwXcd6vQY1oq7SbUiZ9dMNwGW2jQRCHevlTN3iNN3FJJzhL3xS8zlgW2y9QDmaS2x
xT9kGtdUAje0E2pjQJIf4QEB/ln/eXlgdtAB7zJn+1YYRVcvGKtOwXHsFx1+TvmJF3Qi1hu1Cal+
HqVbc8Vl+hfJ9utFQboIhuUw3k3FN/1l4XHMcbGNsohDmjr6t16pb8Qx1bkBSNEeE7IezA0P8TF/
tulQthtP2WsEWIs/TEyYE6TMhrHqxTKKAjCjHt3aQbYv65AHDEnw8dAq7kWzbDuAEwqDY8FZ+72V
QDtjHxOskWi3sJ3/M0ZrvRxVPrSscrzcBVNlJuE5CSOma0f6j6Af9tCbnWZb4rsQ/JDDsMZjrquK
rrHgUskmjS5IrPzVhzGGOZHsJvihT6nZjcO7x6VrfTEKTS+VQZKg6nudEOhd93l9kymGhf0O4rRh
lvUgF2nr1Rh8hFolycjUTv1zXXZG84nQ17QYWKrrl3IWCEqxcy0oYzAOJb34tNPd0VuXgei6f3Op
cGid4EpT1ZPOPz9c8gBfw6k0W3aVXEwwG6N2oBrvROHUWun0hur2yrvi1Gmm37O80mJO9VlFd+9o
WX20reRy4MipAKbnvhhmWYw2UW2Ue9vnrXWp1sAdvarkm8WJmt9irt4ExgxO036BVFE4PUK94v0P
3URCgazlbqMf2B/CVU1z9u8FaXUQhRnqZFDhpjJj3txhNf7SOK1e+4p3p3iAyzTIauu0pZ1elfjq
DE0k++PmFWpAD8WaMAXjkijpVXwrL3BKoggpKco72/lZlL1h/JElMixol+c66fgpytSo7EUhqHmI
MkcwaGKKs+SFEt8NusV+v3e5qWSMw1AWiXe5lvp3zb68F5CxTYJSXJTHdzyl8jL8viRR/5pXbHJ2
y2XDYVL6QVTMo7YYqyK2xlOfoo93JeHDiWmLlNliarGH4jFb4C0yjUk1OSGRoO2kqxcKDMK8r0h3
Pv8OQlEo44C8yBtyDZ11YNQvhFEyNjFiq73KnFp3cVdb5+s89ddLNDbwss1S9JvsA9v+dRaKBjNm
IXxY0NyZKaXOTJz++Twad3rUGOS9TV4RvhcR12uEUNYEvChO6eSTDdpl3h30ZjMELzj4yO7nt8S2
GYeyQGE6/WGgCUfnwmsYfEcJXU39ntPFO5WeQuztTXhMyYF/1GSXlbQhPGPP7JNsbC5/it6sQ/ws
zTSP0uLJt4ZVsClggqDtbfWPK0I9XReRxlFAhYmgZRFsmF9ZjesBOFQkhH2Jk+5ne15t/+5Ygos5
RduFW75MSj8u+fnENcIemb6edhjJjKjvVw1NmROTBncF8fFgcEUx1yOM5tukk3v8Rh29JPVV7Vrw
Sjyd0fnNeCnjH4h26zZL6y1x6gWJ5DmHzK5IMIZTybjn52udCKUlOnqvsXtfp5gHZwegc85QiDX3
hH0nGdMXJqmtAU0nxS5hRSYsrTokbbYilONQbJPlfgKS9T9n/gQEjmK2mAZhe7bu+IVR1p4MOwGr
M/TZ6xwD4HCpqKHITeQiwAKg/lt7kN6ebI9cU+WCcTcYdzHZWXEYW2qL9iDA9y1AyIKECsTmwhnn
pSHzILP+T5ll+0C29u3GfTxW54ZTzdYTyg9bXIpc8ew4/jm3AZUOZkoHLMaR1k43cWF2Y13eFVdL
fFGajIvMZp2F+rcHdMd8yTnxbhwkvEKA7RPgheT2dvjGPsv62QPXbo8ERxI0a+q5kT+9iGzFVlva
j5zFB33T0I2HTmhryahEEFU/lb1puBtH3RShSLLT8YNQdgg66n2epCz7xG+S0flcTzzyDhNwTWei
OHutTHfTcm8N/3lzWbwRsEnG9bKsXQW1fec1XcAAp4NQAiuD3WxHIRA0X8PyedB/QEIJaoIozPQf
wQAbKe18GerLlv7Qx8BhRWDcmHidEq09Kcoh2aKHdewk3pPTzMsoz7fCvMXlf69TDpgMUW6EAtcP
E3ZR0ay1vqG+aH3iQJq+vfJD4xpJFBymo6KT68ruRwYe4XUpiNKat7Vc1LuyDXYqZJym+QGzAtJY
B9CZdRPOTUgamJK0AL+H4KZXOwv3SMlqKD5H2BnTOI51G2z5w7CGc8FT+ykKURFjI8e+Qd/pF+Td
w/bUpkIksx7fbWkzAYJXypKIA4jcvA9/ykECw5cJdqrx4c4gE1m6w7UlTO2KThDp+5l4VH84B8qR
QfiL5TMQDQ8C+wOvVKO3f5jx5eUnH8vqz5egR/xaBfrEFUehmnxmOWrf3DYSYE6GKlwIyipK3OP1
KrNufgItvRlz7EoxwURbF9FegsGx3KCnaAkKCv1LVw8f3Z2BbVc9FjF1Xf12EEdndakILSH0WYEh
FjFCLzrOKZyP425IAfoxogPEAxTON7MrvQkbVpLyUodyveqMSt+E31ft852ktXEXppYfZwjVRs2V
tGk9GBfCOk7RqZfgT+fLMB8zNbE8ywFBmxwoiE3uYIVPmkacQlSrvLQapzsLTaTqzcI7Y9pzs86v
lCp05dnR6cq+zUxn1lL2Ctzc5YN+clg0K84j5derkoCnDiWnLzUAP4FwrySG4AKDZRLVBOcunP+v
AkWgDt2NfN0tdBkbuh2UhP56VtuwGaqngeAohodz3v2Ff3pDNFcUv3DiYA4KU7p2XAeoLxc5bEq6
cjD0pfy6c5QG9RluleooOy6XoMVN27IlRz8AbuBjYuoxkxUKtzg+v4uOnarpgf2F3aXElTz+8E86
UAB/mmaTfB0zQkHOX+RDNnfalH8UxFnSyUS79MSIoNiv5vvkexunmES7D2Be3r35J0drmBrBWDf4
SBj35P1f7YpV7cYoHXQYw8DMe7M9KJ95BTqAHOd0sAGzFliUF02YYDu6EambDtHuNO7mLe6Aa2K3
5mKrig58fCFlm1ySyQ7FPOoT6969bxHi4wdmp4WXOb2fDUF3wA55f5mVM7xWoifveigClJLsP1Xj
vufNZlGIi9fMM8Na3qBlnBIekGuKDEoZpgTncOnnGRrBJHL2q4+EFPHx5233uaZZhWUnyVgHJgRT
EEsXUDjdyajm+jeN/wcZb9bGMzbVORzA9JwzXKvg2V8tn7up/zRr49WdsqVBPi9d9wnb52PTXDQb
rMkTKyDxwZR5847ranl3NCBA2D5eqCNOHGW1u2pQA7AM7jhQHf4rVqnKD6F9Ar4WzjSMAPixM17r
mYM1hHy1MT3eSe0cwBHTFfe+7I505o30bjc0N67KCCQQhM/BhVJG1IMnc8RVXriyky9DddeWokjc
ew0eBvlQl6pwGeHNH/x4NraCOqMHFQrKgiDMMJvQ80yIFHErcLdIjEtCwb8+FP9X2x9DXZFI3/qH
r2Vhq31vN9g0Tk8DHna4I2dQt2t5kzf2el3zg0xCWuPAyHIdo+gWXFNxmgec179g0Otc/zN+DoZN
Inv1heu9Z9rvlT5pLjQ/DZPyH51GGxNEbOWU4TYNa/AdPK0lH+O92MFPJ6VpnqTSfff3qVIl7TYa
3ceH9FwbbRwS6VmiDCkVFvXa026w9cLx7uivVb/KjjLZGjPn2Y4aiyBybFL1mope7YfmvQuo5PUL
9vlEcY7/IZWEbetDVpgUKQtPDjYWTyrM1zusMpV8EQCrrInsR88FFyC0Tdk5MV9VOorOlZ66M5Te
k/t1Mw2IOsykleSUQ3AXeoPnZhDluJt1XgtQcNic8JmyUyyS0o5wlSIUfW40j41hkB5qDGzOZyYY
IqRkeBgdJONW+k/jwg6rNePdu0kuoq6Y36WDZjv2hTIfj4K44zPDFnwr8KjMxKGGvuVO6nFwZfpZ
xoxMsVn00i8k8Y3PvPSINIL51LDoBeTyVbhZr5iDel5mXJ1Qa6DPFCGkl1XlY1YJt0tapfSFDPh/
zTRKgK/e6Op3KbPr0kzbhTVoTW2nND9Img8uGMI7E2iFdL/V82HRajwbXh23AhJOf2ck27vTrBEt
UJBMGxd9+v4+g01bK6hsmiI51rlJAla3Q2dK31DGFpXqBsa3MiXZHmlMlRnwVjhpXIZsExUakUW1
Bxvh6iLBRW3zQhVTzFM9C706qFuD+T/22yWVhIMeRdEwZ1lPYrYGIGolR+TyKuFXNt5KgUYjZ2AT
G8zhPXbZ/dRNUzTuGszAgVXp9UQ+wSQ3MTNQpsc69NWvdxibuWbCSYG1BcNJDxMZ7PtH/XQ6OaTk
CAvVQSpvFFEjLZAfqrLZy1L3lkwlVgW22Slx3jeYpmulWnTEOcM0fJZ5X5DFK0KsCrQ1ica00Ob+
MLefsb+Ws6xydcoZ3v4Q6SKUF5c9VcUrBv5ANO0BsS4/LJFuJT1rp7uMkB0rmT32BMoprWRW6Wrx
QhEtg8djPu5R8nvHgkULl13koGlqQVXLB5CcHuFw0bbsaeFteu0McEgh2Y34kE9BMD+AkVL0F3Gz
bJzBtnQzc+tsERDopdLlo1JcC4C9DEjAzSwWCCYWQJcXApFr8bmT5BwL9agCVkflxU1PXAqVsN0a
+eK5Oy0Ex/HzqULf7tTN9Jz5CsGXh4Hwz9zd54fcNImgK8GlU5xQbVZzyuK3xRF5FHAu5VCinVO/
2aDY19l+4mwhFrTtb7YMJaK3b7b0u63PYZEcmWCkdlU+BI77IcjBWDYKaKQNz/UXSAcQZyzkLYUj
brkgIAAMsrQ881dbJTYTQMESQgfvEoIY/8PI5OXO0nZANcMLegspOh7J4q7gTbY07/4Z5Vb7cCOB
C2aIxWuH09hYiDv4D6Bxm2bzVFaL/M23dSkszP3ikX0WYqXFISiKJjdklqU5fSr+5EDMTg2aW5UC
ZXnTGZ0i7AVkvjCTrxsPnQmXreac7zZhXzu4JSgYdpJufnQZstDrlQ6zx5ZsP62kBcqjlebRVYf9
51T9ONkayKM8ZjOMLEE92kB5KADWUYplbfkcax8DmrWeR/CqC81ZIU8Cj0i4LK5zWnMSYxEZj8UZ
vinxWU/2NF12hhCKFj5fqbEzhURVCMF+IeopthDNn4YNAE81bqso6QHzXePeffhvSC5R9HczOU5C
CvPWPcmK5WjfchbVypKs2UiIzzlYKklQdC22bgaQrLfCAqI0/otCpx7eHvJ3RL2jXghwm6asFwux
cQyEfFst8g13omkI0VXKa070ajLH5yeKSuKe51nNT4G59kcdVLdo3tkro6i4iAOElGOo4JjInHWv
PfNDEiMJHoHpXuPZ31LTKg4PrahGJB1Adx+wXeHREgP2DkDRiKWIE2hXRAKUbuP7WHLlZSZtY9X3
n3Zh5dGs3WJTLYR2vmCo4pkfPXYrmPvBflw3kJq8GgAl/dUhc58U1v1+Q0L93Ca0GeZW+mSf0oMw
DDBZjoS8/LJlSuF5ohsgH+f73YpEh1/MoYtdrasQdJZlbw/QRfHCQHAitBS2zgTSTKTwSsARnHpo
P+fV60Y1RMZC3HSqTJLS+wjH8B1RQxfJMb0Ihz+BvqBmJHTYBLXHHf7K3HsBRTIv/lhc1aKuSnFG
Z7eRX0FFQL1XBQ9GXDoCeou9z1FvPssS1fDIQXjPV9KtdJfcJPjWEXXRnaas3uRthuCjKN9VsGLa
u6WRtKK7GWU2IE5wOPbxkt7o+kYq5dDjn0y9vEPsc0BhJDUYBNgc7s+YsQkocYcMgdbqbpFMoFmG
n5PMtPEGFiy5yHSTbjM6BgJ1WpH6N0jZZhEe1AtMesY3GR2iP9BAGxzOLaiSLsd6qX1AB6j/kVsu
PbsyVWhAZVGIUytgucpGiiFqi1W26hZI44Yg3mTzygFY4SSZMmZvSnzYaOhZEJkuOifVXnGDkxXM
Af1SnuaFGVPGSX7IwWO/tZ/g5IyoxjuNfyrCtjibnouDIBMcr1j7MLknCJHKokVgCnTIWdWQYJwe
lpu00hVXbKPYDAH0uki83EElzBrsJZ290ngHne18Ggag5CG6S1/DXbAzyNlwmZ46iNEkChAwYgxB
ap6oAuijQvhbZj88EiwogCBNEqEZD40aKG64HwBQgxZ9Ap94KZHfFACnGgZi1b1Rrw4HDvXupcoD
cZi5DXn8cVhKp8TkG+JViegdNUAG8HHgrUj/zREM3bTzuLZYeoPqATrS7mVnQk+Us9OInYy6VCSD
N8IkMhtAfHpekNvrnCz91z/K1MI88K3YXGE+h4tpLjfjgi31A1E5YQljQYz10+VFqetb2mlETsfA
vPVs39QJsgeYhm4T+TQK/3rRs/9sOELoLpg2f+P+kQ4vxwAhaKFeHl9iDXB1+9D2fukUi0gOqDZZ
qJZPIFa3PgyJ1fAI/7qQPazdpwcgsUcIE6/mV7e2KHCTHETM7aa1mvZqfIrE8ZBvPI87nAIOk1Ty
+S2aIngaRwGfpHJqRzqeH78cweJxfEwtGlFhBSamI6yRNnFQwUEcZk5aWX+nvg3gO+8HZxLuuunH
IEe5448iWpVGiC0PeEZy8QQkeOL3SAHVmMI8S799rXSUHIRsccEmqysnNaez+0LYma8LQ8UBbg/i
5gfYCNQNQFulzoZNiaYQx8t4U1rIGce6HN/FpSPX1+sWmZw0C36UCliPj9vXDQA1WTNsz7gJJSf+
h9dW/rH95FIiNKhlnotspNnfG0L/B+kSWbcm78InRFCOxpDjxnNUZ2LSydE6apwxWrJrnifVjsny
MRUVHBYiBJ+KQv34pEEDm9ctFK0/1GdBF/VmNmf6vJdJMpRXLxDU9okb9oxYOMjzX4Co3L5FBMVt
8RHsTYZgkvCvisINDYy8WuG+7U/ol/MkZNvJLBL7nQ0lzgCgGKN3CbMSjaWwSirB2PCJmaQDMlqu
64L/1Bhaw4+rdpSQ+H/1VAzITIl/oSgcJJWIaTQmnlK6jB53UClnY/JJRI1NeCjKze2OGnPOFdZm
+naaj59/oRvKMO2geHaPfcHY86v+mrqIkmLSb4zEnb0763VFt/3aO4rvgGuEdRYZ1GNpvnzu5DJP
r94RBdJVVjkX+EkW62QMtJWIKyFK9ENZQC1TlM+pWRJXdGkPWurqGqd/2eB3ud4yv4HJTKkdrEGW
jrDMfT3/+nXLqHQggz1D9Mj+weSPFYbftUygrA+lT0C8nazv+UQC/I/8l+PsauJ6T5iGMdXgnMOf
SIqR4Lw8AHDtv3wdN00RwfFp4NNFxUscOvMy5pC9bnh5rzVNi6mrFuOSAW+SCV7ebYgisnCT96DE
RV7s2kwugvf+CgZ947mOcaUm/RxsHR+vaZodqzUZIdydVUJOfC+rEl2LhpTSdEmU8CjKu+NprqMT
DEbiPtc8jqE+QPFFaIKiVC+BhQeUHdS35ggrncQ9pYS9l2XM1FqkLxIomko+qMeFhZyVUfen0040
TxN5IwZPwH7AKc/1LV8q8Lzno+rUMaof0MzYgciZKqR5NyYL1PiHUiLsIdRxOp9TQjx4TjL3lOVg
A7YVN2OKoTfM/lNw89VeDRKFc1h9tA7mIaHO2FgbskC3BfMQfuI550Rsf2zyBkoCumEeVk1/YIo9
JIrKN7vCh8hynGymbYwFgdaf8sujMU9OWajM1PdTDmfqDHEda9p7F+lBDGST2aPQnPEBI+LYLSE/
zS4/NzIZvbbZEP6a+p+pwkB29NMa7XyPzhl97EMqNn3RLRM2I+tSv2rDEm3WcUYpBp6YYMCtDyhO
KsOP6N0BFReIS1/Ikr82ipeuvGQfH89eIpc0Lwehc6+U4XjeQqDSFS2pmdoQn5RXby8Pv6KHhv2g
G5pD3yQPYKoNvqExH9+HBQNbgl7C4Tir6x06KN1FWB9mY3XY9fhV8IXe4Nn2pG8OxBKx/iKcpm7B
1Xbdcs87YTFByMMAIU3bjufjdIAwppCK4xoOduc0clG2J37yxUgsR4OF1RQINFvH982UWDhVqPN0
3EUGk9UJ0I0rObD/sDB+0NO8pFnBSZV/umR0MXP1gtgyceTpxka4pz7iABgo1fDGmBTTZY2xf63U
6LwnrxYkNhHAwdr7AOxciMhWbjkF0CnEPhiDdSyMf+7X4K/9OAGem5ZBL2CH96pWcLDTh7cH0bLs
1YZ/lP9CGLNDiZ3SLA/pgET9G5AO7et78y37N4xzrE+XLga1FNgAHCvsUV5dUhpd5M437upJAZXy
Kj9VK+JcR/Edg5MEE++IxGyJjqjhsBSgbXWrNIQOySIfAk3JDRW4wWSsZnCrD+lHhYQcQZeI/yzQ
yYmUqkPzhtvoextUf8iokENXenZPhJU3t6vp8D7Q4trgb4hB4r8FtjxFF6N2mpOvFxtoqKl+8mQ7
4NWgQ2QiXzfWZy02HXbIYHu2hPEGld/pQiEFS/yI4W4s3j+g2FBEULBxBKIl27osCEryvjCAboiP
la7Vd/kq7Z5+g5KCQ8Jj2v7Y+E9PZHPRAJiASXrCbumryfaCISUqK2/FlHWGQbEn8DV01XK8eW3j
GV9kmVEfLT+FhaK5TdL0U+PX3K7HqZ/noAGifqWSmDzqA7TJGitA9/gZNfHWipXSAKs3BRSz7pFV
SwmgQK+d99GjJ0sTIL4cYKOIlFhR+IcbvRHuGZ7vVnPjwEoz+0izlyXewi472E7hK5s7cdFjNdq9
fAne89PXSDrC0abwsWdR/QV9kbvuK1dFZjEdk3M82/rLPRExYGaPukfG2AB4GYoqn6P1+7dJ5KLh
XItpW7kLWWzg4RxIlbPOHb61pq3+jtA6lFtcXKQo2ol/n3kCzWGiEGgJGkR0m4kPa+Hsbg+USjAW
jw8sqKUxvHKRWZgNrPh5koBaR1PATEbdxGt2sCQJ+vYdE+m7WOajJxWeD/1e8JFKLU2d6TXISM+i
Y6QYpoytEIX7WWK/ccN0PLQo052fyMjvdM8ArggvdTwErVYD94WJzOp1UBs+AmHDsy/UiYF+F9cF
6x9R+kJsR9gT9NHpG8dZgMRcjtzYvKjn+eVWI1H5xWIywt+qRLHVXurK9FH070Bh28tbABp5PW6n
QLqudAT4q5U3p5G4UOM+r4KtxqjI8AV8M7ExZwl+UiqTBzV/YFNIqB12Ip3je4ngUZ0kovrfItUl
Oe9SivSW+xV0mQH3NACdx6w7Y3QYo82tmWb4SvEuO3OrLFFE76Pf/hMZQ4R5pBh7heNX9A4vElWX
IoY1E4z+DjKi9aB7Gv2ltTLGU1g9mA1mCysko9sUV/MSeK47ChLFtccqX3YKDb3dD6ND7peHOAlu
4Jlli+eAnnId2Igc4ZOhCYdV7c43mGffDJPMJhpSlaGyd15x7jd97yzNP/96tOc0t0kHAhd+6iLg
e68owUuIOA1DJNymg8Izzk1lywTGcQr0ScJHMDcwM8UzBcN0l9/dGRUlt6SGXE4upfgwpfJj6RqY
llnEVRARc8dI2O29yjcPWkas8XmOhq9nmk2xEdDWVVjwF96+UqlPgbPTVkP4XYsOnxKz/cjoBUAd
E2Tw9mqTmMIyt2C3yxIPQ8mzHmEDd/0zhviwzcMqY3/aXs9FHLG+6+9ChnMt3H+y/HCabDtsM1v3
Bgkz5cW/WgQBAj0giKArgHfpOrdWSVBJfUGNtRCmXy5sZUp5iRANgpjBVTRJUvYBaGRBc6YPTjOt
y9eit1mPjwwPdKxHXV9Xc4aTgowBJAonl8EoA7jpvEMOcSWVe0AQlCun6hmE8Hhw/+/DpBLNmUN8
ByVcx809Fm9/n3+tt0d7XRrVjWM24ONfa3qCCBQ1iSMEETPe6BPs60LY3B1bPBQkHICrgxYfX70p
YnlNgRRwhyi2HdMBw51WaqvEr0doUbBCKKbhKdZ7whZfsSy2DJnHo94PTddMjKYHKvFVh5eq6Uml
deUmC+EyFyFouSftuMCTLtnyfy4WMjTEbzErDHQ/i1vdZvvA4G7mrqsWL5b8SyMaePVfz0AIYkNz
T41xDplgYguOLikEy3XbZwBzeJwq1XJrNEZLNsEoPqpiNy32PGtOJ3GmlX3A/FBWTnCicmAgxziW
i3/bVN40ttDmDNnBWgF1ifaEdSX20kSm6OkGNhdomyykRnmCTMPkGfnO2i1ZtW3mcEHLK8NNTrrg
0kQbZH8R5GXYFmizFfSl5hLFcUev7qTdGwZuRoWYZyxODH9kcl+1pUBYJaDvSPQkylMMJH4cg2XD
1S7uipE/DBtHSmPqBAF461UM3pG1R9p7wAPLBPapa0FPkgW3yhitXCBrkn1R6pifEgNW8BysB0rD
3g7guKKhzTgoBB/GzdadElwIm7sPo8ZK2cOosfO88d6NNL896NQUSSb6GmtYDXp31sIIDEifsVXt
u3o4jjE328uLSYqbWANTzNTYgV2C6mYcuQ9rsOsHrUY/HgtIavEkTzpxcPDzfQrIwlC+ON4zKJbV
d/tqa2+1zR260mLwXn/foJNHlVXUBawg2zsrQQDKLTllujG+nllefXi41Z7lMwBr8o/fd2Dm6Are
J6o878QPt+5mSwR3D7Zxr/y0lmg+yMlLFPJarwiSHi7nHHwDuLY61Mn30jjZkw+pOEdwb9ePlkAr
xXLIc931zWN+nx9LL8GgVJimR6HfY/Zd3YF0WU310geuHX4PzKhqGtzmV7QzRSIrTbigJbfsk3md
IOdKbTpV6/G2D8bXw3NvrnaSXf6IkgBSU9fdeI1Pzn/2rBDoDvQdpjzpq7pR02GGZh8kfmrUClhB
Tg920Yd8WB21RQ1JwVHzweu2sPCmK2rszv6baevRBgz5hyg1hp1CWw7MJTyeo0TTHcBKKQdnwWxJ
vu3dC0qugpIgb8j0V+z4SxEondWWlRyqAn0lPcWyPjz6wzGH9FLCZfwIZGGt35Oo5VdsNNhwYeGz
OuIXWncPASkRaGmuAGnT1/eVU0O6A2LAow3IC6QsvWmto0lnf3jZrDec9QosIJum2tAmmC49ZEQB
dnKbETYl4vNhT3wi4QDwCNZ1/SVtejJmXLFQvI1dfB3rcqI616+Wi6ExCGg8AWfqCTNGhxQMP71H
Vbui7fRjP57GwlDBeua3r+4cKr3BWrEmANqD2fFe2XmjUXv8wJGiVT45ShU74Iubr6MpUsAYBPvY
kxQKECoA135dj8Y16FWiCOV60TG6l2XIGYv9+kkWQ6ftR8jplww8Pmdk8jQrX8MaXBx89HiEmFA2
hR6Lx8Y0Jbl8OnWIwUqbUfkyYEFKI+dx0EZAVqRwrpHYM/cS0erqHsABTRHz8lq/zvzfM85Rjvd8
kuA1ORQh5bpz0a97Dyv5gYKnMQ/9d0UsJ8RhZqszCqnvxMlOZWh1Wn4/Bz/rMeTcufKWOpeGXKy/
1vhfgBaaBbOKwCTM1THe0Bf27hcXhaj5fT9nglXdf2ojTbZ/NM+eX1Pe6+gjCpDIaXYEZZrkH4sc
jLl5bs+zEqb0DC9ZHWIP3aDV/Yd42bFCgByFYy1udW2ZmFpXri2UMRwh7TswP5O8t3DSAR/zkymj
x0D1WuWwir0Xg7Vp214KPNPMkLwKjhmIx5nwBxKleb34ptBSQP2+9KNDKwV/xPUoQKXe3Ie6V4cd
n3yOGdTKh6bIUR0/sR1fHerR1BLDNciESQiXFXloI2Dz0RenmUA5LnNW5WYMTml9/NvPKWlaPHW/
oNkrQFrmS5oZazK1HVVzrdf8uQAUlMGP5Z7/2CcBeXsBiJVv799Xz0nv/+CV8bN7TG83g0oVe3Cx
VPutsoy6e3iFDu8ICyt2vf0Hs5KCNfOD/84STY+1fDTQ6e0x/Kjd2R6nYmOcdRbWGTWZe1rkYPrm
sX5kj1bHTfww8vEukz2b1RJC6boYbSj5Cmcf4F1A/WCYQfN5+bdbg6QqI+iy9PR0lUhk0qmMEi86
tNpbz/n0mJhRAV9E/rVSpoqummxWAQ28vrdiVmF49qPcoJjuNK3QVXX2kziIJQh3QHedC3HtyySa
Pqd4PwCCz2QfAHDsrivTQVFfbFydjkm4ykRGDMwxrNoJhSwuJUHTUd/Nw5n5q/uZwxTQKQVWBCcz
fPozDui1XJf50wY2dwVouaWCDJwZc2JITGKO9etZMii1s4KN4P0AnG+17lf80caDlAPZcHcZuBB3
xplnYdXYnEst/MF2nmCfg481GG4UeTz8+SmDBXHJTeq4xqRDw5UUnICddmottAlYKmGqhzzGGdsS
KpvCvD0HXWJgxJE7ndUUs+GVVrnwffPgACdEQA2rUum2gauuzLa6ez3fO1JZ5AQCRl5cU6iZA2Vd
/ZqKgHC9FdfbxMB4s3WkQUlLutCU1A8ITIZhSh0IvqrcrahDnFheUXdWk348YXMedpu7HjeQhXzk
VWIOCQ/g+0dq4u4We5+aArBj1xG/HdeHvwRRWCWGCMUErr+qYCTS+6iK5nQTkqcu68pN83EugTR3
PxYxlKHTObFsCWbB6WPFCO54jUn78sWamr9QTODTo4yoNwLso7kG8fN/ExvcmIUXcZh1htCmYLBX
0JyHwxSkAqL25Q4lb7GqOoTkSKOSEpHKiHrHid/rZAE3TLQINdeN707kNXYPr/T6/Mtng655AiLk
x7Z3xP8gj0+cJaudyxwc1SI7gdx+JEHkwLi18ADaTdqTAOz6Yk8EXtoZb5lY09siv9XbDGEaiKJ9
RkifcLQR3P0+1aU8NeLOHpvRYHpJTS1ZaPOj2yOiMCbFxTrmToHCJkcatmA3VfFe8Ao5y/wEgDJU
GegiR0701kmAU8NIDl+3+/JYQzmE4O7OIWGuPanPvgQATbSaNPrwSQI0yO7oD8VrrdVUsXFI9/HJ
/jRrgBz22zgYh33vMYo/ItM30OiT4FnqKhP0gstL18D4YXW34XXSBv7jGxna3KZUiBGiafaYwMkm
E+u7iRYD3FaA83V6K9xJ1LImQatAdWnzoy/qYvTBe0gApP0Iz3whbt0Z9xr9Qssf0Twlyt+b6IZC
ugqE8U9s1ibZ2HB8A3Z1/tw+V9lP/M+woYnkG6wmjg16owPJsoxRJ6ZUR00npXm9P5Zql7Vm3Xea
xAbR4axCe5JTJQb+N/pg+gdsHsHtx5C+/O3qJCPoY/0GYYKPy3Rj/BS5SouFEALkI9xREelbvlKc
pXtlb2jRlwEtdXGQfnpJj+7eJCyFMBh0G3KnR1mkU+CJkbhZCtNvac4KEaeEdM7egFjyarV7UFw7
0lP6CnPJFp3xw5ls7nCmnjrWR3hPM6r5TvhNb//i8bMqWp3B1lmmNOXij/MKm3K3I6vvKEKZT8/J
aTw0nUThM2K/dnI+hwFX4wGQdbtUAX/9dpzoJkGpE6ydPTOQHkOCELbWt2E9kCkbTgi88logiKJx
+wxQTDNpHkF9qkdQu82DomfVEzqTA0be/1D97K/+ZzE8ff4SQKLUJmb346Ms4WXoq0r0WpuL/ytv
6foMKUIAUKJtgjwMXjXYo1Yob8voHAiknnrpHjmtdsMsktYxPJg/pjFmwdKRpfCiUyDfZuvtyNxV
2W6qbGMireLx/XWPpxYHGC8HWxvjTLdN4u8PR6nzKbqhfX5KDmZR4q9J/gKmycUX3cPitO8SxGEg
EdXNL9LIz1hU1x7HHEu2pku+q6ONGe9Pg66hs9+6jyIjCF1i5k+ZhZmqLCGnBp69VzOmnZhid/3X
eUc/mfhcsJglYC//YxfjqNTR1ZWhCCyJvQgpkyZdQYMcUDgpEkwWpjn7h/lw1lSoeofa4e8ILXO4
9AfQz7D/dx1rZw8MSlPW0Fj1j4EsdtwwwnA73vF3buOlizLP5Dr5YbGABXrVYAMVvb5mum2Yilnp
QtGZ22j3RK5iqjdujn16sTPrwLdDVMNrubOMKomcoc0ixS7DmM1uivmrMJn19ISjYo29g/qyZLAW
gYbYKEzu6NeCDUL84hQE7NVwAQ2eBRlcuGG+cMuqi8NcrjZwtKlF2UofVrLcegTyE2OWaUdyW7mh
2ZLOLJte7ohcUsWIv/jrD68S6Zmh2tBqM5PicYJokVjJn79avA84sBdZbMdH55L3I35T6y/sgRwl
vgVHA0zAx6I8u9oH2hEpTx/AVf34Axt8xJt2sK5rvTx8JqvsBWZO3Z43Z6xIoM/DwhrOBAv3Kf3B
a9CZok3BJYP4L0RagOWeWaxWqa3Z/Q1H7erTWO+pSaOz/PaKnB6/7bxI++qbyHci7DyBU0iFcCwZ
viAcOoFZ/zqMFgYyazLQQpOHXydi45nWMwRVnkZ0acWrD209NdmSKw+7vL1vkqT3brPnWJSRpPBt
bE2+8gNUvsGPJvj23jpOIg2kFoWs+xIZhSp5PWg27gOyDACz27TzaHs5XeZs6e5l4YyPCKY3k5H6
ALR/eF7T5Eiyy2tNtwAKqxOuFkU1K1yesx8fBKDbEE8ljR2CKEzVS2Y4tMCxch3N/LvvzEkrkn17
Ykf5qfhms2o3WaL+/cB6EApRlfyaoVSV12ZSDf8guUalYfztdq/H6cCilyy+WiKv4MuKp0KQs3l9
L60Z+rhduNBpUd5lmIN/zA+QCADiMnjmf05SxVOIxfUrgHIC1ulkP06ft6K+dTF/v7AVob5DuBMm
kijgrqGYGQLZYk3L3pX2x65kq6/WRKJK5iKFrJ2qQ8x4zlZyzIAGrH7AlP6bYrvoXgOgGK++apcs
PrgQPKpBD03pJd7wtVpq+5A/LV1k3UemnQbBwtAnwpiux3F/vcKoAIYbmIgji1IllpIwOjvvkRLM
DoAFHVLuJlkswgigK4Ikckyr0j90rBJD9jOuZC/lc7HN2DGqfoxFc8+icEzHXr/vnoFdLCP3SEAX
Xdc9VA3+WK7HetW86Y5AB2lGcreDR32CRZDYBC2XIh1H7X4xuVn8nwsJALI+W3LwH329QfEQqBWZ
j6fCAPgS58eGIXr0Y9mBrW3d33RI/yZS4tR3wibpL3vurSFrfbloMbcrScL5RbsESvjbwCZ0Tzvs
M15pbsdoOAQ2pay7psMWGDvrbM1V1Nyzh6xseSpmY8iO0Os1oLcoL/egIZaiRpr9X7K2eOQmbmjt
SgewWovIZnW6VCAtvh67n+JeYdTgGwf300L+3wKnppdNyb2zS/Xxo6LOIqm9t/3bbgpHvmpuluGw
CrYXBUjsUPSJ2kXgOKqp9q5N0ldCaTKxbthFeDB3BfNxeqL6LyOuMa1Ryd9ZmONBZdDYa+c+jzX+
fD8NlcKllOaBukNq4ubKNyXimjrMoQ01bZU1EMbs1XxVYr2cwhR5IIzFDOoeQgz/Jp3CIiPrhAaZ
8uunmyyOtDCZR3q1ooW04kC4WRxN1Y7ySkcsLGVIcla8olW+o5/SAWLnL4yBb1KnfqSICw4iMwJy
kx0er5Wg60DU/yqP8yrXB4Wvi3weAeJPyOAZkXKOJzvTM3WNJAd2r7MnSl8xVStR66qCvRZ7Z2gV
aB1m2QqJcj7yORWqWVLocQXZHqesP6qQdzSQN9cahFwuaWbJxJ7XkXU8H5Ai4FYSd8BaljEOHY44
Q71IIgS/n1NiR9jWkYrb2bilTRLW+DUy238SraGavNGSj8HJRubJSaBjriUw9sJU5f42t+i/Fr+F
RkVAxZdRVfJ+CfSZqvJTzxP/MUtPJ2Lmnw4RVtojMuOPd3K981Ew0iFDH6x7h1itvZaX0updR/O+
LtvRP9Y1+aGOhmWCOvxuW9oIixpvqs9OjRtcALk3Q0pwXNjrOSkLvB6se0lFW1Rh1qNw++nmhUbS
kVperJxX+L6ITHRl90fRfmumzHHqihy6XOF1SfPCH94SzMaAGXZX+AEqMQOYlha9NRmXnXEZ7A/M
aNX3B7GlYM2AwcWnzY93Q0hO8TVBq0FxSV8Hr3AwCrNdVqyX2oxH/6bKSe2F8kuG5RTQ1043uTvn
LLipfaxFqLEAuam9/UcFVivoMGN+l0ZFdTKUH81r53UkTkyiX7B2Jj0RymR5TYV1JgEiKNrg8nDl
UbHs556XAIrxcrTrEB5Zh7LT/3FoO/QEA+GGwi6qLVSLdzeuUxn3SFv+zUC2uIg0Bvq5UGfSskBU
/810gv2k7VH96BqkOgV8tmuFw1pYgv3gtm9YrNdevCegbL6iIQJpaS96IbgFATRPFI2Jb6Akg65L
27fRhsEEMffFKlMavmgABDK+T1Ao8NSVepf4YJvZTdvaRKUNEUpJdn30ZnERE9qPnRcRV0OHK88n
NRkkb5+sEfg6jT1vaV/6k23u92GxcR37np+98ilJ4bfAaX1fo1ZvyTtpd9Mh0P61POmayGCVcT4i
B8jLaocecQe3+hlXuWXVw6Ky5JEU6njFS3N1JxB0D5dkFvjUrGKT0hdomuoq+wQ82tSFmX1KU6EL
8y4C5YBMAhLIz6uf8Yvw8I2Cn6PmblyVLTphfKuGMV9ABGYBUs3KOVoRru7NA/fTmRyWU5fLyPFc
g3pqo2D4HaQcPPXCwNmdafM/Bk89hOyX/j3gEbU+nJ99w5NqDzdPD+qcpm+yUSFBd7GW/3ykqZvA
PH5PliRZveXXbulhZclV3dsV6xvP30TcHZhbqrwqLVVUF26ZoaB2kNfm82IX1qtzg8Gk3aL4OuGd
otlhWqS6NkfLqrdQSmnZz5zMuMYADD8gV6yeESY+CJ7p6hsT2XECc/STAAJPs6vrRWWaElvx22rY
iWJgLZkFpYM7WsfAoy+6L6L3Rs3VUPJX/MoRxRU3ZxKzmv23Ya55bxlpp1Xk6Nj7I/ZfqqiBwEnR
RmNEeDH15nIMnfrW5W31Cn2y3i6ke/x4KT854zjmvvjRZa6DZ5ZMqmoGbw0RzJ1IM9vBDEwrVa5c
rc9netZEIebV3dfbpO7pfWflpErMarMJuzIIm7/0/x5Svzz8GKbVIzumR+C76LrNVJevEJWPk0vq
co4K3gKIPpBqcZJre2QsfxhT4M6M1CFn/USmtN+TGq9+BT4LLuUdPgmu5HctBIHTSbFUSJVrAv0H
1NyDJ7JUKVr6GujIkwfNQ9YyzYvCn8sV5FW4eJWCJPWsm8FmS21+8lvfhq5sjH2t6Vi5ea/VNKcr
3ChgiYz2xttj7Hk3+YeswI58J4Tntk7gPfNsfyAByaaBmCN1/ttAPabkVe7LqJ1cn2mqJxulpbLi
LTYcC3wP+qvouDmIfT188JcAiN2bo6DEJOTgGaeyIIE9ku+S0JnmY2BoOxo8XqrJZj4wx1jB1PBl
sHDHySu2/PaVJJsJqBr5CTr8bAHlZ+s0VBzR0YYpjwFjJGbYqCx78laks9fFrUmNI4RnK6OjZHhb
vNhKSOMEzg8DcmIICVF+t/6+bW244v+Uq1hcJOvAUlbbGcy5OQon2aGK+a0rMH9RgW+ep/UyCCjv
MxdOoWH3P+BoWSZYBAutD52KNnEmAYk8W/i87SulhAMGeKs7ekNykAzmqCu7+m5qPqUxBtTqWnW1
qa6eDBRfEA+s3MB6TFDQCGN2/AyMboR5n9SejG/Dlf/A7AL6VpbaGgcsE0DU3+lf5tfl7WqKeIeT
BR1shYCrF+/ffdmsf60VdLE2/3gIYnk3y504yWAeQzrd7PPSBkWq41K1BswdObji5jock4MEtrtn
5rW1gciLcVUoA0MDj5PsRQ8E70upygJZEdr/ySM66LPa9MvKTil69VJrd+8n7ZkFY76Zgb3HY76F
JuSj20fPe/W1bBwtZ4t6D6aLDxyoT3kShtzKTRIlKtFGBy5oEnViKjUng4QGGGPwHPfaR4qOxz/L
hZJS9tz03Yd2KvT4n0TCR4jY+WWTWIeCgD0txrnIsY5jFlPuTLNuYNlTAhZG5qS1arlfTPL0tpRD
hPA2Ux1SUSt09aAzPt19+5p8WVan2Z2cqenC0iyfm3IrvmQQbR9NsYf1bL7/GMuAoC5xPft6FxVQ
//GBJBWFsf6ASnJshbc8QOVr1VwNjj/vRW3cBm7eupEBotJ/17ISshD4frj2gg0FXXj+v+BwlGUe
lF7kfA/VgD1AvQWilSuaPsaIM6+1zqoaUzuCrXY4mZ/Kloh2pi9lXHqcxgQ3z6B4ZD+6wBriNPdT
oLgEUkFf/8sCjnIPC/qaE6RbNUwbRF6krtHpPORz46uDNcqfwfDFL4N3igSe2EpMwq5lCbl5Vc6B
pXbOY5f8mQHtXKAiGp4RfU7s5yWj3R8DPS3NBqkjcUA8EGo34MFEwYLT4UaXvEZMIuaeT2jhmV9w
76Jsgrbc1QM8F3n59qJQBiGjCUIcEuCdC6QwGdOxDyvJ2HHu4E0loK0urUd5sONytxoudp76PFlN
PBXb9a46xCApYug9cNqQ85kX098RZpWt+nZilTMnK1134NBxY6+kYnDdiZL3xF7gTo0vuRA0Fo/n
MgMyDycGO98xieArKiqk6d8n84D5gFAuMwrJ/Vu5uuZxYL0yZPZvN4j/UWEU21NRUAShbGwBuoRU
ewcDXJ6qpdrEOEtuzwJE10PKjcSJW74T0qkiMknkpZvBiE4W7JZBZOhnfc/Zld0wH5T4JCmD9TQr
d70jhCiZpNPUHBcWuZIgTl9wJTqRiRMFi2ew5eNRiavMm/b0ZJhjN4oESsUhRKdHMxKBYLC7TM6J
qLfAHlA+omYogii/QBvgToak5cBhCVbkMsM0j8n0/OTRIKZQgCxmesUUqUzl6dii4KLPJUmpQr9s
lgErsrRI1YAeY2LT7Sr32uALVE2rdCxoOSXwv3M4LhV+TXJ5uWth5a0hw5Cczjpr5QicIO5YH0xp
3KVWIViC3B11wCoLiYxyJvW7IyogKJGn3cIKL71Ah60BJVdnB0nMkRAmL/XPbW+4T6ohU9Vi9AvR
XTOLsn71N6divXO4uDDHJ/POV7u+6OMJa7wSBdvi7tuMglGg/trQyHI97u+GF/RpGXGDoH3aKK9Y
jaXnH7gd7d3C7kY7QIt55hBjd3dV4q0QhW/OTmLxIzHMuGiaVvjF3Nd9MCAberDAoKUiRoeekiyR
PmbV76pODjf4YEjgnqns1RS2e+XdbvTMJjuR56EOP7qFeEw1Y9yHgkSGtpUNnas3OEnJoxN3R3ZC
UI/J3UWwc5CurK0NzHqOHG/7u8z2Kgq4SrmJGEUwWEbjObTBn5oVaxhbSbe73Ukq2Y81FaOGmznd
zPQfMOb/dsCCud/D9qiLTshEyC/A9+edQx1ccQl2+9H+HbrsNykZKmQFK63bp4agbdKKQeADCBjm
3ELM0WIh/xJIFlnlixkt2UPJmjHS7GvamluH3J0FHg5K/UAmyY7lsk6JOXMC0WBb97uaj2iS4F2Z
kf34LEXA6J3b8ToygCYG1pAXpulPKYEkn1qHqkqIcCNpP7c3dUkxToXoirTZ/+w9FOsi3wQjNP7Q
pw6MVSgrEBVEWKhqYuqI9lETwAoYAnbrv4wjiJAj7RyRxb/16uVIsDP+HeXr0Q4STQDwATgMRKYR
RsWU6OSZGuypiM/ePvabHIPlD2xxbdIl1xig2UFSMM7vdR629V6nezcoIxzm+AEqtOPGyvqDy/b0
7nAD1lgywlR/FIMLXkvkudB1036DkrvA5BetSPiB8/fSs8OGsxCZjGyYZt4oVQNxQzSt6F5sxGML
G7vvQGE8I4iYm5vyvWVonk0BcZE8/MK2WQ3i1Jc/XgfRHJ52F7TRfZBECUplaWowtjAYSJZjkuIH
Pd3iGnF/ABPoa7zule+ZINc6M1Tc8OuSmJIiRlq8udw0NNTq8uV0zgkOKwVlphfQ7zKJPfd9l+yn
NjAaYxqMuJd0aQEZQ83II8gwq4m3ZPQrgx9/aRhsFOqt4u/vgnBxEFhf1rvHjuT6Rt7MBSslq0tV
+zBFOpboZv94O7sXanov4XHotq/64y5gKGds1BvLrjOMJ38WFkhkaqMLciWo7Rl+gslOaKqX8NjM
51MHGVcKUyh/k7SUjoYkrpQJr2QA8ITvLUoNOyBDwS53vGIflhm2aqvFp3c3MjYq98osCUb5ZnO0
Za0S30t6e5KvkflfIoFhdq+kWEVWHRvKm5Ip1fcp78zoQgQlHChrDPHr8VcCXhSuxbhuW3RG5wNG
KiXrcKwK/rSkrYhZB1+iBJzIV52QXav0S3GvyBRmdXDptZvhRVhApVcvcfzhGhRNrwRa5OzX0Yq2
owXw0wf/eAqPIsRgAcUMu1HNOmg5QdsuwRO2wZGEt87k8283s9WC3Te+9y2y9IJiiHoFR0I5Y4Wh
JjrLRhZrKEQpR87WzOCxHmxaa5iq0emPLKjhBrw25RdsD8nGuqJVJDJfVFinUZUIQPYA09zA3tEg
QS3d/Ve5swrfAvjAdrN+bJi/D/Y0auOWOSTzqHYjPmafRd7JjNQSKn5dNHC2xzXTXOw/olyvWVlf
TEzv9MMlt/0/MVvgAD9KUbdcGzGaBPwx7GwdEkJxFPdpGN57SOSA5GWfpJd1zVxKDRLEjCAvB9Z8
YxEslKr/AWc8wcJnm1ZnQq588Lc0nHj6hf4YLaFO4FTVZZ4LXDgxcA3hQ8Q4cB/8daxV1MS8U9JU
rrsLMdDbiwe4s3otUo7dWBZXYIxajVlCSHLjeG31ZEnoIjtJleTSGHqetX9XKsAmqudQ5upr9HAK
eXIPIIjgD/gqMmOXCiJ1l0uFNo655dA1ejJY2hfb3TaE6gYR0a8SsQGy6J7Ufht9+deo1Ojt0/JB
GJSr+qPjtMmYPh6mUeUF+aYkwl9PGA9sZkFUQshNlnNNVQbi/mERW/whPw7tS50kDp168dW6YxqN
LDSukAT2eazz5mTd9nZx2dN2w2DLPmPaFr76wRT0p65MoYtLDfJ0F3TOgWmZJAUD1E+WSn0HfVNP
VEJjTKkab4fTDXjZGdDIx9GgWOgTay+q3/G4D3Kepe/1XdeIeAAu59N7GYQQIxA0+ZnEPFkZwQO2
lVwLpBng7UEBtJY0XKbrkoseNwSg/UkON7Kx4dmZ0TlSPVlfL7JyLLjFNfHmGAubIcmqp1RCMpk6
QuLuRdhgmqeOcOFSlF2R9YFBpfZ2G17DNt9XxBykClhukxZPRDvln2BcIJFSX/fVUlExkUBeS9VF
5bphdyZz1D0E8xlpk7utoNpkAqeJM7NEY6m5yKNYOvBWt6wpnC9ktYeJ9kwZWMcl+LOUSTqIm9Py
x1r4j4MdK2r0DLgYnDtNrdsThtlR4Mrv/3gONSJ+zMP5SP0FFOCu2q424m50Tt3ixWBJgx6MB505
p/7BsFC0SOC411LEioZ6ii7n5cx380IukAJxjB0y7tDv8IW2dLD0v2O3+tYMfSpWzU1IhrL7Kz7m
TL39tp0gkih2ui4NQkFcMo1wQq0rioeSx6vIlivi8+FvbFId0BCU+mfKlu5ii/7+KBys3QjS2UJT
YIK4XaAPruXM5EyXLKbRe8Wa8rns972VYucHeX8R0BIIhua8fR+yG7ytLKnqgENdhwwR3xpFzcuC
9Egte8Umek3oQ01ATB3EArFUdj6iH4vlZon7rZ5GyycKAyYdN5CgIwq5mdEEAacxyOI52NTHcDmT
bn/m2XXmFkiQu/Rn51jdE+pWldlj5xcv25LA6hBAUkrhCNOzn8PywhMB62HkaZe9J1J2Hg1VBF/D
yfn9nBTSD4f6TjtJ4Ri3mSRwN0n34PiFvJikem0msbkxm8saJfYaHfIwFJh8EuDGp21pdib+2hjb
+NQNRuYE6A08XHKyOXKSc3Qv1owa31+t4c2GKbtdK4St/wsoaVNU+1csAC21XQZ7megzV+LTbiiT
OcSSjh7uaUlGSue1yI1VlIlF9vPDv0eOGJNOaUg/C795o2Epgat0nn47NCkjnbKlSR8fGZBq2dx5
V+keX1KZQfj503F8Guq7hetHllBWLpZIaepDA/UxK/BClT1Rl3bj3bHyPPXxG4DO1pvHF7gJxIj1
YXXor/kOL4hktde9vDztGNiQQw2eiw/nt33YBMdzl/ICTIOOTape2G6DPPfshxED/+7ZqkFNDZwU
7o5gYO+KSwruwpeWgAqqIS4f2bjAm1tOuoOMSTerAJJJkzvWjvqy4haFMhQJY8Q1EVr0MAXrcbty
W4nahIas8rNGRdGVfW2JzwfyrX6zkWohIJKQ3XayHytib/O3FWAJtc77la7j2NtzOX0J4/36tm8U
MdCl4Vf7Q34/WEtPaPbetvw0fyJa66qL768O61+uVTtk+wbt8UEmdt8rA2XpxQ3KOa0H98QhHvCZ
8d1guvLYscaeIu0pO2LCttmLBIyBcRvFbw3V0NvBkcoq1AxtZb4gC+t36k0c0/MaDIVytRU4P28E
EXekZvG5txRayw4c9Kn8JuvCziwm7suoWLEK32zS6hiRaUvWm7RDjYJDpJwAW4qA/7p/z7aWbb5Z
FlppISh9wSXr65V3R8IvlvzuHI7APQoHxTdKdN2WBgF4eUjSWfzG5G4AGApKmuOq8AN88zV0a4hX
sdTMk2CE1l+0kfw8yxPfz4en2UHYVcPoHa3HkJ0X+tomdVLUVdvWRbGok+Twz2jaK7zMdNYRAFPK
kIN0+GHKMGY7Og2+GTvx8yWiqu6jhJNJtdgPYMcffi/Dn7QGRjb3BiKEv05EtGRQXwZWJX+qVQfS
L0wlSYc8nkBJcnyzCq5QAAh6JS74WUIHWpGfALai+lEUU3UVJcDLPvlVSySvhtf5B/WoQiB1qxSp
UexAxScDedrFUufuXtzGERa+vpbkEO8eqfMHC0fhgnea2orZ+M02s90RlK0syjhq0zjaW1KYOAS/
aztLVEsLTvwdmAm5IjO816JfLx5UPCQBXWzHpyOTt0KxeZav2T1YsK2OZJhPTLqE/9rYE5jO0KLk
9bB6bjUg5QwM6rU/ePyryOLbWA/ia6gNW6Gqi9MR9M7g7K9JksxhskIDGIJkXS707TLCfTwvvanr
iLzkkuYCywASvblADEqrxr3fumh/f/tvKHFWbueEFgNbbig217qJcIWpyyhQ9g0Hu/JDwoXfaHsk
ceURRAzaJiaU4cIcrsl81FT+A5lnIuu3bQO5a1PbfmiXetS0RLMqxACaqZl70q4i53eSy/SaDCcF
R+Wt8lpJpBxBRLvhjePFZyRGhuGL8QYqgGh/EizwYL2vSYMqK/IV9KemrvWvO8tbSjC8KTCMOrkQ
HcX1HOwbyHRcUZnxrOCmKmkv41KdLEVGEUXuJ+7qcyVkcVpyTBDsh7WQDuxdz89EElbzyJpLzL3Z
XGeKSdvlSgePRahU2ki7rcN3tKsVcXyn2b0z4yW3geV4qXbdadGoerLU6qZhCepEBqUbv4kvcV0g
Ry2i5HUKto9uc/AWm51Bxh2VXbzPYMp645UoKaiAuAtWsZI/sqdXL/N9YCbX6JnrEDyXZUKppj5I
hZgqCQSvPYzsZruDnarGbamXVsQXHelNKjO6ATtX3SKtvjAIWA6NQGISrxlDdKfzG7RlbJXJUx4v
4WKo28RJGq5EgREWMXrK0k1FOWdAU3+OeGmB4bmwcjoUdODeQovi7wHUbwGzQf2msDDzFmKp7iuB
Kp3ugXjZIUmAVPKTb6cZhCOaxlD+z9hdlqE5samJ/d+yQX/LPOhifq7NtzJvF7VgnDMiSM+gLK5K
DgHstKYZz6aA2heWcLAUTbY4SU45G4Xue9GYmVWY7Ri2bhns4du/zECP2OeYi0W+PAt5sTofHOJq
2amo29+c0PxMWd5ORrR2GpKN3voATAzG1RDTbtsJ37uqOViXg+heGNRrl6n0Zty1cFvdXZhOfp8B
zSZjwoKNpI6eKyabjssz7XO9iXOmF038tu5cyua+m4P8C7FGhmXet2pifGMDWGHqUPl19UAiti9T
jO2eOc+A6zMBFFV8pR8kgHfpcOqKfFmwZLkzFkSqk2I5jOef7KLCs0Ip5ecHI9pKo3eNvtVQUlm6
ek1hdx0Z9WDfbqSb+NlXxqI6s+2NWaL0wzQQ9+aQQ9L1wDlA+jlS6TFb/40hHqI1tQJ9BysEok/K
nNJq0MdVQZ9+lZdggdJY4O1LXVkxNCQyrRAnj11WdfwfH6e4ZcChcXhX2feUULZOpIZwwTKi18G4
2Ut+KaKSXZi/zIpbYT6QnZkK1GlQHfdYFfBR3Dy1f+rnYG1M3ao8mFpL8JY/ioKGCtBIunrM3v0B
c7Vq3+FxMMVtSXWcwHxDgut5ttbTrJZ2Z/spqJDVbYz/aEEZ+CjOQw9URYEW0hlcNZTGIyKLpjTp
9pgvvoGF1Mgj/4XLUONARBFfFW/NeZFIvQY1CfOdv2q1ExnF+h46kx/7EGHtPe8iJSiHD/IrZLjd
yND2T6QSKBw3wiGZyCYcVmIWWAUsJuJH8mzAzASD6EDU6kden2yGHA7b3EtnzwfUC8UbE1h154MY
LaXJME6YSMxjhsdedno08EMjVq+PmdOseX8X+/ANshPVhuhkc22j/f00cHTwHlJ3+glYVeW60A/S
6TbohwQA4TrjvotNum0VmgxFSCBbVgENOaz7yNO1gS6cAMaHaDmH07SzPLqJ/MCovT/712653uzV
HghkSupdUUERibk+ObLt6lhXg5LhActKHdKBtA8KDpCOM8ngl490HuoAYVfXmWBmQ50KdmcZLOfU
YR1CHm6cV4pJoSSWq44WLk7c5jXSYShRgJsiDO+HSPq1y7L4mI2CFMmNpQzGeYBaXBhiie9vUwcH
fypyfEMKBd/GUTOfgIQVhNP9hZPx1iFh+uvKg2EEa2rEbUHG77vORNk2x23R86vZMOevMJ4sm1eS
zyAQFnTTJi0hvTK1LX1so511pWQ8tft4TBWMTHwxKQVt2cuhPfm2unR0f4Fptgn7ffVVr7Oy34Z2
ch3DgTFi1ea/7vJ57MPUehxM08GG577l5Q4kou2qkGbUvqfygEFa2oYWM0vmE/zD/lGdR5DLxmTv
qRVUoxxFN8sgDFYWs4PUf5Av2a9lHcZWBvC/cmWTHLjqnIqMSTXiZHDId+lelJMmQo+fzmfAtf2w
y4pAB9jC4fdWuuGtCdYtKmEbuUFnhLI+Mp66L9vizbn9giyNLSc6pwpgyug3Bqw9kJh9BlU9j1sr
oYLjUXaf9Ff1QLoi12WNPXFWWxoZXukjhdHi+QuWnFEZ4WtcrDEKHJPGH90zOBkCyt1XL3+2rhIo
f01rhOG47b72o4SZhksOFQpqxxGnNikYwCbxVp4IN/88h/46xTFDde8PWzkVXSXoFweGuQlgwkyY
ih0QRpYlII2AGPUdNff0wzFvx3vBjdV99b5lFgUAmqsteTn+JaPWZzxLZIExxF7WtakfEJ4xbweU
105EhDa0fHGXRR5BgcUeaaj1o/eTAWCZzZNoRWBTLc5WyJCUy1RQMqYdfGg2T0Aeff0p7ukyDN1O
nIEzBq9WXJyrXu6bKi2yWtw3RHfQtRLRkt0j3u3HLDYPjoZP5c1gGRZLjEKDk/+6iaazQOQ7i2RA
l8n0RjOIwI2ZcYSlpm0ML2zkxGgXLB0rLyIGDkEPnIAyYTeL03H1NESFn2huCc7bda/2kSN0Dr7Q
DIVOko99E2ZW/Ixzjt04i1kjzg9gTVvHQ7OQa7iUeoK0mk08+3amQmT8NAkeOHyNTlJflWYy5NaQ
kfSRCivamgtG57PV2pr5Mwv9tInllZArpyToB9iBDvQSrbjWV3nIyhEPISsJa8rntDyeLcesUOre
WBChlBsBnVZ0VwV3GCcAbkj9iVN760wxlG601N3NRWqhkcByekAjwkYG+OieMP9rVOj+F3V1FnkS
84MWjhhbdT+63SAx/6DohU7gfYpKXbB34+fLwD+H5vYCE0MQcPjzkXNWLdXdiAyEsHRJTd76Bh/H
QrQzbvRJerm/u6LfdSVhUPjtcVxyONFweJ3WOESoV4by4psqspZDW6XgAD00MDiF4iY/2d1ed/T/
oAQlgN1Em1QMDNZZiTAZ07RNmwpn0vhr0Zac9CZ2Zgfuj0Xqf00ab5+kqDXuDlpQE7GmzfgJYPDb
ZjcVNN9l4sbmkCWA/UAihwI6yZvRibUW9FS2aktW74WPtOSv/h2FfbQnlAiZLBdCHkLHteRkAaJZ
mo6nM1t9KwgZIsaVv2WHUNjjIuuZ4AdGl8kVpVeWQ2FxSKSok+55fzUONU+BZjvqwODAYxD8SfGC
B8DFIV7T/E20RdGlHG+a2ec6Y5Hbk/TVMkWhWXS5S7Adt5ZmqwaZ8dW/AFZ16CodNHeiQwq/PZpE
WnQ9vTPNny5avydt2WhyjzQheBCGOMUQqj0beLt8wRyyue4WXxjhKxkoyEPBo97LaxKQl57UxTlo
cxgZYyT4FbMr7PjIZHIasF4QqFkJzslSM2zcYsl4/vw4EdlcJKEJLtz6AGbA8oDo3nAC3oAU8xJ2
hNH5+qLPA0GBCo+XASo3wGt4vRzspWwGYY+MQCYzWkBpaw4RY4lrVMXuyrsjQ3MfKMPMG79aCOF9
1hNC2ZdzD55t1BTeI8KIahrM4T5F7Ab4k5zN9byDFQBgmXNBA/xqV/00SS5o2CHNv627iJlTLH26
1VIdwSx0GoI+SCQb5bkC4KBoHpnpsdNbhWXsWf2HXYJRHEIUuywrmCTHDStXb1ML2k5K4SlUNtI7
KpnT6mshLr5wVQyqnVLySyI5UzHR61xQ4XO33RAloNH80QQw3YcoDvP8wP+wRR5H8kZEfG9yVHqN
PeYrTJzdAjAK+QpQ8bizSXnNj0GX8Q92H4dS3K6UMPtxtm5aMvp2SZy1XhG2wn37gRfbTRvHko6R
Zy/8sDAXoKAlzVs8Z1OHcRaIk2wdNjbOxqF67QAyxArCh87DaxZtXP0DTw8Bu0Njp/9uJW3gAGWq
ONicH9IiwFxGBqE2FMJfehJ6w3Q+Of/wYjovYLMYKo0KzIp9akg2QoSH2hH/31teq0I+MFndb++c
GMa9EcsmRpjw9e9Z3kJ6nZsFCx7S/bG0enbliEmOPs4magP46NOBNIkYQ+LIVkX8WxiiMYpFCror
1ieUoHyLP+TNw6LF9PfkqGTR3/Sx+L4UKASq7K66o5fLPABW8B/mjkVyEKxONqvsk4t/WZqkvxiS
RsaR/I/iCZPF2pP9O7FU6VKxzSQUMVy/xorJfm3bt/uVeFiUUjfe4eQDqCLv/dmbVjiwKsumw1D+
s9zr9jonsOlVrnlyTRtrOGEPkyUwNM0zDdjrExd/64rzX6tMmpDFHtzMYi2GT4GIrahD+Ho+5VwA
Y1S1BRqnI6hcAQJOvOwLoLF3VKJTX1s+Qj0LCV3zBNm0JLic+qpU1oDAcPnQMgNGGAsEP12x2D61
ArssTCVCieF0PEo2SBxzFSMDRxQHj9jUEhfooATGy8SlH5hFm4Q/mnVz9iDTcVN6dJ6sQOf2jHI5
bpYtpxRlZkqpwzrTxQIrlC4HPGOktNAAPbTLWR9EW2BIWnRBFhABmdnlTXn9EzeD1dpDgYGPliCH
QWDtHsjrNGgRERg3fx6aPltZEx85Y2+YxXQve4GKJpiDPqIIIzbvVHlKKY2hdi4a8JF9BAYrMTx5
vCzbjl1rN7j74omrigV4SDCbOWvbQ7Ci3NxRaLDdNjeEc6J2PbicR5nGzrpGW2kMK1HpcymWWir1
cu4Uic+h22yvuHG+Qvcuo41wfMAOe8fByvfqNeyjOkaUuDVa/baXHqAq5tR3xFWyMRe9D61gTYH1
58RNPsDw3WoPLFspeIMxetnPhGsvRL6VP5nPf+Ffe1pOBnTyt8I2At6Jd8fM0O7vsm79AEYja7vN
NSQkHq5A3gE5QQLQOjd4AnmEG2G3Gu05iv8MbZIrf2Ac0wVztqTRMyi+B+gruTy/Bv0wXK+I7SPl
4dfhGFDJrWzKbPXdWD1NkdL9G9G4Y/YLkV8/6OsvgdJJZkj09eQDVioes+2os3P1ZPmVy8lv+5fo
e3VJb6++MzVDo0Zwl6UcLrutUFU+45F/suSjKBOfF+uAwp1Pc/KrfqtpU87QBiXmsrf4ddYmx39x
30acyYCgAQiECCChMYMQhENT2TQPIlGnvxXlAB7+cScd5+sIXoob+JzK5ltDKNgMDVtX1j1P18RP
ljYjiuHgUPDUHKNYN5qeH4J1Bc85LsbDZKUEYF4QG68aY5Yg7MG4x4ZzJjyKN70muOxvv64+pwK4
Q6+Gg29dtUiqdFusJPVNfUR6Fhv7YrNwUKVLrzohru2oRh6U0T1lzBmGZ7X40YTPypV2MNchynhH
YrSEs+AufCNzrEhz6LltGFZ0KGXLAU7kBwSTzfcEbMggPJQKmiJo1kQHWJJuq98zBZn7II2pHsH9
dkOux/cFUqMSVLEg1DPvFZEuwzY/OnB2m5E6pttAdqvLCrTV6dEmxrRMGFcC82yplESDmmT4xgsf
OBnm38i5Ji63c1qSozOHMsl43Tk2zu2eKJbnpLgzI/d9TZ3pvRB0mXv7ujENgSF+UyqWyA9ixc8+
ilAAKj34RbvnGXZmwXYJ5Efu7l/b3skoRZHMLjaTViPEQ555K/27/vbhdKdvqUr8ykSjqqpnVX+H
CJ1E/oxYwnqOiqNT1zMtDgJ1Hfra6FXgZux4jL5Cx3HiwAbpKzd36TbgkT8aM0xOheb+SZAsvdyR
anj4gjbONq6ghNiP8oWbNQ2007pB+YUAvslijhxCTwglq0IIcr5YR4z3hm6PR8MLhbZ4V6Y2nLJ9
N6qUpIGL41Ocdbb6vyCqZvIq3+zzwYmKoza3L/Vmr2QfPfD0zIWRfzb8+MpdJ9doAM9IqTqczWRf
eMxoQx8JDQSBxPn73LIy2DppJzVJ67Vdg1eyD4TfGtEwMEY9yaJZympVVesNteot+nkDE4zUT4Ij
yc7a5MbXbEVdVjeTCiqNuNjKAaPiGnz7tzUB3+qVtsdWOVypCRNtM0r3HcIQCRGZbUdheygj+UgE
TjiJqCq0CKldhMKVuuueAXYIITU5vtKmhYmTr2fwGP372roHSMrjc6gYmj75UIgL4XDZj2cR/obx
ETmNSk5dYOGo0W1LJQRwsAd2XninJgl+GD3X1tsX/JEcCUJn2BjLsSER5P57+2crzVssHvLkqWVp
BNbodLNK/nyzOfl+ALGq9BbugrLWL48l16r47kwyNOGA1YqvB9w5HGP8ju3L2oPoIqkIXReow2Fu
E/FZaSoEcdmiHvG12iIEoWY6f6UXAUeQL0TGoyK153nIo9HcUrBhoCrLf3PWxxGE/3qldzuli+4o
vp4YvCxDGt5cRzucoQET2kn5hb+Ir/zbUHhK2OcD1pRlL4CetgATzRALIMgxMHDOepb6hDo2vCJN
03Rn54uMYP+OeuHgQzXevQL9TxjtALEvjM3J6UCf7g9wD/KKZT8Xtptft7vBgW4PDiq+ur6Urm2u
Q0NU1P2m6Tilfr5UKx6u/I6NM1EVJmOLpdHrC5qB8qk37//5NLa980fgeUtpdcjvrKv3QDuUqEwr
ha0Ym3q1/8BD82ENm0+AtNOG7pcxCJYbTqJrUeDbn8w14BIR0Mvf8me+jvzqumLTaEcftseefqMH
f8TXKpQhFDMYIFUUcqBchZA6xF+YstcBZpKo0NHbLzhXZa3w0E1XVhyjJ6xWFLAPP8lQUa1HESP4
sAySpdL9llyBA6CvK5442z+pLr4r6g8dv1NVgF6+ERNbQ7Ex5I/uh/7RrJwJ0YWV9FBQItzITlG7
OO42lYSRcjVsHYmwPofvvacBJ76PEkj6034zKR11HYW0yDJgBwLROJqiXM9gwrvo+bHx3K/XQEsO
l2GhVWDyPDUSnqxYsmhnemP7fZxYaZN+ajLersyQ7cYQcdZzwhYvyfpuK+XE9J1jRDtvcAPr1CL8
RRMY9m3OnOY0AlYQDw6QzCQ0lS6gRVPocDIhHcsd/m+M+vmuNvl5B3gRH+dFQkX6NCwWt/H3/jNP
ZQ/leb1m8x+8wYrGZUHN/IuIFQy8+BBWMMo6ZhJih2c53CCvJWfCpJ/ADhldN4e/ASi+6vgVmAp3
Pta8L5/Csn/2fI9K+r49ivoufk/E0NCLRRZrTIy2q6bPsZ88iRetgyeaCm/mneY20VPllSnRZWJ7
l0DGXlQh4FcHgya6/HLY23dUQ6oF1d3h6vyelc+yMwxzHmmuyDzG+vcvDWLrrzBGTfEQGf60rkzL
o4tJ614mvw+hmulJw4iLZRCawyyoymCk4k1zrhCskI+rLG+jiJ53CSw08MS/osoBWVlOaNZ3Q8KJ
AkynigkJlBx9BU0VrWl2ru2n8GfUWdaIRgOcMP5ZgOcvkDQciGjCLRfxIYPOt34W5/cL8P+nv+GO
xidsO6cNOzFq4z3Ze6p/bO5IPMu27x/ri4MFO01ZeA46SYktouhaI4qH0+xa7VE0ea3PhNsiTpi7
o4nMii4G5DcjeY16BM4HnPkRhfrCZRcsPoTVfdIOX5tfQ4IybVBErrzZO4hzDoVo/TKVwlE/22Gm
84rP516Ng3rqYLow4sYP1n5p4bdLQRGtOCkSbvBctTS3HmuNOqpt0pjg0dhXokj5WuGlph5zCClC
qRaJS1iKf0/2wdjbHkcxRafMwGdyxbcCEu/ZXipk53w364N5+AQS6+6dspZ26vii8oG4/81GL/Ai
geP6MvGz3YgGP+Of452uMCOTFDjqxQkyp0/jP0vIcPZIUvJFnYyojn0QjVAR1N6S5Ebiswmk6Sls
YLMeRDFALtUcnHADTnk+uZ04JRNKpadORnhp2EaLK7uRlkBD6FgKKQdVTpgDjMw1VZsnLElqpDPx
LH+zwJtblcLzLl4KrkhrOZBxzFzmcG/Wy0kLh4YH2qk73qh9bCE6gwbmzFVQ6mmgGqqhGybRw2Mh
R7ON2YpmizeePv6N5XCbbBN4M5TKFROfqTlhSzHvuCWJIIgr9W6EPmbmZ9DjIJIL5w5TuIvIkMcz
Hxl2oUXyuG+0/zcbR2ohFZOp/DO2s9TSimENFfAneDoECpFH2RNmPQSb7ZB3uIneSvjXczh4OqyX
hvy4DJMXtx+gg8sPA3ygJle0ZSiCW1USdcQjQy3gTBYv9gfY3sDVR8NpDYOmrjbqHeYaKSV0IuB4
oJv3bSdjbpB9qgFTy7LKDfvJYGeJMvTr7HJgtp0qxFxkwR8klr01B6NoCCf8Bu7AVv6YtVGy88RV
+Yv+YvHrsv6j4+Qmxn8gH/ZjrufH67jKczR+kbalomL+nTlzjZcGjamc5XBrlxDfIoOAI3Hye0GW
IQA2BShXmpNrBNCzFChroZTdE3fk9KTS8jIxOUYkOsMGkKkgTUzeiUA3+q1gzYbtuL9L0Tz5ul+S
ZfzRnJrnMD7ieTisPjFceL1i8iUpXrVb+bt7K+kASgMDSaWwGeK3odLvCwp2SH4LnR6ljQHA/DEG
0w5rfhcz/eL2qwRQTYEJtFJMP4dTZbrtF/F/WimtEoeYlocQWEs/nthekqBed7Ry6jkvqkiidjx7
zT8F0OyY/IXDKeyIDhQfsjDAVIWjRvdMj6mQpjXdXHx1TZhuP6nSkolHfmVnY9MkOMBnf/eyY4kx
6VK12cQtocQAsleHkW9QgoObz/3Wl9JLlpD6a7CV2JVcIWjvrjAfFrXYjo42uI0IUZU+R6ScIwIm
gpMG7+WbUn8kTj9d+S7EKe0Xc7G2hSIBIKd+NO690htK4dvpxCSuUNYenPlnE6zQpRcrnBJ+pgv4
yS4ExYUqoyL9d/8j7k5aEJT1qEoAS0kGpD4vEinP9mQiZq7ZtsxbKuz7A7i+8tnZMJQeBHu8EzrT
gIWJ6j7QISZ1oe3psYoDd42khzGZMYM3ZKa10uLu8aOfUyBuJrarDkLryUR/ZLYYzaCJZ+4hFgcH
AJBQlwmZI5tBn2ipRRuunr0RSmTyhiMKVeeTjGIT+ZB7pnXlWjB4cRDDbypCRFTR9TfwFB5E9j/o
cUXolhl2+7Fp9VAUT196qkin+SU3omX8QpyTrYl54Ro3wuyMzURcZ2pjFgjLg1EoJcRMSEGVNKmZ
GabcEL7piPynOt4MUDn3pRkagVctBNIwfDx2cFmP8aJarO0CMKasgg9hBLeOzcsqpnLYP3PDbx0w
sgs8ibUV1tt82Y/KTgwsdadtDuzUAEUZ2B9ecgDUs5qZMZh12Tggznnp38wiBU/CzPYXKstqxyE3
cfE89n78cvIqEkQjPZUmVl37TySerHjeVxnTY7cc0mzdEusNZmycjS7VrDLgRt5tHdx1vyvEsBev
c/bzX0nxZuazwmtDsEiWhBhsQIVeBMyOLZJauwgHX9L00Zd/oLTWpTX47XCQSOiVASEaZAHPwZaR
NDaWa3DAAMHiGGfv9AamY7bUN0UNPFLj6DOYFBITIrUTlcO44JdsjbpMUtbS7pP8c//vXF3jiKSO
N/jkUVdrB2j/2ZtoTgPDm4sfhrkAzBEVo3fp7j9Bjn3w5pW6Q+sC/IN2XJYu+pAdApw6jlnQbc6g
fP9N6hmCK1ylTCiU1eRBOBEL3eM85H5V+87yiLFkUAZY/4BG1arCS8icWvTJ1TagyYlFDwiTD9D0
kiayGj7xpB/7lDz9+nqNzOBjZi/p3rTV64bToIZ861ssAH+zP231EpDZVkQkR47B5j+KcjISRZ4G
kKY8HiZGE3lE++y1F5grvqtxKIIUdy0dJgB7lrOtSuGT91rAkIhqPyoZZauHMHOH5Dkfv2G5zRHt
nbkPgKEszYK2H4ggrPkGmhHmLzBGuevBumJzjauwN73keDNrW0poJcB5qVZv0lF5z+qgAzh/l//i
9AVgsEci7Dq+d4r1CUxgFkMUzY4G+U5Y1ibLFQLvvjTtCZJcO4HcWZFWmSoh6D8Sj96EmNB/97gR
mxSQiBHW+JtxXBQpeArsWBrXSL6V7T9QaP4rbXbYcCnHIS3BQCRMPlOYAHXEsDw/7ZND5iG/Vm64
XnO/rgFr7DA7Q8BKmJSYnRpDFpz5ZZtOJpLPFnGuP1G8xDmq0IME7glZ3DxBxFN2PA5om+ig/lGB
VOF+GT/0Ei5rMljGdI8s+4OTebTUPCNNX43ZcJRn3IeQFZY/bj/eKjJFXkJIaFm/SfJd9Bhte7+h
brwfBxe9rjXy1TWDU+61MwmOh+vv+pa2TbPFrSmIuwbQw4G3S9YmEFUbUuFvCIUHEiqAj5Lm+Wck
4P4G3OckrDX2EGyhKdpzAlIjIg261UymKvSr3tzcsR1ZT8WNLXaNkSfYXSPmvpwm92aTAM0tvsg0
gLU596PeLkYfhbI2SFT8d27cNRdmwcyz3nt3WuVsnjr+npnkjH4GQnaRojGj/qSDy8untmW1euYF
WKL9COUMdsTgB6eDnYqNz+JmIdHzRXhFFEV0QCoH5tM2CNSZLWH4o1wgqERoWnV1e2i0b0xjtbzL
SgFfXach/MUk36jJuZ4j8pxiLfHxThcmTbYHmAPISvet47NjhElZyfx3IUiVZRBaAuvLqqCYxkmJ
xf32LSzFWE187SXQd/lx0kkGYgeo6I13J6A7238YdOWXTJUkdLmWAxKqqbQ31Ye5ewZLfA7Rs8t0
+dPMR3qG6TnsvqCRhGNRlxgCi3MJXj6i6BbuUdqjCUZi+MjgDxuYGh1L+eIZwfcBfpooXBZhjvMF
NHBJ0DbDC6jUjHiLjn/vh8OAKoSuBAD4BvbDhk4YqV5mu7FttHaScK7NfPVRUox0opVaoO37GarH
CwvnAQqQD27mBUBsuNpx8if6eaZ1QSKkXTCdRdUc6k7wi8DLB5vylkH0YS+0gyL7jIBc4yer1kQR
ZrLhKC/y+te/yeta6IBvhrHizk6vFiXyssAVbOwRpkFOI8owRFCsxf/ITmuIma2NOsuxM9pV3O9+
vPAGRecCSCe0SqmapTK4xU0FBtwp7JZW3ocZeIrMO10VdJSEIBt6LJL8SeOWKH3Qmw2D+DeC6I7j
1DzDKXTgcKDtOp7Us+7B6cg7XU2JmJOlPQf4P1u5Ur985pEtUlprRIJVScP13dN2zb6Fk2UQvT/A
q3mP5kRpZDlgMz2zVgG2b4XYbPJ3R87r+isgqVWGMbvo2Y6lzETNhZfbOD/oy9GQAIjdBpgRtFWP
4gvgpgRRVhCaxQiDV3kAgIvs+5/z49pM/PIQ7Jow3HUOBNiIC4hXp6Q6UJOSfUIn72e8YRvnz1Wv
ihXuE2FBfVfePsQQFXKSNSxyv4CmRRO6VzMBFD2PyuGdG8EztXQPi7zIlBIr3tjvvsOG+JEzuHo9
2sgLZIJBnxBWrxMYvcUsh2KPUG47nfzMQUpitZqrfw2gDBjCAFhPA19J+jz78m1qi+Qo5xLu4HoF
woyVwAUK5RbbQzMhdqe503OcYLOetOtjpwTjh8h9wXkfEJi8Lu/lQH3IP+p9sPFgPwaVzdeAc5pT
m5voFucGZq4UfqpEf7OcZJKKz5WFceC8yKe7YNepfHF9LDoSTu1Dl36EuUfGShGCn71208mWSJz+
cC1tCbldh7a8FMrFyxvopd8vzUwzvC6avdvsk93irQ7crv/QJCPGnHekg45XeFA54Nawhprpyqi0
peC6uKWHZvDd+zabfMrRI45Uk6X/EDhmjMQ5Pf9NBQ7i8SLuYB/k8yExQg0YC/1x4wEDJl3JfZK5
jik+77mHZvwqKcc/3iBF3csT0DxfSmR4VFtHVhFX7C1FburqtpQzJ06IlW+RbOzmkI7W64zc/1Qk
r9393bG/vMrZ8wmk42VJSsWKfrrMtkUGojYUBsTylUmNpaUlFOAOS0XC6ovpui5YMGF6nQW1XSrc
OSl+t+AMnKyOnP0L0itBZUeeRILMBQs2MzEkgjjSHi+covGNqZxwz8eES5oJK2qSl3KiDE1ZG6+v
xrEAoHpt02whhTkvnnGK+xMIDb7kQCs+hfYvLxQNwgcbTfZan4EHb9XHxkTxtkfR7g/yaMJHCT41
Wzr0XB/S01ySDvjZu9l74bWzfiFvqEOCv6usw4TmKJvhdEKvbI2SgQJcQ3WlcBElyTlrvJWmyc4g
9qImw9rJ30RL0WdMoMluQhSzbX6BZcEDgXWQx4SHq6u1it+OOr3pU+HKui7zxKJyW4vWDP2pnxLz
hf2Xcq25CW0G30yPmjIEdFT5tYkOR4nN42R8pEe2VQdpocPVOhjd9mVmfy7cnbmRLJfM8Ww0ArC9
1XM04tv5otvKKLM4w41MWhrK7gKk29kaXrHRMYOVMD0WhVPXAbkVIsa0Cl0LQpfADTu6abE5+Qvz
rne/M10s8mmW2ajy5pzuPwvmJ2HUenih7cLbstr58jC82mGd4N+muEd50FZ6I7aF0FIj00qm1Hr+
Bng9IVG0N7975JMrn8ImMFgM7ubHrKVX33ZXr9eSn64RzkMIYBMIFCUcHdMeeOFwZ0+J+w21hhAA
xyris60IUsG2fThz2sFEtOkc6BzredJjFin6tdy6sUvLlKvMwZmV/cniYugVuwcaItGrjOiyWvxI
tzMAS2iDoBv6ZCIBpFUrQcnc/XbACxX7R9wrFO2MC2USicoILURHYw+VXkzCLMPzZfi1h+g36eUj
KRy+tNsyeDdSHqUD26qIDG9IH4i/hLEzyQHplo9OzobKckDs7KzSwp6lkTgLQiig27GP4fD00GOQ
+hbdlWVfiultC3S+hPjKb4B+Dday4JdoQVU5OMYQVgN0iVw+mWkYgUhSKzNQDwtSx105AeK4oPGb
BTKPklH5HIJ/ueuAOe7dki2fs9xGSI/lYkrsxsA7ySSjNaoOt8RIJEIP61z2bHIvIz+gW9PERcKq
v3R73GMCFmSF7IGBNa491D8uGxvT4VvsCZyy68QhX/DasqasU/3qa6ACdOkowupxUEqYfoxKhn0I
3AVPrM+n4ihf0MDTpRsupiehXWe9eJz0jEyr6NPNYfjrSWLrXTAnoDuucAcDiI6xPyC8DM9M0svW
kM4cMBMTVWd0WIuWPi+BTg9pxdvfZZ7JySkuF+IoPzcACHGiHgUls2vEjZGt++n31RAbUTJ1uwGZ
3M+VVy7kh0M+hnJlDFHTFdM4bSs61wHfq2zbzgziJTYorS5fX+OWy9gY0ci7YzvpRnO+edaMx+sq
CYgq+HE7GC4yuttHMrSwGFSa1FM7vEqKb/VAI93Gs44HKRKmVndCB2S4zp9M6jOhBXWbM68BYRgX
G5V3j20WDBXjBTz9wnGlfRjl+AYUra4rqya4X5/9HdhVR+SDDf9VFUHvkGBO8dqXgPxw8d0oeSrV
xAPPI5QJRca8p8M7K0Y2PG4gsuqTTwbgJBQv3kcwCLYfisf5iN1uB0vtpSdAYDP92jZZHuqpBJx0
j5+SUkTRTmNLArGMuafXV7zrZEM+TA/7yVZreGokKjEayUc3mylElX7Yqz7BsL0vnk5qrjR8DxPo
gbPt6r5YGYX1WcdTBDdM+Gv1VojGQTEgxMg2s3BAsChIXXqsLlEVzz5xLlB43Wywqpf1/bU/uM8J
nEKnabTitcSv85c7oHDEr4RoalM8spUc8PJ888h8c26p0wJKd+ceAegsxwUCPImbs9h5V3oKf7X/
fksDx/ATxYom0MvI5WdxhLQ+F1mLdn0n5sy/6J16sHJOr+ivtl5j4n+LHVo5GEuZdJlqr2n7sFFM
RCofh789bcMVi5LIizLm9GH4d37vQIQhaAR60gOgYdHWE5zl0iLEFTJCIb46GWXntEzbVc2ld1dR
3NuQVmFW3PKptVquSxabaokSGG6vNxENft7h3XiL0u7JGWTBm3/mB0dFXq4BTfwOxvpub/n5nyRZ
2gMb20DSCb4bJ/Z5pWAMvly77O908XhW4MIOEHpgoL53xbC5oWUFCL1lNmYWobgU5QRIAXHX48W/
kFkFCng5ZSXaKuLkQTx4oKcPaJoajqAnmTLdZJhElr12hLYLDaifTj0HTcQlfMrC17i32aw3eQ5h
czTi0ut/sav6bxxEPt7cXe3BMB8491wQ9AiGJV8uGFCPro4BxVc+Uf9D+yXGrtdmCrOlq+DrlnD2
jlJSzR1vYGZNbI/+BpR5UBL5TEvr2I0gkTu5DlL9ce4GcZPAHukm1aCY6ZyPiDuFbMfPrROf5XIR
rhIJmWuDAIYtH7pJQcVIU8uV8DwokVTSIYL1amDS+Pn6XFWmB0P0yzgFduK+zJK7OBgzq/Ea/r3g
DfMq3HxgVBB2n9i5bmeyzcdJHUxmHzD+iKSkwnHs4cwp+pz/zBIxE6phd2k637rXqoeIrYeJhFH/
BtDLzLUCPrBN7DAlwbu9p5g0wOfjcywXESlFWH6I0oAO0LfM4jXmVkCqVKTV8HQa4nI/fRaXOb97
jrJ1tNgrP3FtvQ1wr/wPXOdbmxPNc4FQz5ZhY0SAodrUW+89gfoAXl6eBrnDlwQvntyVR5SYmfln
XfjufXt1k/kyynRc9ucksOGXejPi9D8gNTn764aem3p7tlKtZowJ7henzPRbJ3XrPKfNdZw0fys9
Si6B+cFosJpqcKkpHNbMvRxJQP14E4jsUzoJi1ZX763nvrIifLUZndTw25/SLDNUx5tU7n12r2dN
SolhruU0hRpKcspXoIMEb0GW0gXi/VzN4t4Et2PhknLqf+T/Mc2GivLTSqDEk3ZUYkjAFnmMlAfk
ZOauA3eOeYiFVgFqIZnTSL1mfinP9K4qm4RhZsiulH77I6C+rCh5SxnzDDBaVFC5mZfBhQi/QPKD
Np8jdUHXxy3nzhIkhse7VArY87PfA3mk1HBFZMcBBI1tnKcoWKeUg3FjGIUnysYUOzJGA3IURsNZ
EioGz4jYUVQszjVCunI7YSP3oUVnl3m5jTSTvacQ01BLotA7yyNENO8F3EHN2FUeBRtE4gPF2Gpc
UOPun988Q3xaCmnvX7pn9kxf0mKfkMrphekcOc3iJryLmmWTTiP8eG8je7ZRTbRpGvex3UMw1iNw
Ja31BtVqc3Ax62qS14OgJzDt4f167rjt8GSJeoYrsk0tSEgbjgbiktHEQ8lnR3aM59+ZLKCi1w02
a9ICxRulXv1AwZOtFSLE+W+NRx8zWV+CINllymp1d8IQPsg0GOGJ+fNvp5LsrRjXVsJMJ7zGdHeT
tD5IQM7/5Xr8sM8ZC1sHaxj4lqk+gJ0vAdrZOboKNdeK7rt3NNoD6e4vKkMmYJWYxp5RvOW3kxSu
bu8LpqV3amEag9JfhufpXF232GeDvzKKqn+xSCt7oG/jylzMHQ4EwLouTgRrJ/ZAdmmVu3yJuVBE
/B4mKnUG9mBoK916+Oha0jF2y3mkwrNfXY6UEEThNG2gU4TsWfbkaqNJhdKldo31TaTU2tDeeFlX
Pz+/xnJCZh6q91qXVhDyaJVz1ArfFVUkTQXF0OgjRdTuCWCGVxx3u1w2pF5uFsvWsdGNZiAnTon0
hA/qv1KZw9RfPP27jidJrHXE2kux3IU/fuW0K1dHUYxv/CZm+BrN3Dgcll1B3VcY5hTaAbheYuqi
3UJ0GZhPRe9IDQKwqmZerNblmvsIUPBm7rIKQ+rx7aZi6XEKxrNbCdW64M0LP+CshCbzBeJAdfAE
JF6nS0k5tvG4zIqIS+r/IFdWrJiX0OZbwbFgROnQpJYccDL+GkYpliobSUEJhFKfwp/5jDoKKz21
+zM2KFwNQOvijuyPAT48p2cc5tCItJXOhloz1wfmibjm6sRSBC45AL39LRiMBARKjAz2M0wBY2o6
MNLOTBPMDodU7aPfCYTTrQpZVOd6tTrb5eygBE0kL4uVKWCE3fgWGLdW0Wi4GNIeU4URcn77riTU
vld+Rvhip/z6cFXiu4xficv785MPhlpPAnG8TJxT3s9kECpWaJr5vMidKQ2xVVS5e8mGUNgKHyaz
WxBV0svZrzjbfngrV6puBUDCHyJsKluTM6zUcY0Uahl6EPNO/zOCb/OHhNtDw3UUxl2ztwqymjnL
dY4KrSxnBk9fAf0TvlAK6HiafwaQQOSxorA4SFQDB8B7fLmh/aemmSbWd4Q4WPXuDRhw4CaNyXWI
+IFdG2HpUa7yeeSLbIzaCsHoXIVe+cKRdU99cXTy7CqlG+skJSjT4wJArf6IBZestr7Lc6OtUrJX
KAWUhO6XC70PkUqwOqTdTMLzI3LsfI5NfAtJMZ01yg6fSnPZDrZhTbA7IHSP
`protect end_protected

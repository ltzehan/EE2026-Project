`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.10.2022 17:57:13
// Design Name: 
// Module Name: sim_goertzel_mul
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define assert(signal, value) \
	if (signal !== value) begin \
	    $display("ASSERTION FAILED in %m: signal != value"); \
	    $finish; \
	end

module sim_goertzel_mul(
    );
    
    // 100MHz clock
    reg CLK = 0;
    always begin
        #5 CLK <= ~CLK;
    end
    
    reg signed [60:0] a;
    reg signed [60:0] b;
    wire signed [60:0] y;
    goertzel_mul goertzel_mul(CLK, 1'b0, 1'b1, a, b, y); 
    
    initial begin
        // a = 2619.305006107305
        // b = 2377.677142872972
        // y = 6227861.64323409
        a = 61'b0000000000000000000101000111011010011100001010011100001010101;
        b = 61'b0000000000000000000100101001001101011010101100100111100001111;
        #10;
        $display("Expected = 0000000010111110000011110010101101001001010101011111101010001");
        $display("Actual   = %b", y);
        #10;
        
        // a = 2430.4977668807733
        // b = 2404.3504052031617
        // y = 5843768.290645167
        a = 61'b0000000000000000000100101111110011111110110110110100110011110;
        b = 61'b0000000000000000000100101100100010110011011010000100111110001;
        #10;
        $display("Expected = 0000000010110010010101100111000010010100110011110111000110000");
        $display("Actual   = %b", y);
        #10;
        
        // a = 1108.2091204349908
        // b = 1511.349611345804
        // y = 1674891.4234592987
        a = 61'b0000000000000000000010001010100001101011000100011101010101101;
        b = 61'b0000000000000000000010111100111010110011000000000100001000100;
        #10;
        $display("Expected = 0000000000110011000111010001011011011000110011111010100000111");
        $display("Actual   = %b", y);
        #10;
        
        // a = 1838.1458222179713
        // b = 2991.7721948171525
        // y = 5499313.560931039
        a = 61'b0000000000000000000011100101110001001010101010010011010110110;
        b = 61'b0000000000000000000101110101111110001011010111010001111001111;
        #10;
        $display("Expected = 0000000010100111110100110110001100011111001100100101101001101");
        $display("Actual   = %b", y);
        #10;
    end
    
endmodule
